VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mgmt_core
  CLASS BLOCK ;
  FOREIGN mgmt_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 2250.000 BY 740.000 ;
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 91.490 2244.340 93.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 221.490 2244.340 223.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 351.490 2244.340 353.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 481.490 2244.340 483.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 611.490 2244.340 613.090 ;
    END
    PORT
      LAYER met4 ;
        RECT 96.040 10.640 97.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 146.040 10.640 147.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 196.040 10.640 197.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 246.040 10.640 247.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 296.040 10.640 297.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.040 10.640 347.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 396.040 10.640 397.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 446.040 10.640 447.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 496.040 10.640 497.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 546.040 10.640 547.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 696.040 10.640 697.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 746.040 10.640 747.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 796.040 10.640 797.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 846.040 10.640 847.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 896.040 10.640 897.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 946.040 10.640 947.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 996.040 10.640 997.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1046.040 10.640 1047.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.040 10.640 1097.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1146.040 10.640 1147.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 46.040 10.640 47.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 96.040 518.260 97.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 146.040 518.260 147.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 196.040 518.260 197.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 246.040 518.260 247.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 296.040 518.260 297.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.040 518.260 347.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 396.040 518.260 397.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 446.040 518.260 447.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 496.040 518.260 497.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 546.040 518.260 547.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 596.040 10.640 597.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 646.040 10.640 647.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 696.040 518.260 697.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 746.040 518.260 747.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 796.040 518.260 797.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 846.040 518.260 847.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 896.040 518.260 897.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 946.040 518.260 947.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 996.040 518.260 997.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1046.040 518.260 1047.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.040 518.260 1097.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1146.040 518.260 1147.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1196.040 10.640 1197.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1246.040 10.640 1247.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1296.040 10.640 1297.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1346.040 10.640 1347.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1396.040 10.640 1397.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1446.040 10.640 1447.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1496.040 10.640 1497.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1546.040 10.640 1547.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1596.040 10.640 1597.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1646.040 10.640 1647.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1696.040 10.640 1697.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1746.040 10.640 1747.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1796.040 10.640 1797.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1846.040 10.640 1847.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1896.040 10.640 1897.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1946.040 10.640 1947.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1996.040 10.640 1997.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2046.040 10.640 2047.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2096.040 10.640 2097.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2146.040 10.640 2147.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2196.040 10.640 2197.640 729.200 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 2244.340 28.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 156.490 2244.340 158.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 286.490 2244.340 288.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 416.490 2244.340 418.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 546.490 2244.340 548.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 676.490 2244.340 678.090 ;
    END
    PORT
      LAYER met4 ;
        RECT 121.040 10.640 122.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.040 10.640 172.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 221.040 10.640 222.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 271.040 10.640 272.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 10.640 322.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 371.040 10.640 372.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 421.040 10.640 422.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 471.040 10.640 472.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 521.040 10.640 522.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 571.040 10.640 572.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.040 10.640 672.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 721.040 10.640 722.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 771.040 10.640 772.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 821.040 10.640 822.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 871.040 10.640 872.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.040 10.640 922.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 971.040 10.640 972.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.040 10.640 1022.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1071.040 10.640 1072.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1121.040 10.640 1122.640 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.040 10.640 72.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 121.040 518.260 122.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.040 518.260 172.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 221.040 518.260 222.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 271.040 518.260 272.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 518.260 322.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 371.040 518.260 372.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 421.040 518.260 422.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 471.040 518.260 472.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 521.040 518.260 522.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 571.040 518.260 572.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 621.040 10.640 622.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.040 518.260 672.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 721.040 518.260 722.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 771.040 518.260 772.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 821.040 518.260 822.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 871.040 518.260 872.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.040 518.260 922.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 971.040 518.260 972.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.040 518.260 1022.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1071.040 518.260 1072.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1121.040 518.260 1122.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1171.040 10.640 1172.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1221.040 10.640 1222.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1271.040 10.640 1272.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1321.040 10.640 1322.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1371.040 10.640 1372.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1421.040 10.640 1422.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1471.040 10.640 1472.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1521.040 10.640 1522.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1571.040 10.640 1572.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1621.040 10.640 1622.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1671.040 10.640 1672.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1721.040 10.640 1722.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1771.040 10.640 1772.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1821.040 10.640 1822.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1871.040 10.640 1872.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1921.040 10.640 1922.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1971.040 10.640 1972.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2021.040 10.640 2022.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2071.040 10.640 2072.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2121.040 10.640 2122.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.040 10.640 2172.640 729.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2221.040 10.640 2222.640 729.200 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END clk
  PIN debug_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1980.850 0.000 1981.130 4.000 ;
    END
  END debug_in
  PIN debug_mode
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2000.630 0.000 2000.910 4.000 ;
    END
  END debug_mode
  PIN debug_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2040.190 0.000 2040.470 4.000 ;
    END
  END debug_oeb
  PIN debug_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2020.410 0.000 2020.690 4.000 ;
    END
  END debug_out
  PIN flash_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 0.000 188.970 4.000 ;
    END
  END flash_clk
  PIN flash_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 0.000 169.190 4.000 ;
    END
  END flash_csb
  PIN flash_io0_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 0.000 208.750 4.000 ;
    END
  END flash_io0_di
  PIN flash_io0_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END flash_io0_do
  PIN flash_io0_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 0.000 248.770 4.000 ;
    END
  END flash_io0_oeb
  PIN flash_io1_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 0.000 268.550 4.000 ;
    END
  END flash_io1_di
  PIN flash_io1_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 0.000 288.330 4.000 ;
    END
  END flash_io1_do
  PIN flash_io1_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 0.000 308.570 4.000 ;
    END
  END flash_io1_oeb
  PIN flash_io2_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.070 0.000 328.350 4.000 ;
    END
  END flash_io2_di
  PIN flash_io2_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END flash_io2_do
  PIN flash_io2_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 517.520 4.000 518.120 ;
    END
  END flash_io2_oeb
  PIN flash_io2_oenb_state
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.650 0.000 407.930 4.000 ;
    END
  END flash_io2_oenb_state
  PIN flash_io3_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 0.000 368.370 4.000 ;
    END
  END flash_io3_di
  PIN flash_io3_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.870 0.000 388.150 4.000 ;
    END
  END flash_io3_do
  PIN flash_io3_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 511.400 4.000 512.000 ;
    END
  END flash_io3_oeb
  PIN flash_io3_oenb_state
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.430 0.000 427.710 4.000 ;
    END
  END flash_io3_oenb_state
  PIN gpio_in_pad
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 4.000 ;
    END
  END gpio_in_pad
  PIN gpio_inenb_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END gpio_inenb_pad
  PIN gpio_mode0_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END gpio_mode0_pad
  PIN gpio_mode1_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 0.000 109.390 4.000 ;
    END
  END gpio_mode1_pad
  PIN gpio_out_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END gpio_out_pad
  PIN gpio_outenb_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 0.000 148.950 4.000 ;
    END
  END gpio_outenb_pad
  PIN hk_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.450 0.000 467.730 4.000 ;
    END
  END hk_ack_i
  PIN hk_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.470 0.000 507.750 4.000 ;
    END
  END hk_dat_i[0]
  PIN hk_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.190 0.000 706.470 4.000 ;
    END
  END hk_dat_i[10]
  PIN hk_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.430 0.000 726.710 4.000 ;
    END
  END hk_dat_i[11]
  PIN hk_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.210 0.000 746.490 4.000 ;
    END
  END hk_dat_i[12]
  PIN hk_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.990 0.000 766.270 4.000 ;
    END
  END hk_dat_i[13]
  PIN hk_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.230 0.000 786.510 4.000 ;
    END
  END hk_dat_i[14]
  PIN hk_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.010 0.000 806.290 4.000 ;
    END
  END hk_dat_i[15]
  PIN hk_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 825.790 0.000 826.070 4.000 ;
    END
  END hk_dat_i[16]
  PIN hk_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.570 0.000 845.850 4.000 ;
    END
  END hk_dat_i[17]
  PIN hk_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.810 0.000 866.090 4.000 ;
    END
  END hk_dat_i[18]
  PIN hk_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.590 0.000 885.870 4.000 ;
    END
  END hk_dat_i[19]
  PIN hk_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.250 0.000 527.530 4.000 ;
    END
  END hk_dat_i[1]
  PIN hk_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 905.370 0.000 905.650 4.000 ;
    END
  END hk_dat_i[20]
  PIN hk_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 925.610 0.000 925.890 4.000 ;
    END
  END hk_dat_i[21]
  PIN hk_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 945.390 0.000 945.670 4.000 ;
    END
  END hk_dat_i[22]
  PIN hk_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.170 0.000 965.450 4.000 ;
    END
  END hk_dat_i[23]
  PIN hk_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.950 0.000 985.230 4.000 ;
    END
  END hk_dat_i[24]
  PIN hk_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1005.190 0.000 1005.470 4.000 ;
    END
  END hk_dat_i[25]
  PIN hk_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.970 0.000 1025.250 4.000 ;
    END
  END hk_dat_i[26]
  PIN hk_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1044.750 0.000 1045.030 4.000 ;
    END
  END hk_dat_i[27]
  PIN hk_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1064.990 0.000 1065.270 4.000 ;
    END
  END hk_dat_i[28]
  PIN hk_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.770 0.000 1085.050 4.000 ;
    END
  END hk_dat_i[29]
  PIN hk_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.030 0.000 547.310 4.000 ;
    END
  END hk_dat_i[2]
  PIN hk_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.550 0.000 1104.830 4.000 ;
    END
  END hk_dat_i[30]
  PIN hk_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1124.330 0.000 1124.610 4.000 ;
    END
  END hk_dat_i[31]
  PIN hk_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 0.000 567.090 4.000 ;
    END
  END hk_dat_i[3]
  PIN hk_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.050 0.000 587.330 4.000 ;
    END
  END hk_dat_i[4]
  PIN hk_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.830 0.000 607.110 4.000 ;
    END
  END hk_dat_i[5]
  PIN hk_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.610 0.000 626.890 4.000 ;
    END
  END hk_dat_i[6]
  PIN hk_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.850 0.000 647.130 4.000 ;
    END
  END hk_dat_i[7]
  PIN hk_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 0.000 666.910 4.000 ;
    END
  END hk_dat_i[8]
  PIN hk_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.410 0.000 686.690 4.000 ;
    END
  END hk_dat_i[9]
  PIN hk_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.230 0.000 487.510 4.000 ;
    END
  END hk_stb_o
  PIN irq[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2228.790 736.000 2229.070 740.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2232.470 736.000 2232.750 740.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2236.610 736.000 2236.890 740.000 ;
    END
  END irq[2]
  PIN irq[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2240.290 736.000 2240.570 740.000 ;
    END
  END irq[3]
  PIN irq[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2243.970 736.000 2244.250 740.000 ;
    END
  END irq[4]
  PIN irq[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2247.650 736.000 2247.930 740.000 ;
    END
  END irq[5]
  PIN jtag_oenb_state
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 185.000 2250.000 185.600 ;
    END
  END jtag_oenb_state
  PIN la_iena[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 736.000 2.210 740.000 ;
    END
  END la_iena[0]
  PIN la_iena[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1519.470 736.000 1519.750 740.000 ;
    END
  END la_iena[100]
  PIN la_iena[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1534.650 736.000 1534.930 740.000 ;
    END
  END la_iena[101]
  PIN la_iena[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1549.830 736.000 1550.110 740.000 ;
    END
  END la_iena[102]
  PIN la_iena[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1565.010 736.000 1565.290 740.000 ;
    END
  END la_iena[103]
  PIN la_iena[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.190 736.000 1580.470 740.000 ;
    END
  END la_iena[104]
  PIN la_iena[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1595.370 736.000 1595.650 740.000 ;
    END
  END la_iena[105]
  PIN la_iena[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.550 736.000 1610.830 740.000 ;
    END
  END la_iena[106]
  PIN la_iena[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1625.730 736.000 1626.010 740.000 ;
    END
  END la_iena[107]
  PIN la_iena[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1640.910 736.000 1641.190 740.000 ;
    END
  END la_iena[108]
  PIN la_iena[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1656.090 736.000 1656.370 740.000 ;
    END
  END la_iena[109]
  PIN la_iena[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 736.000 153.550 740.000 ;
    END
  END la_iena[10]
  PIN la_iena[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1671.270 736.000 1671.550 740.000 ;
    END
  END la_iena[110]
  PIN la_iena[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1686.450 736.000 1686.730 740.000 ;
    END
  END la_iena[111]
  PIN la_iena[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1701.630 736.000 1701.910 740.000 ;
    END
  END la_iena[112]
  PIN la_iena[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.810 736.000 1717.090 740.000 ;
    END
  END la_iena[113]
  PIN la_iena[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1731.990 736.000 1732.270 740.000 ;
    END
  END la_iena[114]
  PIN la_iena[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1747.170 736.000 1747.450 740.000 ;
    END
  END la_iena[115]
  PIN la_iena[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1762.350 736.000 1762.630 740.000 ;
    END
  END la_iena[116]
  PIN la_iena[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1777.530 736.000 1777.810 740.000 ;
    END
  END la_iena[117]
  PIN la_iena[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1792.710 736.000 1792.990 740.000 ;
    END
  END la_iena[118]
  PIN la_iena[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1807.430 736.000 1807.710 740.000 ;
    END
  END la_iena[119]
  PIN la_iena[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 736.000 168.730 740.000 ;
    END
  END la_iena[11]
  PIN la_iena[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1822.610 736.000 1822.890 740.000 ;
    END
  END la_iena[120]
  PIN la_iena[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1837.790 736.000 1838.070 740.000 ;
    END
  END la_iena[121]
  PIN la_iena[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1852.970 736.000 1853.250 740.000 ;
    END
  END la_iena[122]
  PIN la_iena[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1868.150 736.000 1868.430 740.000 ;
    END
  END la_iena[123]
  PIN la_iena[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1883.330 736.000 1883.610 740.000 ;
    END
  END la_iena[124]
  PIN la_iena[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1898.510 736.000 1898.790 740.000 ;
    END
  END la_iena[125]
  PIN la_iena[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1913.690 736.000 1913.970 740.000 ;
    END
  END la_iena[126]
  PIN la_iena[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1928.870 736.000 1929.150 740.000 ;
    END
  END la_iena[127]
  PIN la_iena[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 736.000 183.910 740.000 ;
    END
  END la_iena[12]
  PIN la_iena[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 736.000 199.090 740.000 ;
    END
  END la_iena[13]
  PIN la_iena[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 736.000 214.270 740.000 ;
    END
  END la_iena[14]
  PIN la_iena[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 736.000 229.450 740.000 ;
    END
  END la_iena[15]
  PIN la_iena[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 736.000 244.630 740.000 ;
    END
  END la_iena[16]
  PIN la_iena[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 736.000 259.810 740.000 ;
    END
  END la_iena[17]
  PIN la_iena[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 736.000 274.990 740.000 ;
    END
  END la_iena[18]
  PIN la_iena[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 736.000 290.170 740.000 ;
    END
  END la_iena[19]
  PIN la_iena[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 736.000 16.930 740.000 ;
    END
  END la_iena[1]
  PIN la_iena[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 736.000 305.350 740.000 ;
    END
  END la_iena[20]
  PIN la_iena[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.250 736.000 320.530 740.000 ;
    END
  END la_iena[21]
  PIN la_iena[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 736.000 335.710 740.000 ;
    END
  END la_iena[22]
  PIN la_iena[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.610 736.000 350.890 740.000 ;
    END
  END la_iena[23]
  PIN la_iena[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 736.000 366.070 740.000 ;
    END
  END la_iena[24]
  PIN la_iena[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.970 736.000 381.250 740.000 ;
    END
  END la_iena[25]
  PIN la_iena[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 736.000 396.430 740.000 ;
    END
  END la_iena[26]
  PIN la_iena[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.330 736.000 411.610 740.000 ;
    END
  END la_iena[27]
  PIN la_iena[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.510 736.000 426.790 740.000 ;
    END
  END la_iena[28]
  PIN la_iena[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 736.000 441.970 740.000 ;
    END
  END la_iena[29]
  PIN la_iena[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 736.000 32.110 740.000 ;
    END
  END la_iena[2]
  PIN la_iena[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.870 736.000 457.150 740.000 ;
    END
  END la_iena[30]
  PIN la_iena[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.050 736.000 472.330 740.000 ;
    END
  END la_iena[31]
  PIN la_iena[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.230 736.000 487.510 740.000 ;
    END
  END la_iena[32]
  PIN la_iena[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 736.000 502.690 740.000 ;
    END
  END la_iena[33]
  PIN la_iena[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.590 736.000 517.870 740.000 ;
    END
  END la_iena[34]
  PIN la_iena[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.770 736.000 533.050 740.000 ;
    END
  END la_iena[35]
  PIN la_iena[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.950 736.000 548.230 740.000 ;
    END
  END la_iena[36]
  PIN la_iena[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.130 736.000 563.410 740.000 ;
    END
  END la_iena[37]
  PIN la_iena[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.310 736.000 578.590 740.000 ;
    END
  END la_iena[38]
  PIN la_iena[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.490 736.000 593.770 740.000 ;
    END
  END la_iena[39]
  PIN la_iena[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 736.000 47.290 740.000 ;
    END
  END la_iena[3]
  PIN la_iena[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 736.000 608.950 740.000 ;
    END
  END la_iena[40]
  PIN la_iena[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.850 736.000 624.130 740.000 ;
    END
  END la_iena[41]
  PIN la_iena[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.030 736.000 639.310 740.000 ;
    END
  END la_iena[42]
  PIN la_iena[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.210 736.000 654.490 740.000 ;
    END
  END la_iena[43]
  PIN la_iena[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.390 736.000 669.670 740.000 ;
    END
  END la_iena[44]
  PIN la_iena[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.570 736.000 684.850 740.000 ;
    END
  END la_iena[45]
  PIN la_iena[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.750 736.000 700.030 740.000 ;
    END
  END la_iena[46]
  PIN la_iena[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 736.000 715.210 740.000 ;
    END
  END la_iena[47]
  PIN la_iena[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.110 736.000 730.390 740.000 ;
    END
  END la_iena[48]
  PIN la_iena[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.290 736.000 745.570 740.000 ;
    END
  END la_iena[49]
  PIN la_iena[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 736.000 62.470 740.000 ;
    END
  END la_iena[4]
  PIN la_iena[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.470 736.000 760.750 740.000 ;
    END
  END la_iena[50]
  PIN la_iena[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.650 736.000 775.930 740.000 ;
    END
  END la_iena[51]
  PIN la_iena[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.830 736.000 791.110 740.000 ;
    END
  END la_iena[52]
  PIN la_iena[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.010 736.000 806.290 740.000 ;
    END
  END la_iena[53]
  PIN la_iena[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.190 736.000 821.470 740.000 ;
    END
  END la_iena[54]
  PIN la_iena[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 836.370 736.000 836.650 740.000 ;
    END
  END la_iena[55]
  PIN la_iena[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.550 736.000 851.830 740.000 ;
    END
  END la_iena[56]
  PIN la_iena[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.730 736.000 867.010 740.000 ;
    END
  END la_iena[57]
  PIN la_iena[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.910 736.000 882.190 740.000 ;
    END
  END la_iena[58]
  PIN la_iena[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.090 736.000 897.370 740.000 ;
    END
  END la_iena[59]
  PIN la_iena[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 736.000 77.650 740.000 ;
    END
  END la_iena[5]
  PIN la_iena[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.270 736.000 912.550 740.000 ;
    END
  END la_iena[60]
  PIN la_iena[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 736.000 927.730 740.000 ;
    END
  END la_iena[61]
  PIN la_iena[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.630 736.000 942.910 740.000 ;
    END
  END la_iena[62]
  PIN la_iena[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.810 736.000 958.090 740.000 ;
    END
  END la_iena[63]
  PIN la_iena[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.990 736.000 973.270 740.000 ;
    END
  END la_iena[64]
  PIN la_iena[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.170 736.000 988.450 740.000 ;
    END
  END la_iena[65]
  PIN la_iena[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1003.350 736.000 1003.630 740.000 ;
    END
  END la_iena[66]
  PIN la_iena[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.530 736.000 1018.810 740.000 ;
    END
  END la_iena[67]
  PIN la_iena[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.710 736.000 1033.990 740.000 ;
    END
  END la_iena[68]
  PIN la_iena[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.890 736.000 1049.170 740.000 ;
    END
  END la_iena[69]
  PIN la_iena[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 736.000 92.830 740.000 ;
    END
  END la_iena[6]
  PIN la_iena[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1064.070 736.000 1064.350 740.000 ;
    END
  END la_iena[70]
  PIN la_iena[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.250 736.000 1079.530 740.000 ;
    END
  END la_iena[71]
  PIN la_iena[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.430 736.000 1094.710 740.000 ;
    END
  END la_iena[72]
  PIN la_iena[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1109.610 736.000 1109.890 740.000 ;
    END
  END la_iena[73]
  PIN la_iena[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1124.790 736.000 1125.070 740.000 ;
    END
  END la_iena[74]
  PIN la_iena[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.970 736.000 1140.250 740.000 ;
    END
  END la_iena[75]
  PIN la_iena[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1155.150 736.000 1155.430 740.000 ;
    END
  END la_iena[76]
  PIN la_iena[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1170.330 736.000 1170.610 740.000 ;
    END
  END la_iena[77]
  PIN la_iena[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.510 736.000 1185.790 740.000 ;
    END
  END la_iena[78]
  PIN la_iena[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1200.690 736.000 1200.970 740.000 ;
    END
  END la_iena[79]
  PIN la_iena[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 736.000 108.010 740.000 ;
    END
  END la_iena[7]
  PIN la_iena[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1215.870 736.000 1216.150 740.000 ;
    END
  END la_iena[80]
  PIN la_iena[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.050 736.000 1231.330 740.000 ;
    END
  END la_iena[81]
  PIN la_iena[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1246.230 736.000 1246.510 740.000 ;
    END
  END la_iena[82]
  PIN la_iena[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1261.410 736.000 1261.690 740.000 ;
    END
  END la_iena[83]
  PIN la_iena[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1276.590 736.000 1276.870 740.000 ;
    END
  END la_iena[84]
  PIN la_iena[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.770 736.000 1292.050 740.000 ;
    END
  END la_iena[85]
  PIN la_iena[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1306.950 736.000 1307.230 740.000 ;
    END
  END la_iena[86]
  PIN la_iena[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1322.130 736.000 1322.410 740.000 ;
    END
  END la_iena[87]
  PIN la_iena[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1337.310 736.000 1337.590 740.000 ;
    END
  END la_iena[88]
  PIN la_iena[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.490 736.000 1352.770 740.000 ;
    END
  END la_iena[89]
  PIN la_iena[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 736.000 123.190 740.000 ;
    END
  END la_iena[8]
  PIN la_iena[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1367.670 736.000 1367.950 740.000 ;
    END
  END la_iena[90]
  PIN la_iena[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1382.850 736.000 1383.130 740.000 ;
    END
  END la_iena[91]
  PIN la_iena[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1398.030 736.000 1398.310 740.000 ;
    END
  END la_iena[92]
  PIN la_iena[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1413.210 736.000 1413.490 740.000 ;
    END
  END la_iena[93]
  PIN la_iena[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1428.390 736.000 1428.670 740.000 ;
    END
  END la_iena[94]
  PIN la_iena[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1443.570 736.000 1443.850 740.000 ;
    END
  END la_iena[95]
  PIN la_iena[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1458.750 736.000 1459.030 740.000 ;
    END
  END la_iena[96]
  PIN la_iena[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1473.930 736.000 1474.210 740.000 ;
    END
  END la_iena[97]
  PIN la_iena[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1489.110 736.000 1489.390 740.000 ;
    END
  END la_iena[98]
  PIN la_iena[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1504.290 736.000 1504.570 740.000 ;
    END
  END la_iena[99]
  PIN la_iena[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 736.000 138.370 740.000 ;
    END
  END la_iena[9]
  PIN la_input[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 736.000 5.890 740.000 ;
    END
  END la_input[0]
  PIN la_input[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1523.150 736.000 1523.430 740.000 ;
    END
  END la_input[100]
  PIN la_input[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1538.330 736.000 1538.610 740.000 ;
    END
  END la_input[101]
  PIN la_input[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1553.510 736.000 1553.790 740.000 ;
    END
  END la_input[102]
  PIN la_input[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1568.690 736.000 1568.970 740.000 ;
    END
  END la_input[103]
  PIN la_input[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1583.870 736.000 1584.150 740.000 ;
    END
  END la_input[104]
  PIN la_input[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1599.050 736.000 1599.330 740.000 ;
    END
  END la_input[105]
  PIN la_input[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1614.230 736.000 1614.510 740.000 ;
    END
  END la_input[106]
  PIN la_input[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1629.410 736.000 1629.690 740.000 ;
    END
  END la_input[107]
  PIN la_input[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1644.590 736.000 1644.870 740.000 ;
    END
  END la_input[108]
  PIN la_input[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1659.770 736.000 1660.050 740.000 ;
    END
  END la_input[109]
  PIN la_input[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 736.000 157.690 740.000 ;
    END
  END la_input[10]
  PIN la_input[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1674.950 736.000 1675.230 740.000 ;
    END
  END la_input[110]
  PIN la_input[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1690.130 736.000 1690.410 740.000 ;
    END
  END la_input[111]
  PIN la_input[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1705.310 736.000 1705.590 740.000 ;
    END
  END la_input[112]
  PIN la_input[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1720.490 736.000 1720.770 740.000 ;
    END
  END la_input[113]
  PIN la_input[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1735.670 736.000 1735.950 740.000 ;
    END
  END la_input[114]
  PIN la_input[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1750.850 736.000 1751.130 740.000 ;
    END
  END la_input[115]
  PIN la_input[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1766.030 736.000 1766.310 740.000 ;
    END
  END la_input[116]
  PIN la_input[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1781.210 736.000 1781.490 740.000 ;
    END
  END la_input[117]
  PIN la_input[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1796.390 736.000 1796.670 740.000 ;
    END
  END la_input[118]
  PIN la_input[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1811.570 736.000 1811.850 740.000 ;
    END
  END la_input[119]
  PIN la_input[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 736.000 172.870 740.000 ;
    END
  END la_input[11]
  PIN la_input[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1826.750 736.000 1827.030 740.000 ;
    END
  END la_input[120]
  PIN la_input[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1841.930 736.000 1842.210 740.000 ;
    END
  END la_input[121]
  PIN la_input[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1857.110 736.000 1857.390 740.000 ;
    END
  END la_input[122]
  PIN la_input[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1872.290 736.000 1872.570 740.000 ;
    END
  END la_input[123]
  PIN la_input[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1887.470 736.000 1887.750 740.000 ;
    END
  END la_input[124]
  PIN la_input[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1902.650 736.000 1902.930 740.000 ;
    END
  END la_input[125]
  PIN la_input[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1917.830 736.000 1918.110 740.000 ;
    END
  END la_input[126]
  PIN la_input[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1933.010 736.000 1933.290 740.000 ;
    END
  END la_input[127]
  PIN la_input[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 736.000 188.050 740.000 ;
    END
  END la_input[12]
  PIN la_input[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 736.000 203.230 740.000 ;
    END
  END la_input[13]
  PIN la_input[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 736.000 218.410 740.000 ;
    END
  END la_input[14]
  PIN la_input[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 736.000 233.590 740.000 ;
    END
  END la_input[15]
  PIN la_input[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 736.000 248.770 740.000 ;
    END
  END la_input[16]
  PIN la_input[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 736.000 263.950 740.000 ;
    END
  END la_input[17]
  PIN la_input[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.850 736.000 279.130 740.000 ;
    END
  END la_input[18]
  PIN la_input[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 736.000 294.310 740.000 ;
    END
  END la_input[19]
  PIN la_input[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 736.000 21.070 740.000 ;
    END
  END la_input[1]
  PIN la_input[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 736.000 309.490 740.000 ;
    END
  END la_input[20]
  PIN la_input[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.390 736.000 324.670 740.000 ;
    END
  END la_input[21]
  PIN la_input[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 736.000 339.850 740.000 ;
    END
  END la_input[22]
  PIN la_input[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 736.000 355.030 740.000 ;
    END
  END la_input[23]
  PIN la_input[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.930 736.000 370.210 740.000 ;
    END
  END la_input[24]
  PIN la_input[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 736.000 385.390 740.000 ;
    END
  END la_input[25]
  PIN la_input[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.290 736.000 400.570 740.000 ;
    END
  END la_input[26]
  PIN la_input[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 736.000 415.750 740.000 ;
    END
  END la_input[27]
  PIN la_input[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.650 736.000 430.930 740.000 ;
    END
  END la_input[28]
  PIN la_input[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.830 736.000 446.110 740.000 ;
    END
  END la_input[29]
  PIN la_input[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 736.000 36.250 740.000 ;
    END
  END la_input[2]
  PIN la_input[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 736.000 460.830 740.000 ;
    END
  END la_input[30]
  PIN la_input[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.730 736.000 476.010 740.000 ;
    END
  END la_input[31]
  PIN la_input[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.910 736.000 491.190 740.000 ;
    END
  END la_input[32]
  PIN la_input[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.090 736.000 506.370 740.000 ;
    END
  END la_input[33]
  PIN la_input[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.270 736.000 521.550 740.000 ;
    END
  END la_input[34]
  PIN la_input[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.450 736.000 536.730 740.000 ;
    END
  END la_input[35]
  PIN la_input[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.630 736.000 551.910 740.000 ;
    END
  END la_input[36]
  PIN la_input[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 736.000 567.090 740.000 ;
    END
  END la_input[37]
  PIN la_input[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.990 736.000 582.270 740.000 ;
    END
  END la_input[38]
  PIN la_input[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.170 736.000 597.450 740.000 ;
    END
  END la_input[39]
  PIN la_input[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 736.000 51.430 740.000 ;
    END
  END la_input[3]
  PIN la_input[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.350 736.000 612.630 740.000 ;
    END
  END la_input[40]
  PIN la_input[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.530 736.000 627.810 740.000 ;
    END
  END la_input[41]
  PIN la_input[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.710 736.000 642.990 740.000 ;
    END
  END la_input[42]
  PIN la_input[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.890 736.000 658.170 740.000 ;
    END
  END la_input[43]
  PIN la_input[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.070 736.000 673.350 740.000 ;
    END
  END la_input[44]
  PIN la_input[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.250 736.000 688.530 740.000 ;
    END
  END la_input[45]
  PIN la_input[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.430 736.000 703.710 740.000 ;
    END
  END la_input[46]
  PIN la_input[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.610 736.000 718.890 740.000 ;
    END
  END la_input[47]
  PIN la_input[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.790 736.000 734.070 740.000 ;
    END
  END la_input[48]
  PIN la_input[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.970 736.000 749.250 740.000 ;
    END
  END la_input[49]
  PIN la_input[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 736.000 66.610 740.000 ;
    END
  END la_input[4]
  PIN la_input[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.150 736.000 764.430 740.000 ;
    END
  END la_input[50]
  PIN la_input[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 736.000 779.610 740.000 ;
    END
  END la_input[51]
  PIN la_input[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.510 736.000 794.790 740.000 ;
    END
  END la_input[52]
  PIN la_input[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.690 736.000 809.970 740.000 ;
    END
  END la_input[53]
  PIN la_input[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.870 736.000 825.150 740.000 ;
    END
  END la_input[54]
  PIN la_input[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.050 736.000 840.330 740.000 ;
    END
  END la_input[55]
  PIN la_input[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.230 736.000 855.510 740.000 ;
    END
  END la_input[56]
  PIN la_input[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.410 736.000 870.690 740.000 ;
    END
  END la_input[57]
  PIN la_input[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.590 736.000 885.870 740.000 ;
    END
  END la_input[58]
  PIN la_input[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.770 736.000 901.050 740.000 ;
    END
  END la_input[59]
  PIN la_input[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 736.000 81.790 740.000 ;
    END
  END la_input[5]
  PIN la_input[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.950 736.000 916.230 740.000 ;
    END
  END la_input[60]
  PIN la_input[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.130 736.000 931.410 740.000 ;
    END
  END la_input[61]
  PIN la_input[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.310 736.000 946.590 740.000 ;
    END
  END la_input[62]
  PIN la_input[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.490 736.000 961.770 740.000 ;
    END
  END la_input[63]
  PIN la_input[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.670 736.000 976.950 740.000 ;
    END
  END la_input[64]
  PIN la_input[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.850 736.000 992.130 740.000 ;
    END
  END la_input[65]
  PIN la_input[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.030 736.000 1007.310 740.000 ;
    END
  END la_input[66]
  PIN la_input[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1022.210 736.000 1022.490 740.000 ;
    END
  END la_input[67]
  PIN la_input[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.390 736.000 1037.670 740.000 ;
    END
  END la_input[68]
  PIN la_input[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1052.570 736.000 1052.850 740.000 ;
    END
  END la_input[69]
  PIN la_input[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 736.000 96.970 740.000 ;
    END
  END la_input[6]
  PIN la_input[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1067.750 736.000 1068.030 740.000 ;
    END
  END la_input[70]
  PIN la_input[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.930 736.000 1083.210 740.000 ;
    END
  END la_input[71]
  PIN la_input[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.110 736.000 1098.390 740.000 ;
    END
  END la_input[72]
  PIN la_input[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1113.290 736.000 1113.570 740.000 ;
    END
  END la_input[73]
  PIN la_input[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.470 736.000 1128.750 740.000 ;
    END
  END la_input[74]
  PIN la_input[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.650 736.000 1143.930 740.000 ;
    END
  END la_input[75]
  PIN la_input[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1158.830 736.000 1159.110 740.000 ;
    END
  END la_input[76]
  PIN la_input[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1174.010 736.000 1174.290 740.000 ;
    END
  END la_input[77]
  PIN la_input[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1189.190 736.000 1189.470 740.000 ;
    END
  END la_input[78]
  PIN la_input[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1204.370 736.000 1204.650 740.000 ;
    END
  END la_input[79]
  PIN la_input[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 736.000 112.150 740.000 ;
    END
  END la_input[7]
  PIN la_input[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1219.550 736.000 1219.830 740.000 ;
    END
  END la_input[80]
  PIN la_input[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1234.730 736.000 1235.010 740.000 ;
    END
  END la_input[81]
  PIN la_input[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.910 736.000 1250.190 740.000 ;
    END
  END la_input[82]
  PIN la_input[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1265.090 736.000 1265.370 740.000 ;
    END
  END la_input[83]
  PIN la_input[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1280.270 736.000 1280.550 740.000 ;
    END
  END la_input[84]
  PIN la_input[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1295.450 736.000 1295.730 740.000 ;
    END
  END la_input[85]
  PIN la_input[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1310.630 736.000 1310.910 740.000 ;
    END
  END la_input[86]
  PIN la_input[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1325.810 736.000 1326.090 740.000 ;
    END
  END la_input[87]
  PIN la_input[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.990 736.000 1341.270 740.000 ;
    END
  END la_input[88]
  PIN la_input[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.170 736.000 1356.450 740.000 ;
    END
  END la_input[89]
  PIN la_input[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 736.000 127.330 740.000 ;
    END
  END la_input[8]
  PIN la_input[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1371.350 736.000 1371.630 740.000 ;
    END
  END la_input[90]
  PIN la_input[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1386.530 736.000 1386.810 740.000 ;
    END
  END la_input[91]
  PIN la_input[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1401.710 736.000 1401.990 740.000 ;
    END
  END la_input[92]
  PIN la_input[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1416.890 736.000 1417.170 740.000 ;
    END
  END la_input[93]
  PIN la_input[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.070 736.000 1432.350 740.000 ;
    END
  END la_input[94]
  PIN la_input[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1447.250 736.000 1447.530 740.000 ;
    END
  END la_input[95]
  PIN la_input[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.430 736.000 1462.710 740.000 ;
    END
  END la_input[96]
  PIN la_input[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1477.610 736.000 1477.890 740.000 ;
    END
  END la_input[97]
  PIN la_input[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1492.790 736.000 1493.070 740.000 ;
    END
  END la_input[98]
  PIN la_input[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1507.970 736.000 1508.250 740.000 ;
    END
  END la_input[99]
  PIN la_input[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 736.000 142.510 740.000 ;
    END
  END la_input[9]
  PIN la_oenb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 736.000 9.570 740.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1526.830 736.000 1527.110 740.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.010 736.000 1542.290 740.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1557.190 736.000 1557.470 740.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1572.370 736.000 1572.650 740.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1587.550 736.000 1587.830 740.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1602.730 736.000 1603.010 740.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1617.910 736.000 1618.190 740.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1633.090 736.000 1633.370 740.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1648.270 736.000 1648.550 740.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1663.450 736.000 1663.730 740.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 736.000 161.370 740.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1678.630 736.000 1678.910 740.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.810 736.000 1694.090 740.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1708.990 736.000 1709.270 740.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1724.170 736.000 1724.450 740.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1739.350 736.000 1739.630 740.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1754.530 736.000 1754.810 740.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1769.710 736.000 1769.990 740.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1784.890 736.000 1785.170 740.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1800.070 736.000 1800.350 740.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1815.250 736.000 1815.530 740.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 736.000 176.550 740.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1830.430 736.000 1830.710 740.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1845.610 736.000 1845.890 740.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1860.790 736.000 1861.070 740.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1875.970 736.000 1876.250 740.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1891.150 736.000 1891.430 740.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1906.330 736.000 1906.610 740.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1921.510 736.000 1921.790 740.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1936.690 736.000 1936.970 740.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 736.000 191.730 740.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.630 736.000 206.910 740.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 736.000 222.090 740.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 736.000 237.270 740.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 736.000 252.450 740.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 736.000 267.630 740.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 736.000 282.810 740.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.710 736.000 297.990 740.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 736.000 24.750 740.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 736.000 313.170 740.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.070 736.000 328.350 740.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 736.000 343.530 740.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 736.000 358.710 740.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 736.000 373.890 740.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 736.000 389.070 740.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 736.000 404.250 740.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.150 736.000 419.430 740.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.330 736.000 434.610 740.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 736.000 449.790 740.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 736.000 39.930 740.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.690 736.000 464.970 740.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 736.000 480.150 740.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.050 736.000 495.330 740.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.230 736.000 510.510 740.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.410 736.000 525.690 740.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.590 736.000 540.870 740.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.770 736.000 556.050 740.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.950 736.000 571.230 740.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 736.000 586.410 740.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.310 736.000 601.590 740.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 736.000 55.110 740.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.490 736.000 616.770 740.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.670 736.000 631.950 740.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.850 736.000 647.130 740.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.030 736.000 662.310 740.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.210 736.000 677.490 740.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 736.000 692.670 740.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.570 736.000 707.850 740.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.750 736.000 723.030 740.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.930 736.000 738.210 740.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.110 736.000 753.390 740.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 736.000 70.290 740.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.290 736.000 768.570 740.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.470 736.000 783.750 740.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.650 736.000 798.930 740.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.830 736.000 814.110 740.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.010 736.000 829.290 740.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.190 736.000 844.470 740.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.370 736.000 859.650 740.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 874.550 736.000 874.830 740.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.730 736.000 890.010 740.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.450 736.000 904.730 740.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 736.000 85.470 740.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 919.630 736.000 919.910 740.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 934.810 736.000 935.090 740.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.990 736.000 950.270 740.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.170 736.000 965.450 740.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 980.350 736.000 980.630 740.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.530 736.000 995.810 740.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1010.710 736.000 1010.990 740.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.890 736.000 1026.170 740.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1041.070 736.000 1041.350 740.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.250 736.000 1056.530 740.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 736.000 100.650 740.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1071.430 736.000 1071.710 740.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1086.610 736.000 1086.890 740.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1101.790 736.000 1102.070 740.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1116.970 736.000 1117.250 740.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1132.150 736.000 1132.430 740.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1147.330 736.000 1147.610 740.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.510 736.000 1162.790 740.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1177.690 736.000 1177.970 740.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1192.870 736.000 1193.150 740.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.050 736.000 1208.330 740.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 736.000 115.830 740.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1223.230 736.000 1223.510 740.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1238.410 736.000 1238.690 740.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1253.590 736.000 1253.870 740.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1268.770 736.000 1269.050 740.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1283.950 736.000 1284.230 740.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1299.130 736.000 1299.410 740.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1314.310 736.000 1314.590 740.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1329.490 736.000 1329.770 740.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.670 736.000 1344.950 740.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1359.850 736.000 1360.130 740.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 736.000 131.010 740.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.030 736.000 1375.310 740.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1390.210 736.000 1390.490 740.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1405.390 736.000 1405.670 740.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1420.570 736.000 1420.850 740.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1435.750 736.000 1436.030 740.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1450.930 736.000 1451.210 740.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1466.110 736.000 1466.390 740.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1481.290 736.000 1481.570 740.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1496.470 736.000 1496.750 740.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1511.650 736.000 1511.930 740.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 736.000 146.190 740.000 ;
    END
  END la_oenb[9]
  PIN la_output[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 736.000 13.250 740.000 ;
    END
  END la_output[0]
  PIN la_output[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1530.510 736.000 1530.790 740.000 ;
    END
  END la_output[100]
  PIN la_output[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.690 736.000 1545.970 740.000 ;
    END
  END la_output[101]
  PIN la_output[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1560.870 736.000 1561.150 740.000 ;
    END
  END la_output[102]
  PIN la_output[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1576.050 736.000 1576.330 740.000 ;
    END
  END la_output[103]
  PIN la_output[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1591.230 736.000 1591.510 740.000 ;
    END
  END la_output[104]
  PIN la_output[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1606.410 736.000 1606.690 740.000 ;
    END
  END la_output[105]
  PIN la_output[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1621.590 736.000 1621.870 740.000 ;
    END
  END la_output[106]
  PIN la_output[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1636.770 736.000 1637.050 740.000 ;
    END
  END la_output[107]
  PIN la_output[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.950 736.000 1652.230 740.000 ;
    END
  END la_output[108]
  PIN la_output[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1667.130 736.000 1667.410 740.000 ;
    END
  END la_output[109]
  PIN la_output[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 736.000 165.050 740.000 ;
    END
  END la_output[10]
  PIN la_output[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1682.310 736.000 1682.590 740.000 ;
    END
  END la_output[110]
  PIN la_output[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1697.490 736.000 1697.770 740.000 ;
    END
  END la_output[111]
  PIN la_output[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1712.670 736.000 1712.950 740.000 ;
    END
  END la_output[112]
  PIN la_output[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1727.850 736.000 1728.130 740.000 ;
    END
  END la_output[113]
  PIN la_output[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.030 736.000 1743.310 740.000 ;
    END
  END la_output[114]
  PIN la_output[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.210 736.000 1758.490 740.000 ;
    END
  END la_output[115]
  PIN la_output[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1773.390 736.000 1773.670 740.000 ;
    END
  END la_output[116]
  PIN la_output[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1788.570 736.000 1788.850 740.000 ;
    END
  END la_output[117]
  PIN la_output[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1803.750 736.000 1804.030 740.000 ;
    END
  END la_output[118]
  PIN la_output[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1818.930 736.000 1819.210 740.000 ;
    END
  END la_output[119]
  PIN la_output[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 736.000 180.230 740.000 ;
    END
  END la_output[11]
  PIN la_output[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1834.110 736.000 1834.390 740.000 ;
    END
  END la_output[120]
  PIN la_output[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1849.290 736.000 1849.570 740.000 ;
    END
  END la_output[121]
  PIN la_output[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1864.470 736.000 1864.750 740.000 ;
    END
  END la_output[122]
  PIN la_output[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1879.650 736.000 1879.930 740.000 ;
    END
  END la_output[123]
  PIN la_output[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1894.830 736.000 1895.110 740.000 ;
    END
  END la_output[124]
  PIN la_output[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1910.010 736.000 1910.290 740.000 ;
    END
  END la_output[125]
  PIN la_output[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1925.190 736.000 1925.470 740.000 ;
    END
  END la_output[126]
  PIN la_output[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1940.370 736.000 1940.650 740.000 ;
    END
  END la_output[127]
  PIN la_output[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 736.000 195.410 740.000 ;
    END
  END la_output[12]
  PIN la_output[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.310 736.000 210.590 740.000 ;
    END
  END la_output[13]
  PIN la_output[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 736.000 225.770 740.000 ;
    END
  END la_output[14]
  PIN la_output[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 736.000 240.950 740.000 ;
    END
  END la_output[15]
  PIN la_output[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 736.000 256.130 740.000 ;
    END
  END la_output[16]
  PIN la_output[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 736.000 271.310 740.000 ;
    END
  END la_output[17]
  PIN la_output[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 736.000 286.490 740.000 ;
    END
  END la_output[18]
  PIN la_output[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 736.000 301.670 740.000 ;
    END
  END la_output[19]
  PIN la_output[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 736.000 28.430 740.000 ;
    END
  END la_output[1]
  PIN la_output[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 736.000 316.850 740.000 ;
    END
  END la_output[20]
  PIN la_output[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 736.000 332.030 740.000 ;
    END
  END la_output[21]
  PIN la_output[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.930 736.000 347.210 740.000 ;
    END
  END la_output[22]
  PIN la_output[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 736.000 362.390 740.000 ;
    END
  END la_output[23]
  PIN la_output[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 736.000 377.570 740.000 ;
    END
  END la_output[24]
  PIN la_output[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.470 736.000 392.750 740.000 ;
    END
  END la_output[25]
  PIN la_output[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.650 736.000 407.930 740.000 ;
    END
  END la_output[26]
  PIN la_output[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.830 736.000 423.110 740.000 ;
    END
  END la_output[27]
  PIN la_output[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 736.000 438.290 740.000 ;
    END
  END la_output[28]
  PIN la_output[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.190 736.000 453.470 740.000 ;
    END
  END la_output[29]
  PIN la_output[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 736.000 43.610 740.000 ;
    END
  END la_output[2]
  PIN la_output[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.370 736.000 468.650 740.000 ;
    END
  END la_output[30]
  PIN la_output[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.550 736.000 483.830 740.000 ;
    END
  END la_output[31]
  PIN la_output[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.730 736.000 499.010 740.000 ;
    END
  END la_output[32]
  PIN la_output[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.910 736.000 514.190 740.000 ;
    END
  END la_output[33]
  PIN la_output[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.090 736.000 529.370 740.000 ;
    END
  END la_output[34]
  PIN la_output[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 736.000 544.550 740.000 ;
    END
  END la_output[35]
  PIN la_output[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.450 736.000 559.730 740.000 ;
    END
  END la_output[36]
  PIN la_output[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.630 736.000 574.910 740.000 ;
    END
  END la_output[37]
  PIN la_output[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.810 736.000 590.090 740.000 ;
    END
  END la_output[38]
  PIN la_output[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.990 736.000 605.270 740.000 ;
    END
  END la_output[39]
  PIN la_output[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 736.000 58.790 740.000 ;
    END
  END la_output[3]
  PIN la_output[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.170 736.000 620.450 740.000 ;
    END
  END la_output[40]
  PIN la_output[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.350 736.000 635.630 740.000 ;
    END
  END la_output[41]
  PIN la_output[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 736.000 650.810 740.000 ;
    END
  END la_output[42]
  PIN la_output[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.710 736.000 665.990 740.000 ;
    END
  END la_output[43]
  PIN la_output[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.890 736.000 681.170 740.000 ;
    END
  END la_output[44]
  PIN la_output[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.070 736.000 696.350 740.000 ;
    END
  END la_output[45]
  PIN la_output[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.250 736.000 711.530 740.000 ;
    END
  END la_output[46]
  PIN la_output[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.430 736.000 726.710 740.000 ;
    END
  END la_output[47]
  PIN la_output[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.610 736.000 741.890 740.000 ;
    END
  END la_output[48]
  PIN la_output[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 736.000 757.070 740.000 ;
    END
  END la_output[49]
  PIN la_output[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 736.000 73.970 740.000 ;
    END
  END la_output[4]
  PIN la_output[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.970 736.000 772.250 740.000 ;
    END
  END la_output[50]
  PIN la_output[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.150 736.000 787.430 740.000 ;
    END
  END la_output[51]
  PIN la_output[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.330 736.000 802.610 740.000 ;
    END
  END la_output[52]
  PIN la_output[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.510 736.000 817.790 740.000 ;
    END
  END la_output[53]
  PIN la_output[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.690 736.000 832.970 740.000 ;
    END
  END la_output[54]
  PIN la_output[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.870 736.000 848.150 740.000 ;
    END
  END la_output[55]
  PIN la_output[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.050 736.000 863.330 740.000 ;
    END
  END la_output[56]
  PIN la_output[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 878.230 736.000 878.510 740.000 ;
    END
  END la_output[57]
  PIN la_output[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.410 736.000 893.690 740.000 ;
    END
  END la_output[58]
  PIN la_output[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.590 736.000 908.870 740.000 ;
    END
  END la_output[59]
  PIN la_output[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 736.000 89.150 740.000 ;
    END
  END la_output[5]
  PIN la_output[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 923.770 736.000 924.050 740.000 ;
    END
  END la_output[60]
  PIN la_output[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.950 736.000 939.230 740.000 ;
    END
  END la_output[61]
  PIN la_output[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 954.130 736.000 954.410 740.000 ;
    END
  END la_output[62]
  PIN la_output[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.310 736.000 969.590 740.000 ;
    END
  END la_output[63]
  PIN la_output[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.490 736.000 984.770 740.000 ;
    END
  END la_output[64]
  PIN la_output[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 999.670 736.000 999.950 740.000 ;
    END
  END la_output[65]
  PIN la_output[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.850 736.000 1015.130 740.000 ;
    END
  END la_output[66]
  PIN la_output[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.030 736.000 1030.310 740.000 ;
    END
  END la_output[67]
  PIN la_output[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1045.210 736.000 1045.490 740.000 ;
    END
  END la_output[68]
  PIN la_output[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1060.390 736.000 1060.670 740.000 ;
    END
  END la_output[69]
  PIN la_output[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 736.000 104.330 740.000 ;
    END
  END la_output[6]
  PIN la_output[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1075.570 736.000 1075.850 740.000 ;
    END
  END la_output[70]
  PIN la_output[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.750 736.000 1091.030 740.000 ;
    END
  END la_output[71]
  PIN la_output[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1105.930 736.000 1106.210 740.000 ;
    END
  END la_output[72]
  PIN la_output[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1121.110 736.000 1121.390 740.000 ;
    END
  END la_output[73]
  PIN la_output[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.290 736.000 1136.570 740.000 ;
    END
  END la_output[74]
  PIN la_output[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1151.470 736.000 1151.750 740.000 ;
    END
  END la_output[75]
  PIN la_output[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1166.650 736.000 1166.930 740.000 ;
    END
  END la_output[76]
  PIN la_output[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1181.830 736.000 1182.110 740.000 ;
    END
  END la_output[77]
  PIN la_output[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.010 736.000 1197.290 740.000 ;
    END
  END la_output[78]
  PIN la_output[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1212.190 736.000 1212.470 740.000 ;
    END
  END la_output[79]
  PIN la_output[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 736.000 119.510 740.000 ;
    END
  END la_output[7]
  PIN la_output[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1227.370 736.000 1227.650 740.000 ;
    END
  END la_output[80]
  PIN la_output[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1242.550 736.000 1242.830 740.000 ;
    END
  END la_output[81]
  PIN la_output[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.730 736.000 1258.010 740.000 ;
    END
  END la_output[82]
  PIN la_output[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1272.910 736.000 1273.190 740.000 ;
    END
  END la_output[83]
  PIN la_output[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1288.090 736.000 1288.370 740.000 ;
    END
  END la_output[84]
  PIN la_output[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1303.270 736.000 1303.550 740.000 ;
    END
  END la_output[85]
  PIN la_output[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1318.450 736.000 1318.730 740.000 ;
    END
  END la_output[86]
  PIN la_output[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1333.630 736.000 1333.910 740.000 ;
    END
  END la_output[87]
  PIN la_output[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1348.810 736.000 1349.090 740.000 ;
    END
  END la_output[88]
  PIN la_output[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1363.530 736.000 1363.810 740.000 ;
    END
  END la_output[89]
  PIN la_output[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 736.000 134.690 740.000 ;
    END
  END la_output[8]
  PIN la_output[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1378.710 736.000 1378.990 740.000 ;
    END
  END la_output[90]
  PIN la_output[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1393.890 736.000 1394.170 740.000 ;
    END
  END la_output[91]
  PIN la_output[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1409.070 736.000 1409.350 740.000 ;
    END
  END la_output[92]
  PIN la_output[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1424.250 736.000 1424.530 740.000 ;
    END
  END la_output[93]
  PIN la_output[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.430 736.000 1439.710 740.000 ;
    END
  END la_output[94]
  PIN la_output[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1454.610 736.000 1454.890 740.000 ;
    END
  END la_output[95]
  PIN la_output[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1469.790 736.000 1470.070 740.000 ;
    END
  END la_output[96]
  PIN la_output[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.970 736.000 1485.250 740.000 ;
    END
  END la_output[97]
  PIN la_output[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.150 736.000 1500.430 740.000 ;
    END
  END la_output[98]
  PIN la_output[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1515.330 736.000 1515.610 740.000 ;
    END
  END la_output[99]
  PIN la_output[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 736.000 149.870 740.000 ;
    END
  END la_output[9]
  PIN mem_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.840 4.000 432.440 ;
    END
  END mem_addr[0]
  PIN mem_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 438.640 4.000 439.240 ;
    END
  END mem_addr[1]
  PIN mem_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.760 4.000 445.360 ;
    END
  END mem_addr[2]
  PIN mem_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 451.560 4.000 452.160 ;
    END
  END mem_addr[3]
  PIN mem_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 458.360 4.000 458.960 ;
    END
  END mem_addr[4]
  PIN mem_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.160 4.000 465.760 ;
    END
  END mem_addr[5]
  PIN mem_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.280 4.000 471.880 ;
    END
  END mem_addr[6]
  PIN mem_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.080 4.000 478.680 ;
    END
  END mem_addr[7]
  PIN mem_ena
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END mem_ena
  PIN mem_rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END mem_rdata[0]
  PIN mem_rdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END mem_rdata[10]
  PIN mem_rdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END mem_rdata[11]
  PIN mem_rdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END mem_rdata[12]
  PIN mem_rdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END mem_rdata[13]
  PIN mem_rdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 4.000 101.960 ;
    END
  END mem_rdata[14]
  PIN mem_rdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 4.000 108.760 ;
    END
  END mem_rdata[15]
  PIN mem_rdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.960 4.000 115.560 ;
    END
  END mem_rdata[16]
  PIN mem_rdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END mem_rdata[17]
  PIN mem_rdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END mem_rdata[18]
  PIN mem_rdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END mem_rdata[19]
  PIN mem_rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 4.000 16.280 ;
    END
  END mem_rdata[1]
  PIN mem_rdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END mem_rdata[20]
  PIN mem_rdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 147.600 4.000 148.200 ;
    END
  END mem_rdata[21]
  PIN mem_rdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 154.400 4.000 155.000 ;
    END
  END mem_rdata[22]
  PIN mem_rdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.200 4.000 161.800 ;
    END
  END mem_rdata[23]
  PIN mem_rdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END mem_rdata[24]
  PIN mem_rdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END mem_rdata[25]
  PIN mem_rdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END mem_rdata[26]
  PIN mem_rdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END mem_rdata[27]
  PIN mem_rdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END mem_rdata[28]
  PIN mem_rdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END mem_rdata[29]
  PIN mem_rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 4.000 23.080 ;
    END
  END mem_rdata[2]
  PIN mem_rdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END mem_rdata[30]
  PIN mem_rdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END mem_rdata[31]
  PIN mem_rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END mem_rdata[3]
  PIN mem_rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END mem_rdata[4]
  PIN mem_rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END mem_rdata[5]
  PIN mem_rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END mem_rdata[6]
  PIN mem_rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.120 4.000 55.720 ;
    END
  END mem_rdata[7]
  PIN mem_rdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.920 4.000 62.520 ;
    END
  END mem_rdata[8]
  PIN mem_rdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 4.000 69.320 ;
    END
  END mem_rdata[9]
  PIN mem_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END mem_wdata[0]
  PIN mem_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 286.320 4.000 286.920 ;
    END
  END mem_wdata[10]
  PIN mem_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.120 4.000 293.720 ;
    END
  END mem_wdata[11]
  PIN mem_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.920 4.000 300.520 ;
    END
  END mem_wdata[12]
  PIN mem_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END mem_wdata[13]
  PIN mem_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END mem_wdata[14]
  PIN mem_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END mem_wdata[15]
  PIN mem_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END mem_wdata[16]
  PIN mem_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 332.560 4.000 333.160 ;
    END
  END mem_wdata[17]
  PIN mem_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 339.360 4.000 339.960 ;
    END
  END mem_wdata[18]
  PIN mem_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.160 4.000 346.760 ;
    END
  END mem_wdata[19]
  PIN mem_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END mem_wdata[1]
  PIN mem_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.280 4.000 352.880 ;
    END
  END mem_wdata[20]
  PIN mem_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.080 4.000 359.680 ;
    END
  END mem_wdata[21]
  PIN mem_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 4.000 366.480 ;
    END
  END mem_wdata[22]
  PIN mem_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 4.000 373.280 ;
    END
  END mem_wdata[23]
  PIN mem_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.800 4.000 379.400 ;
    END
  END mem_wdata[24]
  PIN mem_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 385.600 4.000 386.200 ;
    END
  END mem_wdata[25]
  PIN mem_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 392.400 4.000 393.000 ;
    END
  END mem_wdata[26]
  PIN mem_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END mem_wdata[27]
  PIN mem_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 405.320 4.000 405.920 ;
    END
  END mem_wdata[28]
  PIN mem_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.120 4.000 412.720 ;
    END
  END mem_wdata[29]
  PIN mem_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END mem_wdata[2]
  PIN mem_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.920 4.000 419.520 ;
    END
  END mem_wdata[30]
  PIN mem_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.040 4.000 425.640 ;
    END
  END mem_wdata[31]
  PIN mem_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.080 4.000 240.680 ;
    END
  END mem_wdata[3]
  PIN mem_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.880 4.000 247.480 ;
    END
  END mem_wdata[4]
  PIN mem_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.680 4.000 254.280 ;
    END
  END mem_wdata[5]
  PIN mem_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END mem_wdata[6]
  PIN mem_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END mem_wdata[7]
  PIN mem_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END mem_wdata[8]
  PIN mem_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.200 4.000 280.800 ;
    END
  END mem_wdata[9]
  PIN mem_wen[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 484.880 4.000 485.480 ;
    END
  END mem_wen[0]
  PIN mem_wen[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.000 4.000 491.600 ;
    END
  END mem_wen[1]
  PIN mem_wen[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 497.800 4.000 498.400 ;
    END
  END mem_wen[2]
  PIN mem_wen[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 504.600 4.000 505.200 ;
    END
  END mem_wen[3]
  PIN mprj_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 735.800 4.000 736.400 ;
    END
  END mprj_ack_i
  PIN mprj_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1955.550 736.000 1955.830 740.000 ;
    END
  END mprj_adr_o[0]
  PIN mprj_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2046.630 736.000 2046.910 740.000 ;
    END
  END mprj_adr_o[10]
  PIN mprj_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2054.450 736.000 2054.730 740.000 ;
    END
  END mprj_adr_o[11]
  PIN mprj_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2061.810 736.000 2062.090 740.000 ;
    END
  END mprj_adr_o[12]
  PIN mprj_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2069.630 736.000 2069.910 740.000 ;
    END
  END mprj_adr_o[13]
  PIN mprj_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2076.990 736.000 2077.270 740.000 ;
    END
  END mprj_adr_o[14]
  PIN mprj_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2084.810 736.000 2085.090 740.000 ;
    END
  END mprj_adr_o[15]
  PIN mprj_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2092.170 736.000 2092.450 740.000 ;
    END
  END mprj_adr_o[16]
  PIN mprj_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2099.990 736.000 2100.270 740.000 ;
    END
  END mprj_adr_o[17]
  PIN mprj_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2107.350 736.000 2107.630 740.000 ;
    END
  END mprj_adr_o[18]
  PIN mprj_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2115.170 736.000 2115.450 740.000 ;
    END
  END mprj_adr_o[19]
  PIN mprj_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1967.050 736.000 1967.330 740.000 ;
    END
  END mprj_adr_o[1]
  PIN mprj_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2122.530 736.000 2122.810 740.000 ;
    END
  END mprj_adr_o[20]
  PIN mprj_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2130.350 736.000 2130.630 740.000 ;
    END
  END mprj_adr_o[21]
  PIN mprj_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2137.710 736.000 2137.990 740.000 ;
    END
  END mprj_adr_o[22]
  PIN mprj_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2145.530 736.000 2145.810 740.000 ;
    END
  END mprj_adr_o[23]
  PIN mprj_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2152.890 736.000 2153.170 740.000 ;
    END
  END mprj_adr_o[24]
  PIN mprj_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2160.710 736.000 2160.990 740.000 ;
    END
  END mprj_adr_o[25]
  PIN mprj_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2168.070 736.000 2168.350 740.000 ;
    END
  END mprj_adr_o[26]
  PIN mprj_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2175.890 736.000 2176.170 740.000 ;
    END
  END mprj_adr_o[27]
  PIN mprj_adr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2183.250 736.000 2183.530 740.000 ;
    END
  END mprj_adr_o[28]
  PIN mprj_adr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2191.070 736.000 2191.350 740.000 ;
    END
  END mprj_adr_o[29]
  PIN mprj_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1978.550 736.000 1978.830 740.000 ;
    END
  END mprj_adr_o[2]
  PIN mprj_adr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2198.430 736.000 2198.710 740.000 ;
    END
  END mprj_adr_o[30]
  PIN mprj_adr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2206.250 736.000 2206.530 740.000 ;
    END
  END mprj_adr_o[31]
  PIN mprj_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1989.590 736.000 1989.870 740.000 ;
    END
  END mprj_adr_o[3]
  PIN mprj_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2001.090 736.000 2001.370 740.000 ;
    END
  END mprj_adr_o[4]
  PIN mprj_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2008.910 736.000 2009.190 740.000 ;
    END
  END mprj_adr_o[5]
  PIN mprj_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2016.270 736.000 2016.550 740.000 ;
    END
  END mprj_adr_o[6]
  PIN mprj_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2024.090 736.000 2024.370 740.000 ;
    END
  END mprj_adr_o[7]
  PIN mprj_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2031.450 736.000 2031.730 740.000 ;
    END
  END mprj_adr_o[8]
  PIN mprj_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2039.270 736.000 2039.550 740.000 ;
    END
  END mprj_adr_o[9]
  PIN mprj_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1944.050 736.000 1944.330 740.000 ;
    END
  END mprj_cyc_o
  PIN mprj_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 524.320 4.000 524.920 ;
    END
  END mprj_dat_i[0]
  PIN mprj_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.280 4.000 590.880 ;
    END
  END mprj_dat_i[10]
  PIN mprj_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 597.080 4.000 597.680 ;
    END
  END mprj_dat_i[11]
  PIN mprj_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 603.880 4.000 604.480 ;
    END
  END mprj_dat_i[12]
  PIN mprj_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 610.000 4.000 610.600 ;
    END
  END mprj_dat_i[13]
  PIN mprj_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 616.800 4.000 617.400 ;
    END
  END mprj_dat_i[14]
  PIN mprj_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 623.600 4.000 624.200 ;
    END
  END mprj_dat_i[15]
  PIN mprj_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.720 4.000 630.320 ;
    END
  END mprj_dat_i[16]
  PIN mprj_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 636.520 4.000 637.120 ;
    END
  END mprj_dat_i[17]
  PIN mprj_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 643.320 4.000 643.920 ;
    END
  END mprj_dat_i[18]
  PIN mprj_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 650.120 4.000 650.720 ;
    END
  END mprj_dat_i[19]
  PIN mprj_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.120 4.000 531.720 ;
    END
  END mprj_dat_i[1]
  PIN mprj_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 656.240 4.000 656.840 ;
    END
  END mprj_dat_i[20]
  PIN mprj_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.040 4.000 663.640 ;
    END
  END mprj_dat_i[21]
  PIN mprj_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.840 4.000 670.440 ;
    END
  END mprj_dat_i[22]
  PIN mprj_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 675.960 4.000 676.560 ;
    END
  END mprj_dat_i[23]
  PIN mprj_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 682.760 4.000 683.360 ;
    END
  END mprj_dat_i[24]
  PIN mprj_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 689.560 4.000 690.160 ;
    END
  END mprj_dat_i[25]
  PIN mprj_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 696.360 4.000 696.960 ;
    END
  END mprj_dat_i[26]
  PIN mprj_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 702.480 4.000 703.080 ;
    END
  END mprj_dat_i[27]
  PIN mprj_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 709.280 4.000 709.880 ;
    END
  END mprj_dat_i[28]
  PIN mprj_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 716.080 4.000 716.680 ;
    END
  END mprj_dat_i[29]
  PIN mprj_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END mprj_dat_i[2]
  PIN mprj_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 722.200 4.000 722.800 ;
    END
  END mprj_dat_i[30]
  PIN mprj_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 729.000 4.000 729.600 ;
    END
  END mprj_dat_i[31]
  PIN mprj_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.040 4.000 544.640 ;
    END
  END mprj_dat_i[3]
  PIN mprj_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END mprj_dat_i[4]
  PIN mprj_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END mprj_dat_i[5]
  PIN mprj_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 563.760 4.000 564.360 ;
    END
  END mprj_dat_i[6]
  PIN mprj_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 570.560 4.000 571.160 ;
    END
  END mprj_dat_i[7]
  PIN mprj_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 577.360 4.000 577.960 ;
    END
  END mprj_dat_i[8]
  PIN mprj_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 583.480 4.000 584.080 ;
    END
  END mprj_dat_i[9]
  PIN mprj_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1959.230 736.000 1959.510 740.000 ;
    END
  END mprj_dat_o[0]
  PIN mprj_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2050.310 736.000 2050.590 740.000 ;
    END
  END mprj_dat_o[10]
  PIN mprj_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2058.130 736.000 2058.410 740.000 ;
    END
  END mprj_dat_o[11]
  PIN mprj_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2065.490 736.000 2065.770 740.000 ;
    END
  END mprj_dat_o[12]
  PIN mprj_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2073.310 736.000 2073.590 740.000 ;
    END
  END mprj_dat_o[13]
  PIN mprj_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2080.670 736.000 2080.950 740.000 ;
    END
  END mprj_dat_o[14]
  PIN mprj_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2088.490 736.000 2088.770 740.000 ;
    END
  END mprj_dat_o[15]
  PIN mprj_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2095.850 736.000 2096.130 740.000 ;
    END
  END mprj_dat_o[16]
  PIN mprj_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2103.670 736.000 2103.950 740.000 ;
    END
  END mprj_dat_o[17]
  PIN mprj_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2111.030 736.000 2111.310 740.000 ;
    END
  END mprj_dat_o[18]
  PIN mprj_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2118.850 736.000 2119.130 740.000 ;
    END
  END mprj_dat_o[19]
  PIN mprj_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1970.730 736.000 1971.010 740.000 ;
    END
  END mprj_dat_o[1]
  PIN mprj_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2126.210 736.000 2126.490 740.000 ;
    END
  END mprj_dat_o[20]
  PIN mprj_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2134.030 736.000 2134.310 740.000 ;
    END
  END mprj_dat_o[21]
  PIN mprj_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2141.390 736.000 2141.670 740.000 ;
    END
  END mprj_dat_o[22]
  PIN mprj_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2149.210 736.000 2149.490 740.000 ;
    END
  END mprj_dat_o[23]
  PIN mprj_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2156.570 736.000 2156.850 740.000 ;
    END
  END mprj_dat_o[24]
  PIN mprj_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2164.390 736.000 2164.670 740.000 ;
    END
  END mprj_dat_o[25]
  PIN mprj_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2171.750 736.000 2172.030 740.000 ;
    END
  END mprj_dat_o[26]
  PIN mprj_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2179.570 736.000 2179.850 740.000 ;
    END
  END mprj_dat_o[27]
  PIN mprj_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2186.930 736.000 2187.210 740.000 ;
    END
  END mprj_dat_o[28]
  PIN mprj_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2194.750 736.000 2195.030 740.000 ;
    END
  END mprj_dat_o[29]
  PIN mprj_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1982.230 736.000 1982.510 740.000 ;
    END
  END mprj_dat_o[2]
  PIN mprj_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2202.110 736.000 2202.390 740.000 ;
    END
  END mprj_dat_o[30]
  PIN mprj_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2209.930 736.000 2210.210 740.000 ;
    END
  END mprj_dat_o[31]
  PIN mprj_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1993.730 736.000 1994.010 740.000 ;
    END
  END mprj_dat_o[3]
  PIN mprj_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2004.770 736.000 2005.050 740.000 ;
    END
  END mprj_dat_o[4]
  PIN mprj_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2012.590 736.000 2012.870 740.000 ;
    END
  END mprj_dat_o[5]
  PIN mprj_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2019.950 736.000 2020.230 740.000 ;
    END
  END mprj_dat_o[6]
  PIN mprj_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2027.770 736.000 2028.050 740.000 ;
    END
  END mprj_dat_o[7]
  PIN mprj_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2035.130 736.000 2035.410 740.000 ;
    END
  END mprj_dat_o[8]
  PIN mprj_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2042.950 736.000 2043.230 740.000 ;
    END
  END mprj_dat_o[9]
  PIN mprj_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1963.370 736.000 1963.650 740.000 ;
    END
  END mprj_sel_o[0]
  PIN mprj_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1974.410 736.000 1974.690 740.000 ;
    END
  END mprj_sel_o[1]
  PIN mprj_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1985.910 736.000 1986.190 740.000 ;
    END
  END mprj_sel_o[2]
  PIN mprj_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1997.410 736.000 1997.690 740.000 ;
    END
  END mprj_sel_o[3]
  PIN mprj_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1948.190 736.000 1948.470 740.000 ;
    END
  END mprj_stb_o
  PIN mprj_wb_iena
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2213.610 736.000 2213.890 740.000 ;
    END
  END mprj_wb_iena
  PIN mprj_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1951.870 736.000 1952.150 740.000 ;
    END
  END mprj_we_o
  PIN qspi_enabled
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 0.000 447.950 4.000 ;
    END
  END qspi_enabled
  PIN resetn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END resetn
  PIN sdo_oenb_state
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2246.000 554.920 2250.000 555.520 ;
    END
  END sdo_oenb_state
  PIN ser_rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2239.370 0.000 2239.650 4.000 ;
    END
  END ser_rx
  PIN ser_tx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2199.810 0.000 2200.090 4.000 ;
    END
  END ser_tx
  PIN spi_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2060.430 0.000 2060.710 4.000 ;
    END
  END spi_csb
  PIN spi_enabled
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2080.210 0.000 2080.490 4.000 ;
    END
  END spi_enabled
  PIN spi_sck
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2099.990 0.000 2100.270 4.000 ;
    END
  END spi_sck
  PIN spi_sdi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2120.230 0.000 2120.510 4.000 ;
    END
  END spi_sdi
  PIN spi_sdo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2140.010 0.000 2140.290 4.000 ;
    END
  END spi_sdo
  PIN spi_sdoenb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2159.790 0.000 2160.070 4.000 ;
    END
  END spi_sdoenb
  PIN sram_ro_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1184.130 0.000 1184.410 4.000 ;
    END
  END sram_ro_addr[0]
  PIN sram_ro_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1203.910 0.000 1204.190 4.000 ;
    END
  END sram_ro_addr[1]
  PIN sram_ro_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1224.150 0.000 1224.430 4.000 ;
    END
  END sram_ro_addr[2]
  PIN sram_ro_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.930 0.000 1244.210 4.000 ;
    END
  END sram_ro_addr[3]
  PIN sram_ro_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1263.710 0.000 1263.990 4.000 ;
    END
  END sram_ro_addr[4]
  PIN sram_ro_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1283.950 0.000 1284.230 4.000 ;
    END
  END sram_ro_addr[5]
  PIN sram_ro_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1303.730 0.000 1304.010 4.000 ;
    END
  END sram_ro_addr[6]
  PIN sram_ro_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.510 0.000 1323.790 4.000 ;
    END
  END sram_ro_addr[7]
  PIN sram_ro_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1144.570 0.000 1144.850 4.000 ;
    END
  END sram_ro_clk
  PIN sram_ro_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1164.350 0.000 1164.630 4.000 ;
    END
  END sram_ro_csb
  PIN sram_ro_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1343.290 0.000 1343.570 4.000 ;
    END
  END sram_ro_data[0]
  PIN sram_ro_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.470 0.000 1542.750 4.000 ;
    END
  END sram_ro_data[10]
  PIN sram_ro_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1562.710 0.000 1562.990 4.000 ;
    END
  END sram_ro_data[11]
  PIN sram_ro_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1582.490 0.000 1582.770 4.000 ;
    END
  END sram_ro_data[12]
  PIN sram_ro_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1602.270 0.000 1602.550 4.000 ;
    END
  END sram_ro_data[13]
  PIN sram_ro_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1622.050 0.000 1622.330 4.000 ;
    END
  END sram_ro_data[14]
  PIN sram_ro_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1642.290 0.000 1642.570 4.000 ;
    END
  END sram_ro_data[15]
  PIN sram_ro_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1662.070 0.000 1662.350 4.000 ;
    END
  END sram_ro_data[16]
  PIN sram_ro_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1681.850 0.000 1682.130 4.000 ;
    END
  END sram_ro_data[17]
  PIN sram_ro_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1702.090 0.000 1702.370 4.000 ;
    END
  END sram_ro_data[18]
  PIN sram_ro_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1721.870 0.000 1722.150 4.000 ;
    END
  END sram_ro_data[19]
  PIN sram_ro_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1363.530 0.000 1363.810 4.000 ;
    END
  END sram_ro_data[1]
  PIN sram_ro_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1741.650 0.000 1741.930 4.000 ;
    END
  END sram_ro_data[20]
  PIN sram_ro_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1761.430 0.000 1761.710 4.000 ;
    END
  END sram_ro_data[21]
  PIN sram_ro_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1781.670 0.000 1781.950 4.000 ;
    END
  END sram_ro_data[22]
  PIN sram_ro_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1801.450 0.000 1801.730 4.000 ;
    END
  END sram_ro_data[23]
  PIN sram_ro_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1821.230 0.000 1821.510 4.000 ;
    END
  END sram_ro_data[24]
  PIN sram_ro_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1841.470 0.000 1841.750 4.000 ;
    END
  END sram_ro_data[25]
  PIN sram_ro_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1861.250 0.000 1861.530 4.000 ;
    END
  END sram_ro_data[26]
  PIN sram_ro_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1881.030 0.000 1881.310 4.000 ;
    END
  END sram_ro_data[27]
  PIN sram_ro_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1900.810 0.000 1901.090 4.000 ;
    END
  END sram_ro_data[28]
  PIN sram_ro_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1921.050 0.000 1921.330 4.000 ;
    END
  END sram_ro_data[29]
  PIN sram_ro_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1383.310 0.000 1383.590 4.000 ;
    END
  END sram_ro_data[2]
  PIN sram_ro_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1940.830 0.000 1941.110 4.000 ;
    END
  END sram_ro_data[30]
  PIN sram_ro_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1960.610 0.000 1960.890 4.000 ;
    END
  END sram_ro_data[31]
  PIN sram_ro_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1403.090 0.000 1403.370 4.000 ;
    END
  END sram_ro_data[3]
  PIN sram_ro_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1423.330 0.000 1423.610 4.000 ;
    END
  END sram_ro_data[4]
  PIN sram_ro_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1443.110 0.000 1443.390 4.000 ;
    END
  END sram_ro_data[5]
  PIN sram_ro_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.890 0.000 1463.170 4.000 ;
    END
  END sram_ro_data[6]
  PIN sram_ro_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1482.670 0.000 1482.950 4.000 ;
    END
  END sram_ro_data[7]
  PIN sram_ro_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1502.910 0.000 1503.190 4.000 ;
    END
  END sram_ro_data[8]
  PIN sram_ro_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1522.690 0.000 1522.970 4.000 ;
    END
  END sram_ro_data[9]
  PIN trap
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2179.570 0.000 2179.850 4.000 ;
    END
  END trap
  PIN uart_enabled
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2219.590 0.000 2219.870 4.000 ;
    END
  END uart_enabled
  PIN user_irq_ena[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2217.290 736.000 2217.570 740.000 ;
    END
  END user_irq_ena[0]
  PIN user_irq_ena[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2221.430 736.000 2221.710 740.000 ;
    END
  END user_irq_ena[1]
  PIN user_irq_ena[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2225.110 736.000 2225.390 740.000 ;
    END
  END user_irq_ena[2]
  OBS
      LAYER li1 ;
        RECT 5.520 7.905 2244.340 739.755 ;
      LAYER met1 ;
        RECT 1.450 0.720 2247.950 739.800 ;
      LAYER met2 ;
        RECT 1.480 735.720 1.650 739.830 ;
        RECT 2.490 735.720 5.330 739.830 ;
        RECT 6.170 735.720 9.010 739.830 ;
        RECT 9.850 735.720 12.690 739.830 ;
        RECT 13.530 735.720 16.370 739.830 ;
        RECT 17.210 735.720 20.510 739.830 ;
        RECT 21.350 735.720 24.190 739.830 ;
        RECT 25.030 735.720 27.870 739.830 ;
        RECT 28.710 735.720 31.550 739.830 ;
        RECT 32.390 735.720 35.690 739.830 ;
        RECT 36.530 735.720 39.370 739.830 ;
        RECT 40.210 735.720 43.050 739.830 ;
        RECT 43.890 735.720 46.730 739.830 ;
        RECT 47.570 735.720 50.870 739.830 ;
        RECT 51.710 735.720 54.550 739.830 ;
        RECT 55.390 735.720 58.230 739.830 ;
        RECT 59.070 735.720 61.910 739.830 ;
        RECT 62.750 735.720 66.050 739.830 ;
        RECT 66.890 735.720 69.730 739.830 ;
        RECT 70.570 735.720 73.410 739.830 ;
        RECT 74.250 735.720 77.090 739.830 ;
        RECT 77.930 735.720 81.230 739.830 ;
        RECT 82.070 735.720 84.910 739.830 ;
        RECT 85.750 735.720 88.590 739.830 ;
        RECT 89.430 735.720 92.270 739.830 ;
        RECT 93.110 735.720 96.410 739.830 ;
        RECT 97.250 735.720 100.090 739.830 ;
        RECT 100.930 735.720 103.770 739.830 ;
        RECT 104.610 735.720 107.450 739.830 ;
        RECT 108.290 735.720 111.590 739.830 ;
        RECT 112.430 735.720 115.270 739.830 ;
        RECT 116.110 735.720 118.950 739.830 ;
        RECT 119.790 735.720 122.630 739.830 ;
        RECT 123.470 735.720 126.770 739.830 ;
        RECT 127.610 735.720 130.450 739.830 ;
        RECT 131.290 735.720 134.130 739.830 ;
        RECT 134.970 735.720 137.810 739.830 ;
        RECT 138.650 735.720 141.950 739.830 ;
        RECT 142.790 735.720 145.630 739.830 ;
        RECT 146.470 735.720 149.310 739.830 ;
        RECT 150.150 735.720 152.990 739.830 ;
        RECT 153.830 735.720 157.130 739.830 ;
        RECT 157.970 735.720 160.810 739.830 ;
        RECT 161.650 735.720 164.490 739.830 ;
        RECT 165.330 735.720 168.170 739.830 ;
        RECT 169.010 735.720 172.310 739.830 ;
        RECT 173.150 735.720 175.990 739.830 ;
        RECT 176.830 735.720 179.670 739.830 ;
        RECT 180.510 735.720 183.350 739.830 ;
        RECT 184.190 735.720 187.490 739.830 ;
        RECT 188.330 735.720 191.170 739.830 ;
        RECT 192.010 735.720 194.850 739.830 ;
        RECT 195.690 735.720 198.530 739.830 ;
        RECT 199.370 735.720 202.670 739.830 ;
        RECT 203.510 735.720 206.350 739.830 ;
        RECT 207.190 735.720 210.030 739.830 ;
        RECT 210.870 735.720 213.710 739.830 ;
        RECT 214.550 735.720 217.850 739.830 ;
        RECT 218.690 735.720 221.530 739.830 ;
        RECT 222.370 735.720 225.210 739.830 ;
        RECT 226.050 735.720 228.890 739.830 ;
        RECT 229.730 735.720 233.030 739.830 ;
        RECT 233.870 735.720 236.710 739.830 ;
        RECT 237.550 735.720 240.390 739.830 ;
        RECT 241.230 735.720 244.070 739.830 ;
        RECT 244.910 735.720 248.210 739.830 ;
        RECT 249.050 735.720 251.890 739.830 ;
        RECT 252.730 735.720 255.570 739.830 ;
        RECT 256.410 735.720 259.250 739.830 ;
        RECT 260.090 735.720 263.390 739.830 ;
        RECT 264.230 735.720 267.070 739.830 ;
        RECT 267.910 735.720 270.750 739.830 ;
        RECT 271.590 735.720 274.430 739.830 ;
        RECT 275.270 735.720 278.570 739.830 ;
        RECT 279.410 735.720 282.250 739.830 ;
        RECT 283.090 735.720 285.930 739.830 ;
        RECT 286.770 735.720 289.610 739.830 ;
        RECT 290.450 735.720 293.750 739.830 ;
        RECT 294.590 735.720 297.430 739.830 ;
        RECT 298.270 735.720 301.110 739.830 ;
        RECT 301.950 735.720 304.790 739.830 ;
        RECT 305.630 735.720 308.930 739.830 ;
        RECT 309.770 735.720 312.610 739.830 ;
        RECT 313.450 735.720 316.290 739.830 ;
        RECT 317.130 735.720 319.970 739.830 ;
        RECT 320.810 735.720 324.110 739.830 ;
        RECT 324.950 735.720 327.790 739.830 ;
        RECT 328.630 735.720 331.470 739.830 ;
        RECT 332.310 735.720 335.150 739.830 ;
        RECT 335.990 735.720 339.290 739.830 ;
        RECT 340.130 735.720 342.970 739.830 ;
        RECT 343.810 735.720 346.650 739.830 ;
        RECT 347.490 735.720 350.330 739.830 ;
        RECT 351.170 735.720 354.470 739.830 ;
        RECT 355.310 735.720 358.150 739.830 ;
        RECT 358.990 735.720 361.830 739.830 ;
        RECT 362.670 735.720 365.510 739.830 ;
        RECT 366.350 735.720 369.650 739.830 ;
        RECT 370.490 735.720 373.330 739.830 ;
        RECT 374.170 735.720 377.010 739.830 ;
        RECT 377.850 735.720 380.690 739.830 ;
        RECT 381.530 735.720 384.830 739.830 ;
        RECT 385.670 735.720 388.510 739.830 ;
        RECT 389.350 735.720 392.190 739.830 ;
        RECT 393.030 735.720 395.870 739.830 ;
        RECT 396.710 735.720 400.010 739.830 ;
        RECT 400.850 735.720 403.690 739.830 ;
        RECT 404.530 735.720 407.370 739.830 ;
        RECT 408.210 735.720 411.050 739.830 ;
        RECT 411.890 735.720 415.190 739.830 ;
        RECT 416.030 735.720 418.870 739.830 ;
        RECT 419.710 735.720 422.550 739.830 ;
        RECT 423.390 735.720 426.230 739.830 ;
        RECT 427.070 735.720 430.370 739.830 ;
        RECT 431.210 735.720 434.050 739.830 ;
        RECT 434.890 735.720 437.730 739.830 ;
        RECT 438.570 735.720 441.410 739.830 ;
        RECT 442.250 735.720 445.550 739.830 ;
        RECT 446.390 735.720 449.230 739.830 ;
        RECT 450.070 735.720 452.910 739.830 ;
        RECT 453.750 735.720 456.590 739.830 ;
        RECT 457.430 735.720 460.270 739.830 ;
        RECT 461.110 735.720 464.410 739.830 ;
        RECT 465.250 735.720 468.090 739.830 ;
        RECT 468.930 735.720 471.770 739.830 ;
        RECT 472.610 735.720 475.450 739.830 ;
        RECT 476.290 735.720 479.590 739.830 ;
        RECT 480.430 735.720 483.270 739.830 ;
        RECT 484.110 735.720 486.950 739.830 ;
        RECT 487.790 735.720 490.630 739.830 ;
        RECT 491.470 735.720 494.770 739.830 ;
        RECT 495.610 735.720 498.450 739.830 ;
        RECT 499.290 735.720 502.130 739.830 ;
        RECT 502.970 735.720 505.810 739.830 ;
        RECT 506.650 735.720 509.950 739.830 ;
        RECT 510.790 735.720 513.630 739.830 ;
        RECT 514.470 735.720 517.310 739.830 ;
        RECT 518.150 735.720 520.990 739.830 ;
        RECT 521.830 735.720 525.130 739.830 ;
        RECT 525.970 735.720 528.810 739.830 ;
        RECT 529.650 735.720 532.490 739.830 ;
        RECT 533.330 735.720 536.170 739.830 ;
        RECT 537.010 735.720 540.310 739.830 ;
        RECT 541.150 735.720 543.990 739.830 ;
        RECT 544.830 735.720 547.670 739.830 ;
        RECT 548.510 735.720 551.350 739.830 ;
        RECT 552.190 735.720 555.490 739.830 ;
        RECT 556.330 735.720 559.170 739.830 ;
        RECT 560.010 735.720 562.850 739.830 ;
        RECT 563.690 735.720 566.530 739.830 ;
        RECT 567.370 735.720 570.670 739.830 ;
        RECT 571.510 735.720 574.350 739.830 ;
        RECT 575.190 735.720 578.030 739.830 ;
        RECT 578.870 735.720 581.710 739.830 ;
        RECT 582.550 735.720 585.850 739.830 ;
        RECT 586.690 735.720 589.530 739.830 ;
        RECT 590.370 735.720 593.210 739.830 ;
        RECT 594.050 735.720 596.890 739.830 ;
        RECT 597.730 735.720 601.030 739.830 ;
        RECT 601.870 735.720 604.710 739.830 ;
        RECT 605.550 735.720 608.390 739.830 ;
        RECT 609.230 735.720 612.070 739.830 ;
        RECT 612.910 735.720 616.210 739.830 ;
        RECT 617.050 735.720 619.890 739.830 ;
        RECT 620.730 735.720 623.570 739.830 ;
        RECT 624.410 735.720 627.250 739.830 ;
        RECT 628.090 735.720 631.390 739.830 ;
        RECT 632.230 735.720 635.070 739.830 ;
        RECT 635.910 735.720 638.750 739.830 ;
        RECT 639.590 735.720 642.430 739.830 ;
        RECT 643.270 735.720 646.570 739.830 ;
        RECT 647.410 735.720 650.250 739.830 ;
        RECT 651.090 735.720 653.930 739.830 ;
        RECT 654.770 735.720 657.610 739.830 ;
        RECT 658.450 735.720 661.750 739.830 ;
        RECT 662.590 735.720 665.430 739.830 ;
        RECT 666.270 735.720 669.110 739.830 ;
        RECT 669.950 735.720 672.790 739.830 ;
        RECT 673.630 735.720 676.930 739.830 ;
        RECT 677.770 735.720 680.610 739.830 ;
        RECT 681.450 735.720 684.290 739.830 ;
        RECT 685.130 735.720 687.970 739.830 ;
        RECT 688.810 735.720 692.110 739.830 ;
        RECT 692.950 735.720 695.790 739.830 ;
        RECT 696.630 735.720 699.470 739.830 ;
        RECT 700.310 735.720 703.150 739.830 ;
        RECT 703.990 735.720 707.290 739.830 ;
        RECT 708.130 735.720 710.970 739.830 ;
        RECT 711.810 735.720 714.650 739.830 ;
        RECT 715.490 735.720 718.330 739.830 ;
        RECT 719.170 735.720 722.470 739.830 ;
        RECT 723.310 735.720 726.150 739.830 ;
        RECT 726.990 735.720 729.830 739.830 ;
        RECT 730.670 735.720 733.510 739.830 ;
        RECT 734.350 735.720 737.650 739.830 ;
        RECT 738.490 735.720 741.330 739.830 ;
        RECT 742.170 735.720 745.010 739.830 ;
        RECT 745.850 735.720 748.690 739.830 ;
        RECT 749.530 735.720 752.830 739.830 ;
        RECT 753.670 735.720 756.510 739.830 ;
        RECT 757.350 735.720 760.190 739.830 ;
        RECT 761.030 735.720 763.870 739.830 ;
        RECT 764.710 735.720 768.010 739.830 ;
        RECT 768.850 735.720 771.690 739.830 ;
        RECT 772.530 735.720 775.370 739.830 ;
        RECT 776.210 735.720 779.050 739.830 ;
        RECT 779.890 735.720 783.190 739.830 ;
        RECT 784.030 735.720 786.870 739.830 ;
        RECT 787.710 735.720 790.550 739.830 ;
        RECT 791.390 735.720 794.230 739.830 ;
        RECT 795.070 735.720 798.370 739.830 ;
        RECT 799.210 735.720 802.050 739.830 ;
        RECT 802.890 735.720 805.730 739.830 ;
        RECT 806.570 735.720 809.410 739.830 ;
        RECT 810.250 735.720 813.550 739.830 ;
        RECT 814.390 735.720 817.230 739.830 ;
        RECT 818.070 735.720 820.910 739.830 ;
        RECT 821.750 735.720 824.590 739.830 ;
        RECT 825.430 735.720 828.730 739.830 ;
        RECT 829.570 735.720 832.410 739.830 ;
        RECT 833.250 735.720 836.090 739.830 ;
        RECT 836.930 735.720 839.770 739.830 ;
        RECT 840.610 735.720 843.910 739.830 ;
        RECT 844.750 735.720 847.590 739.830 ;
        RECT 848.430 735.720 851.270 739.830 ;
        RECT 852.110 735.720 854.950 739.830 ;
        RECT 855.790 735.720 859.090 739.830 ;
        RECT 859.930 735.720 862.770 739.830 ;
        RECT 863.610 735.720 866.450 739.830 ;
        RECT 867.290 735.720 870.130 739.830 ;
        RECT 870.970 735.720 874.270 739.830 ;
        RECT 875.110 735.720 877.950 739.830 ;
        RECT 878.790 735.720 881.630 739.830 ;
        RECT 882.470 735.720 885.310 739.830 ;
        RECT 886.150 735.720 889.450 739.830 ;
        RECT 890.290 735.720 893.130 739.830 ;
        RECT 893.970 735.720 896.810 739.830 ;
        RECT 897.650 735.720 900.490 739.830 ;
        RECT 901.330 735.720 904.170 739.830 ;
        RECT 905.010 735.720 908.310 739.830 ;
        RECT 909.150 735.720 911.990 739.830 ;
        RECT 912.830 735.720 915.670 739.830 ;
        RECT 916.510 735.720 919.350 739.830 ;
        RECT 920.190 735.720 923.490 739.830 ;
        RECT 924.330 735.720 927.170 739.830 ;
        RECT 928.010 735.720 930.850 739.830 ;
        RECT 931.690 735.720 934.530 739.830 ;
        RECT 935.370 735.720 938.670 739.830 ;
        RECT 939.510 735.720 942.350 739.830 ;
        RECT 943.190 735.720 946.030 739.830 ;
        RECT 946.870 735.720 949.710 739.830 ;
        RECT 950.550 735.720 953.850 739.830 ;
        RECT 954.690 735.720 957.530 739.830 ;
        RECT 958.370 735.720 961.210 739.830 ;
        RECT 962.050 735.720 964.890 739.830 ;
        RECT 965.730 735.720 969.030 739.830 ;
        RECT 969.870 735.720 972.710 739.830 ;
        RECT 973.550 735.720 976.390 739.830 ;
        RECT 977.230 735.720 980.070 739.830 ;
        RECT 980.910 735.720 984.210 739.830 ;
        RECT 985.050 735.720 987.890 739.830 ;
        RECT 988.730 735.720 991.570 739.830 ;
        RECT 992.410 735.720 995.250 739.830 ;
        RECT 996.090 735.720 999.390 739.830 ;
        RECT 1000.230 735.720 1003.070 739.830 ;
        RECT 1003.910 735.720 1006.750 739.830 ;
        RECT 1007.590 735.720 1010.430 739.830 ;
        RECT 1011.270 735.720 1014.570 739.830 ;
        RECT 1015.410 735.720 1018.250 739.830 ;
        RECT 1019.090 735.720 1021.930 739.830 ;
        RECT 1022.770 735.720 1025.610 739.830 ;
        RECT 1026.450 735.720 1029.750 739.830 ;
        RECT 1030.590 735.720 1033.430 739.830 ;
        RECT 1034.270 735.720 1037.110 739.830 ;
        RECT 1037.950 735.720 1040.790 739.830 ;
        RECT 1041.630 735.720 1044.930 739.830 ;
        RECT 1045.770 735.720 1048.610 739.830 ;
        RECT 1049.450 735.720 1052.290 739.830 ;
        RECT 1053.130 735.720 1055.970 739.830 ;
        RECT 1056.810 735.720 1060.110 739.830 ;
        RECT 1060.950 735.720 1063.790 739.830 ;
        RECT 1064.630 735.720 1067.470 739.830 ;
        RECT 1068.310 735.720 1071.150 739.830 ;
        RECT 1071.990 735.720 1075.290 739.830 ;
        RECT 1076.130 735.720 1078.970 739.830 ;
        RECT 1079.810 735.720 1082.650 739.830 ;
        RECT 1083.490 735.720 1086.330 739.830 ;
        RECT 1087.170 735.720 1090.470 739.830 ;
        RECT 1091.310 735.720 1094.150 739.830 ;
        RECT 1094.990 735.720 1097.830 739.830 ;
        RECT 1098.670 735.720 1101.510 739.830 ;
        RECT 1102.350 735.720 1105.650 739.830 ;
        RECT 1106.490 735.720 1109.330 739.830 ;
        RECT 1110.170 735.720 1113.010 739.830 ;
        RECT 1113.850 735.720 1116.690 739.830 ;
        RECT 1117.530 735.720 1120.830 739.830 ;
        RECT 1121.670 735.720 1124.510 739.830 ;
        RECT 1125.350 735.720 1128.190 739.830 ;
        RECT 1129.030 735.720 1131.870 739.830 ;
        RECT 1132.710 735.720 1136.010 739.830 ;
        RECT 1136.850 735.720 1139.690 739.830 ;
        RECT 1140.530 735.720 1143.370 739.830 ;
        RECT 1144.210 735.720 1147.050 739.830 ;
        RECT 1147.890 735.720 1151.190 739.830 ;
        RECT 1152.030 735.720 1154.870 739.830 ;
        RECT 1155.710 735.720 1158.550 739.830 ;
        RECT 1159.390 735.720 1162.230 739.830 ;
        RECT 1163.070 735.720 1166.370 739.830 ;
        RECT 1167.210 735.720 1170.050 739.830 ;
        RECT 1170.890 735.720 1173.730 739.830 ;
        RECT 1174.570 735.720 1177.410 739.830 ;
        RECT 1178.250 735.720 1181.550 739.830 ;
        RECT 1182.390 735.720 1185.230 739.830 ;
        RECT 1186.070 735.720 1188.910 739.830 ;
        RECT 1189.750 735.720 1192.590 739.830 ;
        RECT 1193.430 735.720 1196.730 739.830 ;
        RECT 1197.570 735.720 1200.410 739.830 ;
        RECT 1201.250 735.720 1204.090 739.830 ;
        RECT 1204.930 735.720 1207.770 739.830 ;
        RECT 1208.610 735.720 1211.910 739.830 ;
        RECT 1212.750 735.720 1215.590 739.830 ;
        RECT 1216.430 735.720 1219.270 739.830 ;
        RECT 1220.110 735.720 1222.950 739.830 ;
        RECT 1223.790 735.720 1227.090 739.830 ;
        RECT 1227.930 735.720 1230.770 739.830 ;
        RECT 1231.610 735.720 1234.450 739.830 ;
        RECT 1235.290 735.720 1238.130 739.830 ;
        RECT 1238.970 735.720 1242.270 739.830 ;
        RECT 1243.110 735.720 1245.950 739.830 ;
        RECT 1246.790 735.720 1249.630 739.830 ;
        RECT 1250.470 735.720 1253.310 739.830 ;
        RECT 1254.150 735.720 1257.450 739.830 ;
        RECT 1258.290 735.720 1261.130 739.830 ;
        RECT 1261.970 735.720 1264.810 739.830 ;
        RECT 1265.650 735.720 1268.490 739.830 ;
        RECT 1269.330 735.720 1272.630 739.830 ;
        RECT 1273.470 735.720 1276.310 739.830 ;
        RECT 1277.150 735.720 1279.990 739.830 ;
        RECT 1280.830 735.720 1283.670 739.830 ;
        RECT 1284.510 735.720 1287.810 739.830 ;
        RECT 1288.650 735.720 1291.490 739.830 ;
        RECT 1292.330 735.720 1295.170 739.830 ;
        RECT 1296.010 735.720 1298.850 739.830 ;
        RECT 1299.690 735.720 1302.990 739.830 ;
        RECT 1303.830 735.720 1306.670 739.830 ;
        RECT 1307.510 735.720 1310.350 739.830 ;
        RECT 1311.190 735.720 1314.030 739.830 ;
        RECT 1314.870 735.720 1318.170 739.830 ;
        RECT 1319.010 735.720 1321.850 739.830 ;
        RECT 1322.690 735.720 1325.530 739.830 ;
        RECT 1326.370 735.720 1329.210 739.830 ;
        RECT 1330.050 735.720 1333.350 739.830 ;
        RECT 1334.190 735.720 1337.030 739.830 ;
        RECT 1337.870 735.720 1340.710 739.830 ;
        RECT 1341.550 735.720 1344.390 739.830 ;
        RECT 1345.230 735.720 1348.530 739.830 ;
        RECT 1349.370 735.720 1352.210 739.830 ;
        RECT 1353.050 735.720 1355.890 739.830 ;
        RECT 1356.730 735.720 1359.570 739.830 ;
        RECT 1360.410 735.720 1363.250 739.830 ;
        RECT 1364.090 735.720 1367.390 739.830 ;
        RECT 1368.230 735.720 1371.070 739.830 ;
        RECT 1371.910 735.720 1374.750 739.830 ;
        RECT 1375.590 735.720 1378.430 739.830 ;
        RECT 1379.270 735.720 1382.570 739.830 ;
        RECT 1383.410 735.720 1386.250 739.830 ;
        RECT 1387.090 735.720 1389.930 739.830 ;
        RECT 1390.770 735.720 1393.610 739.830 ;
        RECT 1394.450 735.720 1397.750 739.830 ;
        RECT 1398.590 735.720 1401.430 739.830 ;
        RECT 1402.270 735.720 1405.110 739.830 ;
        RECT 1405.950 735.720 1408.790 739.830 ;
        RECT 1409.630 735.720 1412.930 739.830 ;
        RECT 1413.770 735.720 1416.610 739.830 ;
        RECT 1417.450 735.720 1420.290 739.830 ;
        RECT 1421.130 735.720 1423.970 739.830 ;
        RECT 1424.810 735.720 1428.110 739.830 ;
        RECT 1428.950 735.720 1431.790 739.830 ;
        RECT 1432.630 735.720 1435.470 739.830 ;
        RECT 1436.310 735.720 1439.150 739.830 ;
        RECT 1439.990 735.720 1443.290 739.830 ;
        RECT 1444.130 735.720 1446.970 739.830 ;
        RECT 1447.810 735.720 1450.650 739.830 ;
        RECT 1451.490 735.720 1454.330 739.830 ;
        RECT 1455.170 735.720 1458.470 739.830 ;
        RECT 1459.310 735.720 1462.150 739.830 ;
        RECT 1462.990 735.720 1465.830 739.830 ;
        RECT 1466.670 735.720 1469.510 739.830 ;
        RECT 1470.350 735.720 1473.650 739.830 ;
        RECT 1474.490 735.720 1477.330 739.830 ;
        RECT 1478.170 735.720 1481.010 739.830 ;
        RECT 1481.850 735.720 1484.690 739.830 ;
        RECT 1485.530 735.720 1488.830 739.830 ;
        RECT 1489.670 735.720 1492.510 739.830 ;
        RECT 1493.350 735.720 1496.190 739.830 ;
        RECT 1497.030 735.720 1499.870 739.830 ;
        RECT 1500.710 735.720 1504.010 739.830 ;
        RECT 1504.850 735.720 1507.690 739.830 ;
        RECT 1508.530 735.720 1511.370 739.830 ;
        RECT 1512.210 735.720 1515.050 739.830 ;
        RECT 1515.890 735.720 1519.190 739.830 ;
        RECT 1520.030 735.720 1522.870 739.830 ;
        RECT 1523.710 735.720 1526.550 739.830 ;
        RECT 1527.390 735.720 1530.230 739.830 ;
        RECT 1531.070 735.720 1534.370 739.830 ;
        RECT 1535.210 735.720 1538.050 739.830 ;
        RECT 1538.890 735.720 1541.730 739.830 ;
        RECT 1542.570 735.720 1545.410 739.830 ;
        RECT 1546.250 735.720 1549.550 739.830 ;
        RECT 1550.390 735.720 1553.230 739.830 ;
        RECT 1554.070 735.720 1556.910 739.830 ;
        RECT 1557.750 735.720 1560.590 739.830 ;
        RECT 1561.430 735.720 1564.730 739.830 ;
        RECT 1565.570 735.720 1568.410 739.830 ;
        RECT 1569.250 735.720 1572.090 739.830 ;
        RECT 1572.930 735.720 1575.770 739.830 ;
        RECT 1576.610 735.720 1579.910 739.830 ;
        RECT 1580.750 735.720 1583.590 739.830 ;
        RECT 1584.430 735.720 1587.270 739.830 ;
        RECT 1588.110 735.720 1590.950 739.830 ;
        RECT 1591.790 735.720 1595.090 739.830 ;
        RECT 1595.930 735.720 1598.770 739.830 ;
        RECT 1599.610 735.720 1602.450 739.830 ;
        RECT 1603.290 735.720 1606.130 739.830 ;
        RECT 1606.970 735.720 1610.270 739.830 ;
        RECT 1611.110 735.720 1613.950 739.830 ;
        RECT 1614.790 735.720 1617.630 739.830 ;
        RECT 1618.470 735.720 1621.310 739.830 ;
        RECT 1622.150 735.720 1625.450 739.830 ;
        RECT 1626.290 735.720 1629.130 739.830 ;
        RECT 1629.970 735.720 1632.810 739.830 ;
        RECT 1633.650 735.720 1636.490 739.830 ;
        RECT 1637.330 735.720 1640.630 739.830 ;
        RECT 1641.470 735.720 1644.310 739.830 ;
        RECT 1645.150 735.720 1647.990 739.830 ;
        RECT 1648.830 735.720 1651.670 739.830 ;
        RECT 1652.510 735.720 1655.810 739.830 ;
        RECT 1656.650 735.720 1659.490 739.830 ;
        RECT 1660.330 735.720 1663.170 739.830 ;
        RECT 1664.010 735.720 1666.850 739.830 ;
        RECT 1667.690 735.720 1670.990 739.830 ;
        RECT 1671.830 735.720 1674.670 739.830 ;
        RECT 1675.510 735.720 1678.350 739.830 ;
        RECT 1679.190 735.720 1682.030 739.830 ;
        RECT 1682.870 735.720 1686.170 739.830 ;
        RECT 1687.010 735.720 1689.850 739.830 ;
        RECT 1690.690 735.720 1693.530 739.830 ;
        RECT 1694.370 735.720 1697.210 739.830 ;
        RECT 1698.050 735.720 1701.350 739.830 ;
        RECT 1702.190 735.720 1705.030 739.830 ;
        RECT 1705.870 735.720 1708.710 739.830 ;
        RECT 1709.550 735.720 1712.390 739.830 ;
        RECT 1713.230 735.720 1716.530 739.830 ;
        RECT 1717.370 735.720 1720.210 739.830 ;
        RECT 1721.050 735.720 1723.890 739.830 ;
        RECT 1724.730 735.720 1727.570 739.830 ;
        RECT 1728.410 735.720 1731.710 739.830 ;
        RECT 1732.550 735.720 1735.390 739.830 ;
        RECT 1736.230 735.720 1739.070 739.830 ;
        RECT 1739.910 735.720 1742.750 739.830 ;
        RECT 1743.590 735.720 1746.890 739.830 ;
        RECT 1747.730 735.720 1750.570 739.830 ;
        RECT 1751.410 735.720 1754.250 739.830 ;
        RECT 1755.090 735.720 1757.930 739.830 ;
        RECT 1758.770 735.720 1762.070 739.830 ;
        RECT 1762.910 735.720 1765.750 739.830 ;
        RECT 1766.590 735.720 1769.430 739.830 ;
        RECT 1770.270 735.720 1773.110 739.830 ;
        RECT 1773.950 735.720 1777.250 739.830 ;
        RECT 1778.090 735.720 1780.930 739.830 ;
        RECT 1781.770 735.720 1784.610 739.830 ;
        RECT 1785.450 735.720 1788.290 739.830 ;
        RECT 1789.130 735.720 1792.430 739.830 ;
        RECT 1793.270 735.720 1796.110 739.830 ;
        RECT 1796.950 735.720 1799.790 739.830 ;
        RECT 1800.630 735.720 1803.470 739.830 ;
        RECT 1804.310 735.720 1807.150 739.830 ;
        RECT 1807.990 735.720 1811.290 739.830 ;
        RECT 1812.130 735.720 1814.970 739.830 ;
        RECT 1815.810 735.720 1818.650 739.830 ;
        RECT 1819.490 735.720 1822.330 739.830 ;
        RECT 1823.170 735.720 1826.470 739.830 ;
        RECT 1827.310 735.720 1830.150 739.830 ;
        RECT 1830.990 735.720 1833.830 739.830 ;
        RECT 1834.670 735.720 1837.510 739.830 ;
        RECT 1838.350 735.720 1841.650 739.830 ;
        RECT 1842.490 735.720 1845.330 739.830 ;
        RECT 1846.170 735.720 1849.010 739.830 ;
        RECT 1849.850 735.720 1852.690 739.830 ;
        RECT 1853.530 735.720 1856.830 739.830 ;
        RECT 1857.670 735.720 1860.510 739.830 ;
        RECT 1861.350 735.720 1864.190 739.830 ;
        RECT 1865.030 735.720 1867.870 739.830 ;
        RECT 1868.710 735.720 1872.010 739.830 ;
        RECT 1872.850 735.720 1875.690 739.830 ;
        RECT 1876.530 735.720 1879.370 739.830 ;
        RECT 1880.210 735.720 1883.050 739.830 ;
        RECT 1883.890 735.720 1887.190 739.830 ;
        RECT 1888.030 735.720 1890.870 739.830 ;
        RECT 1891.710 735.720 1894.550 739.830 ;
        RECT 1895.390 735.720 1898.230 739.830 ;
        RECT 1899.070 735.720 1902.370 739.830 ;
        RECT 1903.210 735.720 1906.050 739.830 ;
        RECT 1906.890 735.720 1909.730 739.830 ;
        RECT 1910.570 735.720 1913.410 739.830 ;
        RECT 1914.250 735.720 1917.550 739.830 ;
        RECT 1918.390 735.720 1921.230 739.830 ;
        RECT 1922.070 735.720 1924.910 739.830 ;
        RECT 1925.750 735.720 1928.590 739.830 ;
        RECT 1929.430 735.720 1932.730 739.830 ;
        RECT 1933.570 735.720 1936.410 739.830 ;
        RECT 1937.250 735.720 1940.090 739.830 ;
        RECT 1940.930 735.720 1943.770 739.830 ;
        RECT 1944.610 735.720 1947.910 739.830 ;
        RECT 1948.750 735.720 1951.590 739.830 ;
        RECT 1952.430 735.720 1955.270 739.830 ;
        RECT 1956.110 735.720 1958.950 739.830 ;
        RECT 1959.790 735.720 1963.090 739.830 ;
        RECT 1963.930 735.720 1966.770 739.830 ;
        RECT 1967.610 735.720 1970.450 739.830 ;
        RECT 1971.290 735.720 1974.130 739.830 ;
        RECT 1974.970 735.720 1978.270 739.830 ;
        RECT 1979.110 735.720 1981.950 739.830 ;
        RECT 1982.790 735.720 1985.630 739.830 ;
        RECT 1986.470 735.720 1989.310 739.830 ;
        RECT 1990.150 735.720 1993.450 739.830 ;
        RECT 1994.290 735.720 1997.130 739.830 ;
        RECT 1997.970 735.720 2000.810 739.830 ;
        RECT 2001.650 735.720 2004.490 739.830 ;
        RECT 2005.330 735.720 2008.630 739.830 ;
        RECT 2009.470 735.720 2012.310 739.830 ;
        RECT 2013.150 735.720 2015.990 739.830 ;
        RECT 2016.830 735.720 2019.670 739.830 ;
        RECT 2020.510 735.720 2023.810 739.830 ;
        RECT 2024.650 735.720 2027.490 739.830 ;
        RECT 2028.330 735.720 2031.170 739.830 ;
        RECT 2032.010 735.720 2034.850 739.830 ;
        RECT 2035.690 735.720 2038.990 739.830 ;
        RECT 2039.830 735.720 2042.670 739.830 ;
        RECT 2043.510 735.720 2046.350 739.830 ;
        RECT 2047.190 735.720 2050.030 739.830 ;
        RECT 2050.870 735.720 2054.170 739.830 ;
        RECT 2055.010 735.720 2057.850 739.830 ;
        RECT 2058.690 735.720 2061.530 739.830 ;
        RECT 2062.370 735.720 2065.210 739.830 ;
        RECT 2066.050 735.720 2069.350 739.830 ;
        RECT 2070.190 735.720 2073.030 739.830 ;
        RECT 2073.870 735.720 2076.710 739.830 ;
        RECT 2077.550 735.720 2080.390 739.830 ;
        RECT 2081.230 735.720 2084.530 739.830 ;
        RECT 2085.370 735.720 2088.210 739.830 ;
        RECT 2089.050 735.720 2091.890 739.830 ;
        RECT 2092.730 735.720 2095.570 739.830 ;
        RECT 2096.410 735.720 2099.710 739.830 ;
        RECT 2100.550 735.720 2103.390 739.830 ;
        RECT 2104.230 735.720 2107.070 739.830 ;
        RECT 2107.910 735.720 2110.750 739.830 ;
        RECT 2111.590 735.720 2114.890 739.830 ;
        RECT 2115.730 735.720 2118.570 739.830 ;
        RECT 2119.410 735.720 2122.250 739.830 ;
        RECT 2123.090 735.720 2125.930 739.830 ;
        RECT 2126.770 735.720 2130.070 739.830 ;
        RECT 2130.910 735.720 2133.750 739.830 ;
        RECT 2134.590 735.720 2137.430 739.830 ;
        RECT 2138.270 735.720 2141.110 739.830 ;
        RECT 2141.950 735.720 2145.250 739.830 ;
        RECT 2146.090 735.720 2148.930 739.830 ;
        RECT 2149.770 735.720 2152.610 739.830 ;
        RECT 2153.450 735.720 2156.290 739.830 ;
        RECT 2157.130 735.720 2160.430 739.830 ;
        RECT 2161.270 735.720 2164.110 739.830 ;
        RECT 2164.950 735.720 2167.790 739.830 ;
        RECT 2168.630 735.720 2171.470 739.830 ;
        RECT 2172.310 735.720 2175.610 739.830 ;
        RECT 2176.450 735.720 2179.290 739.830 ;
        RECT 2180.130 735.720 2182.970 739.830 ;
        RECT 2183.810 735.720 2186.650 739.830 ;
        RECT 2187.490 735.720 2190.790 739.830 ;
        RECT 2191.630 735.720 2194.470 739.830 ;
        RECT 2195.310 735.720 2198.150 739.830 ;
        RECT 2198.990 735.720 2201.830 739.830 ;
        RECT 2202.670 735.720 2205.970 739.830 ;
        RECT 2206.810 735.720 2209.650 739.830 ;
        RECT 2210.490 735.720 2213.330 739.830 ;
        RECT 2214.170 735.720 2217.010 739.830 ;
        RECT 2217.850 735.720 2221.150 739.830 ;
        RECT 2221.990 735.720 2224.830 739.830 ;
        RECT 2225.670 735.720 2228.510 739.830 ;
        RECT 2229.350 735.720 2232.190 739.830 ;
        RECT 2233.030 735.720 2236.330 739.830 ;
        RECT 2237.170 735.720 2240.010 739.830 ;
        RECT 2240.850 735.720 2243.690 739.830 ;
        RECT 2244.530 735.720 2247.370 739.830 ;
        RECT 1.480 4.280 2247.920 735.720 ;
        RECT 1.480 0.690 9.470 4.280 ;
        RECT 10.310 0.690 29.250 4.280 ;
        RECT 30.090 0.690 49.030 4.280 ;
        RECT 49.870 0.690 68.810 4.280 ;
        RECT 69.650 0.690 89.050 4.280 ;
        RECT 89.890 0.690 108.830 4.280 ;
        RECT 109.670 0.690 128.610 4.280 ;
        RECT 129.450 0.690 148.390 4.280 ;
        RECT 149.230 0.690 168.630 4.280 ;
        RECT 169.470 0.690 188.410 4.280 ;
        RECT 189.250 0.690 208.190 4.280 ;
        RECT 209.030 0.690 228.430 4.280 ;
        RECT 229.270 0.690 248.210 4.280 ;
        RECT 249.050 0.690 267.990 4.280 ;
        RECT 268.830 0.690 287.770 4.280 ;
        RECT 288.610 0.690 308.010 4.280 ;
        RECT 308.850 0.690 327.790 4.280 ;
        RECT 328.630 0.690 347.570 4.280 ;
        RECT 348.410 0.690 367.810 4.280 ;
        RECT 368.650 0.690 387.590 4.280 ;
        RECT 388.430 0.690 407.370 4.280 ;
        RECT 408.210 0.690 427.150 4.280 ;
        RECT 427.990 0.690 447.390 4.280 ;
        RECT 448.230 0.690 467.170 4.280 ;
        RECT 468.010 0.690 486.950 4.280 ;
        RECT 487.790 0.690 507.190 4.280 ;
        RECT 508.030 0.690 526.970 4.280 ;
        RECT 527.810 0.690 546.750 4.280 ;
        RECT 547.590 0.690 566.530 4.280 ;
        RECT 567.370 0.690 586.770 4.280 ;
        RECT 587.610 0.690 606.550 4.280 ;
        RECT 607.390 0.690 626.330 4.280 ;
        RECT 627.170 0.690 646.570 4.280 ;
        RECT 647.410 0.690 666.350 4.280 ;
        RECT 667.190 0.690 686.130 4.280 ;
        RECT 686.970 0.690 705.910 4.280 ;
        RECT 706.750 0.690 726.150 4.280 ;
        RECT 726.990 0.690 745.930 4.280 ;
        RECT 746.770 0.690 765.710 4.280 ;
        RECT 766.550 0.690 785.950 4.280 ;
        RECT 786.790 0.690 805.730 4.280 ;
        RECT 806.570 0.690 825.510 4.280 ;
        RECT 826.350 0.690 845.290 4.280 ;
        RECT 846.130 0.690 865.530 4.280 ;
        RECT 866.370 0.690 885.310 4.280 ;
        RECT 886.150 0.690 905.090 4.280 ;
        RECT 905.930 0.690 925.330 4.280 ;
        RECT 926.170 0.690 945.110 4.280 ;
        RECT 945.950 0.690 964.890 4.280 ;
        RECT 965.730 0.690 984.670 4.280 ;
        RECT 985.510 0.690 1004.910 4.280 ;
        RECT 1005.750 0.690 1024.690 4.280 ;
        RECT 1025.530 0.690 1044.470 4.280 ;
        RECT 1045.310 0.690 1064.710 4.280 ;
        RECT 1065.550 0.690 1084.490 4.280 ;
        RECT 1085.330 0.690 1104.270 4.280 ;
        RECT 1105.110 0.690 1124.050 4.280 ;
        RECT 1124.890 0.690 1144.290 4.280 ;
        RECT 1145.130 0.690 1164.070 4.280 ;
        RECT 1164.910 0.690 1183.850 4.280 ;
        RECT 1184.690 0.690 1203.630 4.280 ;
        RECT 1204.470 0.690 1223.870 4.280 ;
        RECT 1224.710 0.690 1243.650 4.280 ;
        RECT 1244.490 0.690 1263.430 4.280 ;
        RECT 1264.270 0.690 1283.670 4.280 ;
        RECT 1284.510 0.690 1303.450 4.280 ;
        RECT 1304.290 0.690 1323.230 4.280 ;
        RECT 1324.070 0.690 1343.010 4.280 ;
        RECT 1343.850 0.690 1363.250 4.280 ;
        RECT 1364.090 0.690 1383.030 4.280 ;
        RECT 1383.870 0.690 1402.810 4.280 ;
        RECT 1403.650 0.690 1423.050 4.280 ;
        RECT 1423.890 0.690 1442.830 4.280 ;
        RECT 1443.670 0.690 1462.610 4.280 ;
        RECT 1463.450 0.690 1482.390 4.280 ;
        RECT 1483.230 0.690 1502.630 4.280 ;
        RECT 1503.470 0.690 1522.410 4.280 ;
        RECT 1523.250 0.690 1542.190 4.280 ;
        RECT 1543.030 0.690 1562.430 4.280 ;
        RECT 1563.270 0.690 1582.210 4.280 ;
        RECT 1583.050 0.690 1601.990 4.280 ;
        RECT 1602.830 0.690 1621.770 4.280 ;
        RECT 1622.610 0.690 1642.010 4.280 ;
        RECT 1642.850 0.690 1661.790 4.280 ;
        RECT 1662.630 0.690 1681.570 4.280 ;
        RECT 1682.410 0.690 1701.810 4.280 ;
        RECT 1702.650 0.690 1721.590 4.280 ;
        RECT 1722.430 0.690 1741.370 4.280 ;
        RECT 1742.210 0.690 1761.150 4.280 ;
        RECT 1761.990 0.690 1781.390 4.280 ;
        RECT 1782.230 0.690 1801.170 4.280 ;
        RECT 1802.010 0.690 1820.950 4.280 ;
        RECT 1821.790 0.690 1841.190 4.280 ;
        RECT 1842.030 0.690 1860.970 4.280 ;
        RECT 1861.810 0.690 1880.750 4.280 ;
        RECT 1881.590 0.690 1900.530 4.280 ;
        RECT 1901.370 0.690 1920.770 4.280 ;
        RECT 1921.610 0.690 1940.550 4.280 ;
        RECT 1941.390 0.690 1960.330 4.280 ;
        RECT 1961.170 0.690 1980.570 4.280 ;
        RECT 1981.410 0.690 2000.350 4.280 ;
        RECT 2001.190 0.690 2020.130 4.280 ;
        RECT 2020.970 0.690 2039.910 4.280 ;
        RECT 2040.750 0.690 2060.150 4.280 ;
        RECT 2060.990 0.690 2079.930 4.280 ;
        RECT 2080.770 0.690 2099.710 4.280 ;
        RECT 2100.550 0.690 2119.950 4.280 ;
        RECT 2120.790 0.690 2139.730 4.280 ;
        RECT 2140.570 0.690 2159.510 4.280 ;
        RECT 2160.350 0.690 2179.290 4.280 ;
        RECT 2180.130 0.690 2199.530 4.280 ;
        RECT 2200.370 0.690 2219.310 4.280 ;
        RECT 2220.150 0.690 2239.090 4.280 ;
        RECT 2239.930 0.690 2247.920 4.280 ;
      LAYER met3 ;
        RECT 2.365 736.800 2246.000 736.945 ;
        RECT 4.400 735.400 2246.000 736.800 ;
        RECT 2.365 730.000 2246.000 735.400 ;
        RECT 4.400 728.600 2246.000 730.000 ;
        RECT 2.365 723.200 2246.000 728.600 ;
        RECT 4.400 721.800 2246.000 723.200 ;
        RECT 2.365 717.080 2246.000 721.800 ;
        RECT 4.400 715.680 2246.000 717.080 ;
        RECT 2.365 710.280 2246.000 715.680 ;
        RECT 4.400 708.880 2246.000 710.280 ;
        RECT 2.365 703.480 2246.000 708.880 ;
        RECT 4.400 702.080 2246.000 703.480 ;
        RECT 2.365 697.360 2246.000 702.080 ;
        RECT 4.400 695.960 2246.000 697.360 ;
        RECT 2.365 690.560 2246.000 695.960 ;
        RECT 4.400 689.160 2246.000 690.560 ;
        RECT 2.365 683.760 2246.000 689.160 ;
        RECT 4.400 682.360 2246.000 683.760 ;
        RECT 2.365 676.960 2246.000 682.360 ;
        RECT 4.400 675.560 2246.000 676.960 ;
        RECT 2.365 670.840 2246.000 675.560 ;
        RECT 4.400 669.440 2246.000 670.840 ;
        RECT 2.365 664.040 2246.000 669.440 ;
        RECT 4.400 662.640 2246.000 664.040 ;
        RECT 2.365 657.240 2246.000 662.640 ;
        RECT 4.400 655.840 2246.000 657.240 ;
        RECT 2.365 651.120 2246.000 655.840 ;
        RECT 4.400 649.720 2246.000 651.120 ;
        RECT 2.365 644.320 2246.000 649.720 ;
        RECT 4.400 642.920 2246.000 644.320 ;
        RECT 2.365 637.520 2246.000 642.920 ;
        RECT 4.400 636.120 2246.000 637.520 ;
        RECT 2.365 630.720 2246.000 636.120 ;
        RECT 4.400 629.320 2246.000 630.720 ;
        RECT 2.365 624.600 2246.000 629.320 ;
        RECT 4.400 623.200 2246.000 624.600 ;
        RECT 2.365 617.800 2246.000 623.200 ;
        RECT 4.400 616.400 2246.000 617.800 ;
        RECT 2.365 611.000 2246.000 616.400 ;
        RECT 4.400 609.600 2246.000 611.000 ;
        RECT 2.365 604.880 2246.000 609.600 ;
        RECT 4.400 603.480 2246.000 604.880 ;
        RECT 2.365 598.080 2246.000 603.480 ;
        RECT 4.400 596.680 2246.000 598.080 ;
        RECT 2.365 591.280 2246.000 596.680 ;
        RECT 4.400 589.880 2246.000 591.280 ;
        RECT 2.365 584.480 2246.000 589.880 ;
        RECT 4.400 583.080 2246.000 584.480 ;
        RECT 2.365 578.360 2246.000 583.080 ;
        RECT 4.400 576.960 2246.000 578.360 ;
        RECT 2.365 571.560 2246.000 576.960 ;
        RECT 4.400 570.160 2246.000 571.560 ;
        RECT 2.365 564.760 2246.000 570.160 ;
        RECT 4.400 563.360 2246.000 564.760 ;
        RECT 2.365 558.640 2246.000 563.360 ;
        RECT 4.400 557.240 2246.000 558.640 ;
        RECT 2.365 555.920 2246.000 557.240 ;
        RECT 2.365 554.520 2245.600 555.920 ;
        RECT 2.365 551.840 2246.000 554.520 ;
        RECT 4.400 550.440 2246.000 551.840 ;
        RECT 2.365 545.040 2246.000 550.440 ;
        RECT 4.400 543.640 2246.000 545.040 ;
        RECT 2.365 538.240 2246.000 543.640 ;
        RECT 4.400 536.840 2246.000 538.240 ;
        RECT 2.365 532.120 2246.000 536.840 ;
        RECT 4.400 530.720 2246.000 532.120 ;
        RECT 2.365 525.320 2246.000 530.720 ;
        RECT 4.400 523.920 2246.000 525.320 ;
        RECT 2.365 518.520 2246.000 523.920 ;
        RECT 4.400 517.120 2246.000 518.520 ;
        RECT 2.365 512.400 2246.000 517.120 ;
        RECT 4.400 511.000 2246.000 512.400 ;
        RECT 2.365 505.600 2246.000 511.000 ;
        RECT 4.400 504.200 2246.000 505.600 ;
        RECT 2.365 498.800 2246.000 504.200 ;
        RECT 4.400 497.400 2246.000 498.800 ;
        RECT 2.365 492.000 2246.000 497.400 ;
        RECT 4.400 490.600 2246.000 492.000 ;
        RECT 2.365 485.880 2246.000 490.600 ;
        RECT 4.400 484.480 2246.000 485.880 ;
        RECT 2.365 479.080 2246.000 484.480 ;
        RECT 4.400 477.680 2246.000 479.080 ;
        RECT 2.365 472.280 2246.000 477.680 ;
        RECT 4.400 470.880 2246.000 472.280 ;
        RECT 2.365 466.160 2246.000 470.880 ;
        RECT 4.400 464.760 2246.000 466.160 ;
        RECT 2.365 459.360 2246.000 464.760 ;
        RECT 4.400 457.960 2246.000 459.360 ;
        RECT 2.365 452.560 2246.000 457.960 ;
        RECT 4.400 451.160 2246.000 452.560 ;
        RECT 2.365 445.760 2246.000 451.160 ;
        RECT 4.400 444.360 2246.000 445.760 ;
        RECT 2.365 439.640 2246.000 444.360 ;
        RECT 4.400 438.240 2246.000 439.640 ;
        RECT 2.365 432.840 2246.000 438.240 ;
        RECT 4.400 431.440 2246.000 432.840 ;
        RECT 2.365 426.040 2246.000 431.440 ;
        RECT 4.400 424.640 2246.000 426.040 ;
        RECT 2.365 419.920 2246.000 424.640 ;
        RECT 4.400 418.520 2246.000 419.920 ;
        RECT 2.365 413.120 2246.000 418.520 ;
        RECT 4.400 411.720 2246.000 413.120 ;
        RECT 2.365 406.320 2246.000 411.720 ;
        RECT 4.400 404.920 2246.000 406.320 ;
        RECT 2.365 399.520 2246.000 404.920 ;
        RECT 4.400 398.120 2246.000 399.520 ;
        RECT 2.365 393.400 2246.000 398.120 ;
        RECT 4.400 392.000 2246.000 393.400 ;
        RECT 2.365 386.600 2246.000 392.000 ;
        RECT 4.400 385.200 2246.000 386.600 ;
        RECT 2.365 379.800 2246.000 385.200 ;
        RECT 4.400 378.400 2246.000 379.800 ;
        RECT 2.365 373.680 2246.000 378.400 ;
        RECT 4.400 372.280 2246.000 373.680 ;
        RECT 2.365 366.880 2246.000 372.280 ;
        RECT 4.400 365.480 2246.000 366.880 ;
        RECT 2.365 360.080 2246.000 365.480 ;
        RECT 4.400 358.680 2246.000 360.080 ;
        RECT 2.365 353.280 2246.000 358.680 ;
        RECT 4.400 351.880 2246.000 353.280 ;
        RECT 2.365 347.160 2246.000 351.880 ;
        RECT 4.400 345.760 2246.000 347.160 ;
        RECT 2.365 340.360 2246.000 345.760 ;
        RECT 4.400 338.960 2246.000 340.360 ;
        RECT 2.365 333.560 2246.000 338.960 ;
        RECT 4.400 332.160 2246.000 333.560 ;
        RECT 2.365 327.440 2246.000 332.160 ;
        RECT 4.400 326.040 2246.000 327.440 ;
        RECT 2.365 320.640 2246.000 326.040 ;
        RECT 4.400 319.240 2246.000 320.640 ;
        RECT 2.365 313.840 2246.000 319.240 ;
        RECT 4.400 312.440 2246.000 313.840 ;
        RECT 2.365 307.040 2246.000 312.440 ;
        RECT 4.400 305.640 2246.000 307.040 ;
        RECT 2.365 300.920 2246.000 305.640 ;
        RECT 4.400 299.520 2246.000 300.920 ;
        RECT 2.365 294.120 2246.000 299.520 ;
        RECT 4.400 292.720 2246.000 294.120 ;
        RECT 2.365 287.320 2246.000 292.720 ;
        RECT 4.400 285.920 2246.000 287.320 ;
        RECT 2.365 281.200 2246.000 285.920 ;
        RECT 4.400 279.800 2246.000 281.200 ;
        RECT 2.365 274.400 2246.000 279.800 ;
        RECT 4.400 273.000 2246.000 274.400 ;
        RECT 2.365 267.600 2246.000 273.000 ;
        RECT 4.400 266.200 2246.000 267.600 ;
        RECT 2.365 260.800 2246.000 266.200 ;
        RECT 4.400 259.400 2246.000 260.800 ;
        RECT 2.365 254.680 2246.000 259.400 ;
        RECT 4.400 253.280 2246.000 254.680 ;
        RECT 2.365 247.880 2246.000 253.280 ;
        RECT 4.400 246.480 2246.000 247.880 ;
        RECT 2.365 241.080 2246.000 246.480 ;
        RECT 4.400 239.680 2246.000 241.080 ;
        RECT 2.365 234.960 2246.000 239.680 ;
        RECT 4.400 233.560 2246.000 234.960 ;
        RECT 2.365 228.160 2246.000 233.560 ;
        RECT 4.400 226.760 2246.000 228.160 ;
        RECT 2.365 221.360 2246.000 226.760 ;
        RECT 4.400 219.960 2246.000 221.360 ;
        RECT 2.365 214.560 2246.000 219.960 ;
        RECT 4.400 213.160 2246.000 214.560 ;
        RECT 2.365 208.440 2246.000 213.160 ;
        RECT 4.400 207.040 2246.000 208.440 ;
        RECT 2.365 201.640 2246.000 207.040 ;
        RECT 4.400 200.240 2246.000 201.640 ;
        RECT 2.365 194.840 2246.000 200.240 ;
        RECT 4.400 193.440 2246.000 194.840 ;
        RECT 2.365 188.720 2246.000 193.440 ;
        RECT 4.400 187.320 2246.000 188.720 ;
        RECT 2.365 186.000 2246.000 187.320 ;
        RECT 2.365 184.600 2245.600 186.000 ;
        RECT 2.365 181.920 2246.000 184.600 ;
        RECT 4.400 180.520 2246.000 181.920 ;
        RECT 2.365 175.120 2246.000 180.520 ;
        RECT 4.400 173.720 2246.000 175.120 ;
        RECT 2.365 168.320 2246.000 173.720 ;
        RECT 4.400 166.920 2246.000 168.320 ;
        RECT 2.365 162.200 2246.000 166.920 ;
        RECT 4.400 160.800 2246.000 162.200 ;
        RECT 2.365 155.400 2246.000 160.800 ;
        RECT 4.400 154.000 2246.000 155.400 ;
        RECT 2.365 148.600 2246.000 154.000 ;
        RECT 4.400 147.200 2246.000 148.600 ;
        RECT 2.365 142.480 2246.000 147.200 ;
        RECT 4.400 141.080 2246.000 142.480 ;
        RECT 2.365 135.680 2246.000 141.080 ;
        RECT 4.400 134.280 2246.000 135.680 ;
        RECT 2.365 128.880 2246.000 134.280 ;
        RECT 4.400 127.480 2246.000 128.880 ;
        RECT 2.365 122.080 2246.000 127.480 ;
        RECT 4.400 120.680 2246.000 122.080 ;
        RECT 2.365 115.960 2246.000 120.680 ;
        RECT 4.400 114.560 2246.000 115.960 ;
        RECT 2.365 109.160 2246.000 114.560 ;
        RECT 4.400 107.760 2246.000 109.160 ;
        RECT 2.365 102.360 2246.000 107.760 ;
        RECT 4.400 100.960 2246.000 102.360 ;
        RECT 2.365 96.240 2246.000 100.960 ;
        RECT 4.400 94.840 2246.000 96.240 ;
        RECT 2.365 89.440 2246.000 94.840 ;
        RECT 4.400 88.040 2246.000 89.440 ;
        RECT 2.365 82.640 2246.000 88.040 ;
        RECT 4.400 81.240 2246.000 82.640 ;
        RECT 2.365 75.840 2246.000 81.240 ;
        RECT 4.400 74.440 2246.000 75.840 ;
        RECT 2.365 69.720 2246.000 74.440 ;
        RECT 4.400 68.320 2246.000 69.720 ;
        RECT 2.365 62.920 2246.000 68.320 ;
        RECT 4.400 61.520 2246.000 62.920 ;
        RECT 2.365 56.120 2246.000 61.520 ;
        RECT 4.400 54.720 2246.000 56.120 ;
        RECT 2.365 50.000 2246.000 54.720 ;
        RECT 4.400 48.600 2246.000 50.000 ;
        RECT 2.365 43.200 2246.000 48.600 ;
        RECT 4.400 41.800 2246.000 43.200 ;
        RECT 2.365 36.400 2246.000 41.800 ;
        RECT 4.400 35.000 2246.000 36.400 ;
        RECT 2.365 29.600 2246.000 35.000 ;
        RECT 4.400 28.200 2246.000 29.600 ;
        RECT 2.365 23.480 2246.000 28.200 ;
        RECT 4.400 22.080 2246.000 23.480 ;
        RECT 2.365 16.680 2246.000 22.080 ;
        RECT 4.400 15.280 2246.000 16.680 ;
        RECT 2.365 9.880 2246.000 15.280 ;
        RECT 4.400 8.480 2246.000 9.880 ;
        RECT 2.365 3.760 2246.000 8.480 ;
        RECT 4.400 2.360 2246.000 3.760 ;
        RECT 2.365 0.860 2246.000 2.360 ;
      LAYER met4 ;
        RECT 12.750 729.600 2224.690 734.905 ;
        RECT 12.750 10.240 20.640 729.600 ;
        RECT 23.040 10.240 45.640 729.600 ;
        RECT 48.040 10.240 70.640 729.600 ;
        RECT 73.040 517.860 95.640 729.600 ;
        RECT 98.040 517.860 120.640 729.600 ;
        RECT 123.040 517.860 145.640 729.600 ;
        RECT 148.040 517.860 170.640 729.600 ;
        RECT 173.040 517.860 195.640 729.600 ;
        RECT 198.040 517.860 220.640 729.600 ;
        RECT 223.040 517.860 245.640 729.600 ;
        RECT 248.040 517.860 270.640 729.600 ;
        RECT 273.040 517.860 295.640 729.600 ;
        RECT 298.040 517.860 320.640 729.600 ;
        RECT 323.040 517.860 345.640 729.600 ;
        RECT 348.040 517.860 370.640 729.600 ;
        RECT 373.040 517.860 395.640 729.600 ;
        RECT 398.040 517.860 420.640 729.600 ;
        RECT 423.040 517.860 445.640 729.600 ;
        RECT 448.040 517.860 470.640 729.600 ;
        RECT 473.040 517.860 495.640 729.600 ;
        RECT 498.040 517.860 520.640 729.600 ;
        RECT 523.040 517.860 545.640 729.600 ;
        RECT 548.040 517.860 570.640 729.600 ;
        RECT 573.040 517.860 595.640 729.600 ;
        RECT 73.040 101.640 595.640 517.860 ;
        RECT 73.040 10.240 95.640 101.640 ;
        RECT 98.040 10.240 120.640 101.640 ;
        RECT 123.040 10.240 145.640 101.640 ;
        RECT 148.040 10.240 170.640 101.640 ;
        RECT 173.040 10.240 195.640 101.640 ;
        RECT 198.040 10.240 220.640 101.640 ;
        RECT 223.040 10.240 245.640 101.640 ;
        RECT 248.040 10.240 270.640 101.640 ;
        RECT 273.040 10.240 295.640 101.640 ;
        RECT 298.040 10.240 320.640 101.640 ;
        RECT 323.040 10.240 345.640 101.640 ;
        RECT 348.040 10.240 370.640 101.640 ;
        RECT 373.040 10.240 395.640 101.640 ;
        RECT 398.040 10.240 420.640 101.640 ;
        RECT 423.040 10.240 445.640 101.640 ;
        RECT 448.040 10.240 470.640 101.640 ;
        RECT 473.040 10.240 495.640 101.640 ;
        RECT 498.040 10.240 520.640 101.640 ;
        RECT 523.040 10.240 545.640 101.640 ;
        RECT 548.040 10.240 570.640 101.640 ;
        RECT 573.040 10.240 595.640 101.640 ;
        RECT 598.040 10.240 620.640 729.600 ;
        RECT 623.040 10.240 645.640 729.600 ;
        RECT 648.040 517.860 670.640 729.600 ;
        RECT 673.040 517.860 695.640 729.600 ;
        RECT 698.040 517.860 720.640 729.600 ;
        RECT 723.040 517.860 745.640 729.600 ;
        RECT 748.040 517.860 770.640 729.600 ;
        RECT 773.040 517.860 795.640 729.600 ;
        RECT 798.040 517.860 820.640 729.600 ;
        RECT 823.040 517.860 845.640 729.600 ;
        RECT 848.040 517.860 870.640 729.600 ;
        RECT 873.040 517.860 895.640 729.600 ;
        RECT 898.040 517.860 920.640 729.600 ;
        RECT 923.040 517.860 945.640 729.600 ;
        RECT 948.040 517.860 970.640 729.600 ;
        RECT 973.040 517.860 995.640 729.600 ;
        RECT 998.040 517.860 1020.640 729.600 ;
        RECT 1023.040 517.860 1045.640 729.600 ;
        RECT 1048.040 517.860 1070.640 729.600 ;
        RECT 1073.040 517.860 1095.640 729.600 ;
        RECT 1098.040 517.860 1120.640 729.600 ;
        RECT 1123.040 517.860 1145.640 729.600 ;
        RECT 1148.040 517.860 1170.640 729.600 ;
        RECT 648.040 101.640 1170.640 517.860 ;
        RECT 648.040 10.240 670.640 101.640 ;
        RECT 673.040 10.240 695.640 101.640 ;
        RECT 698.040 10.240 720.640 101.640 ;
        RECT 723.040 10.240 745.640 101.640 ;
        RECT 748.040 10.240 770.640 101.640 ;
        RECT 773.040 10.240 795.640 101.640 ;
        RECT 798.040 10.240 820.640 101.640 ;
        RECT 823.040 10.240 845.640 101.640 ;
        RECT 848.040 10.240 870.640 101.640 ;
        RECT 873.040 10.240 895.640 101.640 ;
        RECT 898.040 10.240 920.640 101.640 ;
        RECT 923.040 10.240 945.640 101.640 ;
        RECT 948.040 10.240 970.640 101.640 ;
        RECT 973.040 10.240 995.640 101.640 ;
        RECT 998.040 10.240 1020.640 101.640 ;
        RECT 1023.040 10.240 1045.640 101.640 ;
        RECT 1048.040 10.240 1070.640 101.640 ;
        RECT 1073.040 10.240 1095.640 101.640 ;
        RECT 1098.040 10.240 1120.640 101.640 ;
        RECT 1123.040 10.240 1145.640 101.640 ;
        RECT 1148.040 10.240 1170.640 101.640 ;
        RECT 1173.040 10.240 1195.640 729.600 ;
        RECT 1198.040 10.240 1220.640 729.600 ;
        RECT 1223.040 10.240 1245.640 729.600 ;
        RECT 1248.040 10.240 1270.640 729.600 ;
        RECT 1273.040 10.240 1295.640 729.600 ;
        RECT 1298.040 10.240 1320.640 729.600 ;
        RECT 1323.040 10.240 1345.640 729.600 ;
        RECT 1348.040 10.240 1370.640 729.600 ;
        RECT 1373.040 10.240 1395.640 729.600 ;
        RECT 1398.040 10.240 1420.640 729.600 ;
        RECT 1423.040 10.240 1445.640 729.600 ;
        RECT 1448.040 10.240 1470.640 729.600 ;
        RECT 1473.040 10.240 1495.640 729.600 ;
        RECT 1498.040 10.240 1520.640 729.600 ;
        RECT 1523.040 10.240 1545.640 729.600 ;
        RECT 1548.040 10.240 1570.640 729.600 ;
        RECT 1573.040 10.240 1595.640 729.600 ;
        RECT 1598.040 10.240 1620.640 729.600 ;
        RECT 1623.040 10.240 1645.640 729.600 ;
        RECT 1648.040 10.240 1670.640 729.600 ;
        RECT 1673.040 10.240 1695.640 729.600 ;
        RECT 1698.040 10.240 1720.640 729.600 ;
        RECT 1723.040 10.240 1745.640 729.600 ;
        RECT 1748.040 10.240 1770.640 729.600 ;
        RECT 1773.040 10.240 1795.640 729.600 ;
        RECT 1798.040 10.240 1820.640 729.600 ;
        RECT 1823.040 10.240 1845.640 729.600 ;
        RECT 1848.040 10.240 1870.640 729.600 ;
        RECT 1873.040 10.240 1895.640 729.600 ;
        RECT 1898.040 10.240 1920.640 729.600 ;
        RECT 1923.040 10.240 1945.640 729.600 ;
        RECT 1948.040 10.240 1970.640 729.600 ;
        RECT 1973.040 10.240 1995.640 729.600 ;
        RECT 1998.040 10.240 2020.640 729.600 ;
        RECT 2023.040 10.240 2045.640 729.600 ;
        RECT 2048.040 10.240 2070.640 729.600 ;
        RECT 2073.040 10.240 2095.640 729.600 ;
        RECT 2098.040 10.240 2120.640 729.600 ;
        RECT 2123.040 10.240 2145.640 729.600 ;
        RECT 2148.040 10.240 2170.640 729.600 ;
        RECT 2173.040 10.240 2195.640 729.600 ;
        RECT 2198.040 10.240 2220.640 729.600 ;
        RECT 2223.040 10.240 2224.690 729.600 ;
        RECT 12.750 0.855 2224.690 10.240 ;
      LAYER met5 ;
        RECT 12.540 679.690 2224.900 726.700 ;
        RECT 12.540 614.690 2224.900 674.890 ;
        RECT 12.540 549.690 2224.900 609.890 ;
        RECT 12.540 484.690 2224.900 544.890 ;
        RECT 12.540 419.690 2224.900 479.890 ;
        RECT 12.540 354.690 2224.900 414.890 ;
        RECT 12.540 289.690 2224.900 349.890 ;
        RECT 12.540 224.690 2224.900 284.890 ;
        RECT 12.540 159.690 2224.900 219.890 ;
        RECT 12.540 94.690 2224.900 154.890 ;
        RECT 12.540 29.690 2224.900 89.890 ;
        RECT 12.540 11.100 2224.900 24.890 ;
  END
END mgmt_core
END LIBRARY

