magic
tech sky130A
magscale 1 2
timestamp 1636710988
<< obsli1 >>
rect 5869 4641 539551 163931
<< obsm1 >>
rect 382 1300 539566 163996
<< metal2 >>
rect 386 163200 442 164000
rect 1214 163200 1270 164000
rect 2042 163200 2098 164000
rect 2962 163200 3018 164000
rect 3790 163200 3846 164000
rect 4710 163200 4766 164000
rect 5538 163200 5594 164000
rect 6366 163200 6422 164000
rect 7286 163200 7342 164000
rect 8114 163200 8170 164000
rect 9034 163200 9090 164000
rect 9862 163200 9918 164000
rect 10782 163200 10838 164000
rect 11610 163200 11666 164000
rect 12438 163200 12494 164000
rect 13358 163200 13414 164000
rect 14186 163200 14242 164000
rect 15106 163200 15162 164000
rect 15934 163200 15990 164000
rect 16854 163200 16910 164000
rect 17682 163200 17738 164000
rect 18510 163200 18566 164000
rect 19430 163200 19486 164000
rect 20258 163200 20314 164000
rect 21178 163200 21234 164000
rect 22006 163200 22062 164000
rect 22834 163200 22890 164000
rect 23754 163200 23810 164000
rect 24582 163200 24638 164000
rect 25502 163200 25558 164000
rect 26330 163200 26386 164000
rect 27250 163200 27306 164000
rect 28078 163200 28134 164000
rect 28906 163200 28962 164000
rect 29826 163200 29882 164000
rect 30654 163200 30710 164000
rect 31574 163200 31630 164000
rect 32402 163200 32458 164000
rect 33322 163200 33378 164000
rect 34150 163200 34206 164000
rect 34978 163200 35034 164000
rect 35898 163200 35954 164000
rect 36726 163200 36782 164000
rect 37646 163200 37702 164000
rect 38474 163200 38530 164000
rect 39302 163200 39358 164000
rect 40222 163200 40278 164000
rect 41050 163200 41106 164000
rect 41970 163200 42026 164000
rect 42798 163200 42854 164000
rect 43718 163200 43774 164000
rect 44546 163200 44602 164000
rect 45374 163200 45430 164000
rect 46294 163200 46350 164000
rect 47122 163200 47178 164000
rect 48042 163200 48098 164000
rect 48870 163200 48926 164000
rect 49790 163200 49846 164000
rect 50618 163200 50674 164000
rect 51446 163200 51502 164000
rect 52366 163200 52422 164000
rect 53194 163200 53250 164000
rect 54114 163200 54170 164000
rect 54942 163200 54998 164000
rect 55862 163200 55918 164000
rect 56690 163200 56746 164000
rect 57518 163200 57574 164000
rect 58438 163200 58494 164000
rect 59266 163200 59322 164000
rect 60186 163200 60242 164000
rect 61014 163200 61070 164000
rect 61842 163200 61898 164000
rect 62762 163200 62818 164000
rect 63590 163200 63646 164000
rect 64510 163200 64566 164000
rect 65338 163200 65394 164000
rect 66258 163200 66314 164000
rect 67086 163200 67142 164000
rect 67914 163200 67970 164000
rect 68834 163200 68890 164000
rect 69662 163200 69718 164000
rect 70582 163200 70638 164000
rect 71410 163200 71466 164000
rect 72330 163200 72386 164000
rect 73158 163200 73214 164000
rect 73986 163200 74042 164000
rect 74906 163200 74962 164000
rect 75734 163200 75790 164000
rect 76654 163200 76710 164000
rect 77482 163200 77538 164000
rect 78310 163200 78366 164000
rect 79230 163200 79286 164000
rect 80058 163200 80114 164000
rect 80978 163200 81034 164000
rect 81806 163200 81862 164000
rect 82726 163200 82782 164000
rect 83554 163200 83610 164000
rect 84382 163200 84438 164000
rect 85302 163200 85358 164000
rect 86130 163200 86186 164000
rect 87050 163200 87106 164000
rect 87878 163200 87934 164000
rect 88798 163200 88854 164000
rect 89626 163200 89682 164000
rect 90454 163200 90510 164000
rect 91374 163200 91430 164000
rect 92202 163200 92258 164000
rect 93122 163200 93178 164000
rect 93950 163200 94006 164000
rect 94870 163200 94926 164000
rect 95698 163200 95754 164000
rect 96526 163200 96582 164000
rect 97446 163200 97502 164000
rect 98274 163200 98330 164000
rect 99194 163200 99250 164000
rect 100022 163200 100078 164000
rect 100850 163200 100906 164000
rect 101770 163200 101826 164000
rect 102598 163200 102654 164000
rect 103518 163200 103574 164000
rect 104346 163200 104402 164000
rect 105266 163200 105322 164000
rect 106094 163200 106150 164000
rect 106922 163200 106978 164000
rect 107842 163200 107898 164000
rect 108670 163200 108726 164000
rect 109590 163200 109646 164000
rect 110418 163200 110474 164000
rect 111338 163200 111394 164000
rect 112166 163200 112222 164000
rect 112994 163200 113050 164000
rect 113914 163200 113970 164000
rect 114742 163200 114798 164000
rect 115662 163200 115718 164000
rect 116490 163200 116546 164000
rect 117318 163200 117374 164000
rect 118238 163200 118294 164000
rect 119066 163200 119122 164000
rect 119986 163200 120042 164000
rect 120814 163200 120870 164000
rect 121734 163200 121790 164000
rect 122562 163200 122618 164000
rect 123390 163200 123446 164000
rect 124310 163200 124366 164000
rect 125138 163200 125194 164000
rect 126058 163200 126114 164000
rect 126886 163200 126942 164000
rect 127806 163200 127862 164000
rect 128634 163200 128690 164000
rect 129462 163200 129518 164000
rect 130382 163200 130438 164000
rect 131210 163200 131266 164000
rect 132130 163200 132186 164000
rect 132958 163200 133014 164000
rect 133878 163200 133934 164000
rect 134706 163200 134762 164000
rect 135534 163200 135590 164000
rect 136454 163200 136510 164000
rect 137282 163200 137338 164000
rect 138202 163200 138258 164000
rect 139030 163200 139086 164000
rect 139858 163200 139914 164000
rect 140778 163200 140834 164000
rect 141606 163200 141662 164000
rect 142526 163200 142582 164000
rect 143354 163200 143410 164000
rect 144274 163200 144330 164000
rect 145102 163200 145158 164000
rect 145930 163200 145986 164000
rect 146850 163200 146906 164000
rect 147678 163200 147734 164000
rect 148598 163200 148654 164000
rect 149426 163200 149482 164000
rect 150346 163200 150402 164000
rect 151174 163200 151230 164000
rect 152002 163200 152058 164000
rect 152922 163200 152978 164000
rect 153750 163200 153806 164000
rect 154670 163200 154726 164000
rect 155498 163200 155554 164000
rect 156326 163200 156382 164000
rect 157246 163200 157302 164000
rect 158074 163200 158130 164000
rect 158994 163200 159050 164000
rect 159822 163200 159878 164000
rect 160742 163200 160798 164000
rect 161570 163200 161626 164000
rect 162398 163200 162454 164000
rect 163318 163200 163374 164000
rect 164146 163200 164202 164000
rect 165066 163200 165122 164000
rect 165894 163200 165950 164000
rect 166814 163200 166870 164000
rect 167642 163200 167698 164000
rect 168470 163200 168526 164000
rect 169390 163200 169446 164000
rect 170218 163200 170274 164000
rect 171138 163200 171194 164000
rect 171966 163200 172022 164000
rect 172886 163200 172942 164000
rect 173714 163200 173770 164000
rect 174542 163200 174598 164000
rect 175462 163200 175518 164000
rect 176290 163200 176346 164000
rect 177210 163200 177266 164000
rect 178038 163200 178094 164000
rect 178866 163200 178922 164000
rect 179786 163200 179842 164000
rect 180614 163200 180670 164000
rect 181534 163200 181590 164000
rect 182362 163200 182418 164000
rect 183282 163200 183338 164000
rect 184110 163200 184166 164000
rect 184938 163200 184994 164000
rect 185858 163200 185914 164000
rect 186686 163200 186742 164000
rect 187606 163200 187662 164000
rect 188434 163200 188490 164000
rect 189354 163200 189410 164000
rect 190182 163200 190238 164000
rect 191010 163200 191066 164000
rect 191930 163200 191986 164000
rect 192758 163200 192814 164000
rect 193678 163200 193734 164000
rect 194506 163200 194562 164000
rect 195334 163200 195390 164000
rect 196254 163200 196310 164000
rect 197082 163200 197138 164000
rect 198002 163200 198058 164000
rect 198830 163200 198886 164000
rect 199750 163200 199806 164000
rect 200578 163200 200634 164000
rect 201406 163200 201462 164000
rect 202326 163200 202382 164000
rect 203154 163200 203210 164000
rect 204074 163200 204130 164000
rect 204902 163200 204958 164000
rect 205822 163200 205878 164000
rect 206650 163200 206706 164000
rect 207478 163200 207534 164000
rect 208398 163200 208454 164000
rect 209226 163200 209282 164000
rect 210146 163200 210202 164000
rect 210974 163200 211030 164000
rect 211894 163200 211950 164000
rect 212722 163200 212778 164000
rect 213550 163200 213606 164000
rect 214470 163200 214526 164000
rect 215298 163200 215354 164000
rect 216218 163200 216274 164000
rect 217046 163200 217102 164000
rect 217874 163200 217930 164000
rect 218794 163200 218850 164000
rect 219622 163200 219678 164000
rect 220542 163200 220598 164000
rect 221370 163200 221426 164000
rect 222290 163200 222346 164000
rect 223118 163200 223174 164000
rect 223946 163200 224002 164000
rect 224866 163200 224922 164000
rect 225694 163200 225750 164000
rect 226614 163200 226670 164000
rect 227442 163200 227498 164000
rect 228362 163200 228418 164000
rect 229190 163200 229246 164000
rect 230018 163200 230074 164000
rect 230938 163200 230994 164000
rect 231766 163200 231822 164000
rect 232686 163200 232742 164000
rect 233514 163200 233570 164000
rect 234342 163200 234398 164000
rect 235262 163200 235318 164000
rect 236090 163200 236146 164000
rect 237010 163200 237066 164000
rect 237838 163200 237894 164000
rect 238758 163200 238814 164000
rect 239586 163200 239642 164000
rect 240414 163200 240470 164000
rect 241334 163200 241390 164000
rect 242162 163200 242218 164000
rect 243082 163200 243138 164000
rect 243910 163200 243966 164000
rect 244830 163200 244886 164000
rect 245658 163200 245714 164000
rect 246486 163200 246542 164000
rect 247406 163200 247462 164000
rect 248234 163200 248290 164000
rect 249154 163200 249210 164000
rect 249982 163200 250038 164000
rect 250902 163200 250958 164000
rect 251730 163200 251786 164000
rect 252558 163200 252614 164000
rect 253478 163200 253534 164000
rect 254306 163200 254362 164000
rect 255226 163200 255282 164000
rect 256054 163200 256110 164000
rect 256882 163200 256938 164000
rect 257802 163200 257858 164000
rect 258630 163200 258686 164000
rect 259550 163200 259606 164000
rect 260378 163200 260434 164000
rect 261298 163200 261354 164000
rect 262126 163200 262182 164000
rect 262954 163200 263010 164000
rect 263874 163200 263930 164000
rect 264702 163200 264758 164000
rect 265622 163200 265678 164000
rect 266450 163200 266506 164000
rect 267370 163200 267426 164000
rect 268198 163200 268254 164000
rect 269026 163200 269082 164000
rect 269946 163200 270002 164000
rect 270774 163200 270830 164000
rect 271694 163200 271750 164000
rect 272522 163200 272578 164000
rect 273350 163200 273406 164000
rect 274270 163200 274326 164000
rect 275098 163200 275154 164000
rect 276018 163200 276074 164000
rect 276846 163200 276902 164000
rect 277766 163200 277822 164000
rect 278594 163200 278650 164000
rect 279422 163200 279478 164000
rect 280342 163200 280398 164000
rect 281170 163200 281226 164000
rect 282090 163200 282146 164000
rect 282918 163200 282974 164000
rect 283838 163200 283894 164000
rect 284666 163200 284722 164000
rect 285494 163200 285550 164000
rect 286414 163200 286470 164000
rect 287242 163200 287298 164000
rect 288162 163200 288218 164000
rect 288990 163200 289046 164000
rect 289818 163200 289874 164000
rect 290738 163200 290794 164000
rect 291566 163200 291622 164000
rect 292486 163200 292542 164000
rect 293314 163200 293370 164000
rect 294234 163200 294290 164000
rect 295062 163200 295118 164000
rect 295890 163200 295946 164000
rect 296810 163200 296866 164000
rect 297638 163200 297694 164000
rect 298558 163200 298614 164000
rect 299386 163200 299442 164000
rect 300306 163200 300362 164000
rect 301134 163200 301190 164000
rect 301962 163200 302018 164000
rect 302882 163200 302938 164000
rect 303710 163200 303766 164000
rect 304630 163200 304686 164000
rect 305458 163200 305514 164000
rect 306378 163200 306434 164000
rect 307206 163200 307262 164000
rect 308034 163200 308090 164000
rect 308954 163200 309010 164000
rect 309782 163200 309838 164000
rect 310702 163200 310758 164000
rect 311530 163200 311586 164000
rect 312358 163200 312414 164000
rect 313278 163200 313334 164000
rect 314106 163200 314162 164000
rect 315026 163200 315082 164000
rect 315854 163200 315910 164000
rect 316774 163200 316830 164000
rect 317602 163200 317658 164000
rect 318430 163200 318486 164000
rect 319350 163200 319406 164000
rect 320178 163200 320234 164000
rect 321098 163200 321154 164000
rect 321926 163200 321982 164000
rect 322846 163200 322902 164000
rect 323674 163200 323730 164000
rect 324502 163200 324558 164000
rect 325422 163200 325478 164000
rect 326250 163200 326306 164000
rect 327170 163200 327226 164000
rect 327998 163200 328054 164000
rect 328826 163200 328882 164000
rect 329746 163200 329802 164000
rect 330574 163200 330630 164000
rect 331494 163200 331550 164000
rect 332322 163200 332378 164000
rect 333242 163200 333298 164000
rect 334070 163200 334126 164000
rect 334898 163200 334954 164000
rect 335818 163200 335874 164000
rect 336646 163200 336702 164000
rect 337566 163200 337622 164000
rect 338394 163200 338450 164000
rect 339314 163200 339370 164000
rect 340142 163200 340198 164000
rect 340970 163200 341026 164000
rect 341890 163200 341946 164000
rect 342718 163200 342774 164000
rect 343638 163200 343694 164000
rect 344466 163200 344522 164000
rect 345386 163200 345442 164000
rect 346214 163200 346270 164000
rect 347042 163200 347098 164000
rect 347962 163200 348018 164000
rect 348790 163200 348846 164000
rect 349710 163200 349766 164000
rect 350538 163200 350594 164000
rect 351366 163200 351422 164000
rect 352286 163200 352342 164000
rect 353114 163200 353170 164000
rect 354034 163200 354090 164000
rect 354862 163200 354918 164000
rect 355782 163200 355838 164000
rect 356610 163200 356666 164000
rect 357438 163200 357494 164000
rect 358358 163200 358414 164000
rect 359186 163200 359242 164000
rect 360106 163200 360162 164000
rect 360934 163200 360990 164000
rect 361854 163200 361910 164000
rect 362682 163200 362738 164000
rect 363510 163200 363566 164000
rect 364430 163200 364486 164000
rect 365258 163200 365314 164000
rect 366178 163200 366234 164000
rect 367006 163200 367062 164000
rect 367834 163200 367890 164000
rect 368754 163200 368810 164000
rect 369582 163200 369638 164000
rect 370502 163200 370558 164000
rect 371330 163200 371386 164000
rect 372250 163200 372306 164000
rect 373078 163200 373134 164000
rect 373906 163200 373962 164000
rect 374826 163200 374882 164000
rect 375654 163200 375710 164000
rect 376574 163200 376630 164000
rect 377402 163200 377458 164000
rect 378322 163200 378378 164000
rect 379150 163200 379206 164000
rect 379978 163200 380034 164000
rect 380898 163200 380954 164000
rect 381726 163200 381782 164000
rect 382646 163200 382702 164000
rect 383474 163200 383530 164000
rect 384394 163200 384450 164000
rect 385222 163200 385278 164000
rect 386050 163200 386106 164000
rect 386970 163200 387026 164000
rect 387798 163200 387854 164000
rect 388718 163200 388774 164000
rect 389546 163200 389602 164000
rect 390374 163200 390430 164000
rect 391294 163200 391350 164000
rect 392122 163200 392178 164000
rect 393042 163200 393098 164000
rect 393870 163200 393926 164000
rect 394790 163200 394846 164000
rect 395618 163200 395674 164000
rect 396446 163200 396502 164000
rect 397366 163200 397422 164000
rect 398194 163200 398250 164000
rect 399114 163200 399170 164000
rect 399942 163200 399998 164000
rect 400862 163200 400918 164000
rect 401690 163200 401746 164000
rect 402518 163200 402574 164000
rect 403438 163200 403494 164000
rect 404266 163200 404322 164000
rect 405186 163200 405242 164000
rect 406014 163200 406070 164000
rect 406842 163200 406898 164000
rect 407762 163200 407818 164000
rect 408590 163200 408646 164000
rect 409510 163200 409566 164000
rect 410338 163200 410394 164000
rect 411258 163200 411314 164000
rect 412086 163200 412142 164000
rect 412914 163200 412970 164000
rect 413834 163200 413890 164000
rect 414662 163200 414718 164000
rect 415582 163200 415638 164000
rect 416410 163200 416466 164000
rect 417330 163200 417386 164000
rect 418158 163200 418214 164000
rect 418986 163200 419042 164000
rect 419906 163200 419962 164000
rect 420734 163200 420790 164000
rect 421654 163200 421710 164000
rect 422482 163200 422538 164000
rect 423402 163200 423458 164000
rect 424230 163200 424286 164000
rect 425058 163200 425114 164000
rect 425978 163200 426034 164000
rect 426806 163200 426862 164000
rect 427726 163200 427782 164000
rect 428554 163200 428610 164000
rect 429382 163200 429438 164000
rect 430302 163200 430358 164000
rect 431130 163200 431186 164000
rect 432050 163200 432106 164000
rect 432878 163200 432934 164000
rect 433798 163200 433854 164000
rect 434626 163200 434682 164000
rect 435454 163200 435510 164000
rect 436374 163200 436430 164000
rect 437202 163200 437258 164000
rect 438122 163200 438178 164000
rect 438950 163200 439006 164000
rect 439870 163200 439926 164000
rect 440698 163200 440754 164000
rect 441526 163200 441582 164000
rect 442446 163200 442502 164000
rect 443274 163200 443330 164000
rect 444194 163200 444250 164000
rect 445022 163200 445078 164000
rect 445850 163200 445906 164000
rect 446770 163200 446826 164000
rect 447598 163200 447654 164000
rect 448518 163200 448574 164000
rect 449346 163200 449402 164000
rect 450266 163200 450322 164000
rect 451094 163200 451150 164000
rect 451922 163200 451978 164000
rect 452842 163200 452898 164000
rect 453670 163200 453726 164000
rect 454590 163200 454646 164000
rect 455418 163200 455474 164000
rect 456338 163200 456394 164000
rect 457166 163200 457222 164000
rect 457994 163200 458050 164000
rect 458914 163200 458970 164000
rect 459742 163200 459798 164000
rect 460662 163200 460718 164000
rect 461490 163200 461546 164000
rect 462410 163200 462466 164000
rect 463238 163200 463294 164000
rect 464066 163200 464122 164000
rect 464986 163200 465042 164000
rect 465814 163200 465870 164000
rect 466734 163200 466790 164000
rect 467562 163200 467618 164000
rect 468390 163200 468446 164000
rect 469310 163200 469366 164000
rect 470138 163200 470194 164000
rect 471058 163200 471114 164000
rect 471886 163200 471942 164000
rect 472806 163200 472862 164000
rect 473634 163200 473690 164000
rect 474462 163200 474518 164000
rect 475382 163200 475438 164000
rect 476210 163200 476266 164000
rect 477130 163200 477186 164000
rect 477958 163200 478014 164000
rect 478878 163200 478934 164000
rect 479706 163200 479762 164000
rect 480534 163200 480590 164000
rect 481454 163200 481510 164000
rect 482282 163200 482338 164000
rect 483202 163200 483258 164000
rect 484030 163200 484086 164000
rect 484858 163200 484914 164000
rect 485778 163200 485834 164000
rect 486606 163200 486662 164000
rect 487526 163200 487582 164000
rect 488354 163200 488410 164000
rect 489274 163200 489330 164000
rect 490102 163200 490158 164000
rect 490930 163200 490986 164000
rect 491850 163200 491906 164000
rect 492678 163200 492734 164000
rect 493598 163200 493654 164000
rect 494426 163200 494482 164000
rect 495346 163200 495402 164000
rect 496174 163200 496230 164000
rect 497002 163200 497058 164000
rect 497922 163200 497978 164000
rect 498750 163200 498806 164000
rect 499670 163200 499726 164000
rect 500498 163200 500554 164000
rect 501418 163200 501474 164000
rect 502246 163200 502302 164000
rect 503074 163200 503130 164000
rect 503994 163200 504050 164000
rect 504822 163200 504878 164000
rect 505742 163200 505798 164000
rect 506570 163200 506626 164000
rect 507398 163200 507454 164000
rect 508318 163200 508374 164000
rect 509146 163200 509202 164000
rect 510066 163200 510122 164000
rect 510894 163200 510950 164000
rect 511814 163200 511870 164000
rect 512642 163200 512698 164000
rect 513470 163200 513526 164000
rect 514390 163200 514446 164000
rect 515218 163200 515274 164000
rect 516138 163200 516194 164000
rect 516966 163200 517022 164000
rect 517886 163200 517942 164000
rect 518714 163200 518770 164000
rect 519542 163200 519598 164000
rect 520462 163200 520518 164000
rect 521290 163200 521346 164000
rect 522210 163200 522266 164000
rect 523038 163200 523094 164000
rect 523866 163200 523922 164000
rect 524786 163200 524842 164000
rect 525614 163200 525670 164000
rect 526534 163200 526590 164000
rect 527362 163200 527418 164000
rect 528282 163200 528338 164000
rect 529110 163200 529166 164000
rect 529938 163200 529994 164000
rect 530858 163200 530914 164000
rect 531686 163200 531742 164000
rect 532606 163200 532662 164000
rect 533434 163200 533490 164000
rect 534354 163200 534410 164000
rect 535182 163200 535238 164000
rect 536010 163200 536066 164000
rect 536930 163200 536986 164000
rect 537758 163200 537814 164000
rect 538678 163200 538734 164000
rect 539506 163200 539562 164000
rect 33690 0 33746 800
rect 101126 0 101182 800
rect 168654 0 168710 800
rect 236182 0 236238 800
rect 303710 0 303766 800
rect 371146 0 371202 800
rect 438674 0 438730 800
rect 506202 0 506258 800
<< obsm2 >>
rect 498 163144 1158 163946
rect 1326 163144 1986 163946
rect 2154 163144 2906 163946
rect 3074 163144 3734 163946
rect 3902 163144 4654 163946
rect 4822 163144 5482 163946
rect 5650 163144 6310 163946
rect 6478 163144 7230 163946
rect 7398 163144 8058 163946
rect 8226 163144 8978 163946
rect 9146 163144 9806 163946
rect 9974 163144 10726 163946
rect 10894 163144 11554 163946
rect 11722 163144 12382 163946
rect 12550 163144 13302 163946
rect 13470 163144 14130 163946
rect 14298 163144 15050 163946
rect 15218 163144 15878 163946
rect 16046 163144 16798 163946
rect 16966 163144 17626 163946
rect 17794 163144 18454 163946
rect 18622 163144 19374 163946
rect 19542 163144 20202 163946
rect 20370 163144 21122 163946
rect 21290 163144 21950 163946
rect 22118 163144 22778 163946
rect 22946 163144 23698 163946
rect 23866 163144 24526 163946
rect 24694 163144 25446 163946
rect 25614 163144 26274 163946
rect 26442 163144 27194 163946
rect 27362 163144 28022 163946
rect 28190 163144 28850 163946
rect 29018 163144 29770 163946
rect 29938 163144 30598 163946
rect 30766 163144 31518 163946
rect 31686 163144 32346 163946
rect 32514 163144 33266 163946
rect 33434 163144 34094 163946
rect 34262 163144 34922 163946
rect 35090 163144 35842 163946
rect 36010 163144 36670 163946
rect 36838 163144 37590 163946
rect 37758 163144 38418 163946
rect 38586 163144 39246 163946
rect 39414 163144 40166 163946
rect 40334 163144 40994 163946
rect 41162 163144 41914 163946
rect 42082 163144 42742 163946
rect 42910 163144 43662 163946
rect 43830 163144 44490 163946
rect 44658 163144 45318 163946
rect 45486 163144 46238 163946
rect 46406 163144 47066 163946
rect 47234 163144 47986 163946
rect 48154 163144 48814 163946
rect 48982 163144 49734 163946
rect 49902 163144 50562 163946
rect 50730 163144 51390 163946
rect 51558 163144 52310 163946
rect 52478 163144 53138 163946
rect 53306 163144 54058 163946
rect 54226 163144 54886 163946
rect 55054 163144 55806 163946
rect 55974 163144 56634 163946
rect 56802 163144 57462 163946
rect 57630 163144 58382 163946
rect 58550 163144 59210 163946
rect 59378 163144 60130 163946
rect 60298 163144 60958 163946
rect 61126 163144 61786 163946
rect 61954 163144 62706 163946
rect 62874 163144 63534 163946
rect 63702 163144 64454 163946
rect 64622 163144 65282 163946
rect 65450 163144 66202 163946
rect 66370 163144 67030 163946
rect 67198 163144 67858 163946
rect 68026 163144 68778 163946
rect 68946 163144 69606 163946
rect 69774 163144 70526 163946
rect 70694 163144 71354 163946
rect 71522 163144 72274 163946
rect 72442 163144 73102 163946
rect 73270 163144 73930 163946
rect 74098 163144 74850 163946
rect 75018 163144 75678 163946
rect 75846 163144 76598 163946
rect 76766 163144 77426 163946
rect 77594 163144 78254 163946
rect 78422 163144 79174 163946
rect 79342 163144 80002 163946
rect 80170 163144 80922 163946
rect 81090 163144 81750 163946
rect 81918 163144 82670 163946
rect 82838 163144 83498 163946
rect 83666 163144 84326 163946
rect 84494 163144 85246 163946
rect 85414 163144 86074 163946
rect 86242 163144 86994 163946
rect 87162 163144 87822 163946
rect 87990 163144 88742 163946
rect 88910 163144 89570 163946
rect 89738 163144 90398 163946
rect 90566 163144 91318 163946
rect 91486 163144 92146 163946
rect 92314 163144 93066 163946
rect 93234 163144 93894 163946
rect 94062 163144 94814 163946
rect 94982 163144 95642 163946
rect 95810 163144 96470 163946
rect 96638 163144 97390 163946
rect 97558 163144 98218 163946
rect 98386 163144 99138 163946
rect 99306 163144 99966 163946
rect 100134 163144 100794 163946
rect 100962 163144 101714 163946
rect 101882 163144 102542 163946
rect 102710 163144 103462 163946
rect 103630 163144 104290 163946
rect 104458 163144 105210 163946
rect 105378 163144 106038 163946
rect 106206 163144 106866 163946
rect 107034 163144 107786 163946
rect 107954 163144 108614 163946
rect 108782 163144 109534 163946
rect 109702 163144 110362 163946
rect 110530 163144 111282 163946
rect 111450 163144 112110 163946
rect 112278 163144 112938 163946
rect 113106 163144 113858 163946
rect 114026 163144 114686 163946
rect 114854 163144 115606 163946
rect 115774 163144 116434 163946
rect 116602 163144 117262 163946
rect 117430 163144 118182 163946
rect 118350 163144 119010 163946
rect 119178 163144 119930 163946
rect 120098 163144 120758 163946
rect 120926 163144 121678 163946
rect 121846 163144 122506 163946
rect 122674 163144 123334 163946
rect 123502 163144 124254 163946
rect 124422 163144 125082 163946
rect 125250 163144 126002 163946
rect 126170 163144 126830 163946
rect 126998 163144 127750 163946
rect 127918 163144 128578 163946
rect 128746 163144 129406 163946
rect 129574 163144 130326 163946
rect 130494 163144 131154 163946
rect 131322 163144 132074 163946
rect 132242 163144 132902 163946
rect 133070 163144 133822 163946
rect 133990 163144 134650 163946
rect 134818 163144 135478 163946
rect 135646 163144 136398 163946
rect 136566 163144 137226 163946
rect 137394 163144 138146 163946
rect 138314 163144 138974 163946
rect 139142 163144 139802 163946
rect 139970 163144 140722 163946
rect 140890 163144 141550 163946
rect 141718 163144 142470 163946
rect 142638 163144 143298 163946
rect 143466 163144 144218 163946
rect 144386 163144 145046 163946
rect 145214 163144 145874 163946
rect 146042 163144 146794 163946
rect 146962 163144 147622 163946
rect 147790 163144 148542 163946
rect 148710 163144 149370 163946
rect 149538 163144 150290 163946
rect 150458 163144 151118 163946
rect 151286 163144 151946 163946
rect 152114 163144 152866 163946
rect 153034 163144 153694 163946
rect 153862 163144 154614 163946
rect 154782 163144 155442 163946
rect 155610 163144 156270 163946
rect 156438 163144 157190 163946
rect 157358 163144 158018 163946
rect 158186 163144 158938 163946
rect 159106 163144 159766 163946
rect 159934 163144 160686 163946
rect 160854 163144 161514 163946
rect 161682 163144 162342 163946
rect 162510 163144 163262 163946
rect 163430 163144 164090 163946
rect 164258 163144 165010 163946
rect 165178 163144 165838 163946
rect 166006 163144 166758 163946
rect 166926 163144 167586 163946
rect 167754 163144 168414 163946
rect 168582 163144 169334 163946
rect 169502 163144 170162 163946
rect 170330 163144 171082 163946
rect 171250 163144 171910 163946
rect 172078 163144 172830 163946
rect 172998 163144 173658 163946
rect 173826 163144 174486 163946
rect 174654 163144 175406 163946
rect 175574 163144 176234 163946
rect 176402 163144 177154 163946
rect 177322 163144 177982 163946
rect 178150 163144 178810 163946
rect 178978 163144 179730 163946
rect 179898 163144 180558 163946
rect 180726 163144 181478 163946
rect 181646 163144 182306 163946
rect 182474 163144 183226 163946
rect 183394 163144 184054 163946
rect 184222 163144 184882 163946
rect 185050 163144 185802 163946
rect 185970 163144 186630 163946
rect 186798 163144 187550 163946
rect 187718 163144 188378 163946
rect 188546 163144 189298 163946
rect 189466 163144 190126 163946
rect 190294 163144 190954 163946
rect 191122 163144 191874 163946
rect 192042 163144 192702 163946
rect 192870 163144 193622 163946
rect 193790 163144 194450 163946
rect 194618 163144 195278 163946
rect 195446 163144 196198 163946
rect 196366 163144 197026 163946
rect 197194 163144 197946 163946
rect 198114 163144 198774 163946
rect 198942 163144 199694 163946
rect 199862 163144 200522 163946
rect 200690 163144 201350 163946
rect 201518 163144 202270 163946
rect 202438 163144 203098 163946
rect 203266 163144 204018 163946
rect 204186 163144 204846 163946
rect 205014 163144 205766 163946
rect 205934 163144 206594 163946
rect 206762 163144 207422 163946
rect 207590 163144 208342 163946
rect 208510 163144 209170 163946
rect 209338 163144 210090 163946
rect 210258 163144 210918 163946
rect 211086 163144 211838 163946
rect 212006 163144 212666 163946
rect 212834 163144 213494 163946
rect 213662 163144 214414 163946
rect 214582 163144 215242 163946
rect 215410 163144 216162 163946
rect 216330 163144 216990 163946
rect 217158 163144 217818 163946
rect 217986 163144 218738 163946
rect 218906 163144 219566 163946
rect 219734 163144 220486 163946
rect 220654 163144 221314 163946
rect 221482 163144 222234 163946
rect 222402 163144 223062 163946
rect 223230 163144 223890 163946
rect 224058 163144 224810 163946
rect 224978 163144 225638 163946
rect 225806 163144 226558 163946
rect 226726 163144 227386 163946
rect 227554 163144 228306 163946
rect 228474 163144 229134 163946
rect 229302 163144 229962 163946
rect 230130 163144 230882 163946
rect 231050 163144 231710 163946
rect 231878 163144 232630 163946
rect 232798 163144 233458 163946
rect 233626 163144 234286 163946
rect 234454 163144 235206 163946
rect 235374 163144 236034 163946
rect 236202 163144 236954 163946
rect 237122 163144 237782 163946
rect 237950 163144 238702 163946
rect 238870 163144 239530 163946
rect 239698 163144 240358 163946
rect 240526 163144 241278 163946
rect 241446 163144 242106 163946
rect 242274 163144 243026 163946
rect 243194 163144 243854 163946
rect 244022 163144 244774 163946
rect 244942 163144 245602 163946
rect 245770 163144 246430 163946
rect 246598 163144 247350 163946
rect 247518 163144 248178 163946
rect 248346 163144 249098 163946
rect 249266 163144 249926 163946
rect 250094 163144 250846 163946
rect 251014 163144 251674 163946
rect 251842 163144 252502 163946
rect 252670 163144 253422 163946
rect 253590 163144 254250 163946
rect 254418 163144 255170 163946
rect 255338 163144 255998 163946
rect 256166 163144 256826 163946
rect 256994 163144 257746 163946
rect 257914 163144 258574 163946
rect 258742 163144 259494 163946
rect 259662 163144 260322 163946
rect 260490 163144 261242 163946
rect 261410 163144 262070 163946
rect 262238 163144 262898 163946
rect 263066 163144 263818 163946
rect 263986 163144 264646 163946
rect 264814 163144 265566 163946
rect 265734 163144 266394 163946
rect 266562 163144 267314 163946
rect 267482 163144 268142 163946
rect 268310 163144 268970 163946
rect 269138 163144 269890 163946
rect 270058 163144 270718 163946
rect 270886 163144 271638 163946
rect 271806 163144 272466 163946
rect 272634 163144 273294 163946
rect 273462 163144 274214 163946
rect 274382 163144 275042 163946
rect 275210 163144 275962 163946
rect 276130 163144 276790 163946
rect 276958 163144 277710 163946
rect 277878 163144 278538 163946
rect 278706 163144 279366 163946
rect 279534 163144 280286 163946
rect 280454 163144 281114 163946
rect 281282 163144 282034 163946
rect 282202 163144 282862 163946
rect 283030 163144 283782 163946
rect 283950 163144 284610 163946
rect 284778 163144 285438 163946
rect 285606 163144 286358 163946
rect 286526 163144 287186 163946
rect 287354 163144 288106 163946
rect 288274 163144 288934 163946
rect 289102 163144 289762 163946
rect 289930 163144 290682 163946
rect 290850 163144 291510 163946
rect 291678 163144 292430 163946
rect 292598 163144 293258 163946
rect 293426 163144 294178 163946
rect 294346 163144 295006 163946
rect 295174 163144 295834 163946
rect 296002 163144 296754 163946
rect 296922 163144 297582 163946
rect 297750 163144 298502 163946
rect 298670 163144 299330 163946
rect 299498 163144 300250 163946
rect 300418 163144 301078 163946
rect 301246 163144 301906 163946
rect 302074 163144 302826 163946
rect 302994 163144 303654 163946
rect 303822 163144 304574 163946
rect 304742 163144 305402 163946
rect 305570 163144 306322 163946
rect 306490 163144 307150 163946
rect 307318 163144 307978 163946
rect 308146 163144 308898 163946
rect 309066 163144 309726 163946
rect 309894 163144 310646 163946
rect 310814 163144 311474 163946
rect 311642 163144 312302 163946
rect 312470 163144 313222 163946
rect 313390 163144 314050 163946
rect 314218 163144 314970 163946
rect 315138 163144 315798 163946
rect 315966 163144 316718 163946
rect 316886 163144 317546 163946
rect 317714 163144 318374 163946
rect 318542 163144 319294 163946
rect 319462 163144 320122 163946
rect 320290 163144 321042 163946
rect 321210 163144 321870 163946
rect 322038 163144 322790 163946
rect 322958 163144 323618 163946
rect 323786 163144 324446 163946
rect 324614 163144 325366 163946
rect 325534 163144 326194 163946
rect 326362 163144 327114 163946
rect 327282 163144 327942 163946
rect 328110 163144 328770 163946
rect 328938 163144 329690 163946
rect 329858 163144 330518 163946
rect 330686 163144 331438 163946
rect 331606 163144 332266 163946
rect 332434 163144 333186 163946
rect 333354 163144 334014 163946
rect 334182 163144 334842 163946
rect 335010 163144 335762 163946
rect 335930 163144 336590 163946
rect 336758 163144 337510 163946
rect 337678 163144 338338 163946
rect 338506 163144 339258 163946
rect 339426 163144 340086 163946
rect 340254 163144 340914 163946
rect 341082 163144 341834 163946
rect 342002 163144 342662 163946
rect 342830 163144 343582 163946
rect 343750 163144 344410 163946
rect 344578 163144 345330 163946
rect 345498 163144 346158 163946
rect 346326 163144 346986 163946
rect 347154 163144 347906 163946
rect 348074 163144 348734 163946
rect 348902 163144 349654 163946
rect 349822 163144 350482 163946
rect 350650 163144 351310 163946
rect 351478 163144 352230 163946
rect 352398 163144 353058 163946
rect 353226 163144 353978 163946
rect 354146 163144 354806 163946
rect 354974 163144 355726 163946
rect 355894 163144 356554 163946
rect 356722 163144 357382 163946
rect 357550 163144 358302 163946
rect 358470 163144 359130 163946
rect 359298 163144 360050 163946
rect 360218 163144 360878 163946
rect 361046 163144 361798 163946
rect 361966 163144 362626 163946
rect 362794 163144 363454 163946
rect 363622 163144 364374 163946
rect 364542 163144 365202 163946
rect 365370 163144 366122 163946
rect 366290 163144 366950 163946
rect 367118 163144 367778 163946
rect 367946 163144 368698 163946
rect 368866 163144 369526 163946
rect 369694 163144 370446 163946
rect 370614 163144 371274 163946
rect 371442 163144 372194 163946
rect 372362 163144 373022 163946
rect 373190 163144 373850 163946
rect 374018 163144 374770 163946
rect 374938 163144 375598 163946
rect 375766 163144 376518 163946
rect 376686 163144 377346 163946
rect 377514 163144 378266 163946
rect 378434 163144 379094 163946
rect 379262 163144 379922 163946
rect 380090 163144 380842 163946
rect 381010 163144 381670 163946
rect 381838 163144 382590 163946
rect 382758 163144 383418 163946
rect 383586 163144 384338 163946
rect 384506 163144 385166 163946
rect 385334 163144 385994 163946
rect 386162 163144 386914 163946
rect 387082 163144 387742 163946
rect 387910 163144 388662 163946
rect 388830 163144 389490 163946
rect 389658 163144 390318 163946
rect 390486 163144 391238 163946
rect 391406 163144 392066 163946
rect 392234 163144 392986 163946
rect 393154 163144 393814 163946
rect 393982 163144 394734 163946
rect 394902 163144 395562 163946
rect 395730 163144 396390 163946
rect 396558 163144 397310 163946
rect 397478 163144 398138 163946
rect 398306 163144 399058 163946
rect 399226 163144 399886 163946
rect 400054 163144 400806 163946
rect 400974 163144 401634 163946
rect 401802 163144 402462 163946
rect 402630 163144 403382 163946
rect 403550 163144 404210 163946
rect 404378 163144 405130 163946
rect 405298 163144 405958 163946
rect 406126 163144 406786 163946
rect 406954 163144 407706 163946
rect 407874 163144 408534 163946
rect 408702 163144 409454 163946
rect 409622 163144 410282 163946
rect 410450 163144 411202 163946
rect 411370 163144 412030 163946
rect 412198 163144 412858 163946
rect 413026 163144 413778 163946
rect 413946 163144 414606 163946
rect 414774 163144 415526 163946
rect 415694 163144 416354 163946
rect 416522 163144 417274 163946
rect 417442 163144 418102 163946
rect 418270 163144 418930 163946
rect 419098 163144 419850 163946
rect 420018 163144 420678 163946
rect 420846 163144 421598 163946
rect 421766 163144 422426 163946
rect 422594 163144 423346 163946
rect 423514 163144 424174 163946
rect 424342 163144 425002 163946
rect 425170 163144 425922 163946
rect 426090 163144 426750 163946
rect 426918 163144 427670 163946
rect 427838 163144 428498 163946
rect 428666 163144 429326 163946
rect 429494 163144 430246 163946
rect 430414 163144 431074 163946
rect 431242 163144 431994 163946
rect 432162 163144 432822 163946
rect 432990 163144 433742 163946
rect 433910 163144 434570 163946
rect 434738 163144 435398 163946
rect 435566 163144 436318 163946
rect 436486 163144 437146 163946
rect 437314 163144 438066 163946
rect 438234 163144 438894 163946
rect 439062 163144 439814 163946
rect 439982 163144 440642 163946
rect 440810 163144 441470 163946
rect 441638 163144 442390 163946
rect 442558 163144 443218 163946
rect 443386 163144 444138 163946
rect 444306 163144 444966 163946
rect 445134 163144 445794 163946
rect 445962 163144 446714 163946
rect 446882 163144 447542 163946
rect 447710 163144 448462 163946
rect 448630 163144 449290 163946
rect 449458 163144 450210 163946
rect 450378 163144 451038 163946
rect 451206 163144 451866 163946
rect 452034 163144 452786 163946
rect 452954 163144 453614 163946
rect 453782 163144 454534 163946
rect 454702 163144 455362 163946
rect 455530 163144 456282 163946
rect 456450 163144 457110 163946
rect 457278 163144 457938 163946
rect 458106 163144 458858 163946
rect 459026 163144 459686 163946
rect 459854 163144 460606 163946
rect 460774 163144 461434 163946
rect 461602 163144 462354 163946
rect 462522 163144 463182 163946
rect 463350 163144 464010 163946
rect 464178 163144 464930 163946
rect 465098 163144 465758 163946
rect 465926 163144 466678 163946
rect 466846 163144 467506 163946
rect 467674 163144 468334 163946
rect 468502 163144 469254 163946
rect 469422 163144 470082 163946
rect 470250 163144 471002 163946
rect 471170 163144 471830 163946
rect 471998 163144 472750 163946
rect 472918 163144 473578 163946
rect 473746 163144 474406 163946
rect 474574 163144 475326 163946
rect 475494 163144 476154 163946
rect 476322 163144 477074 163946
rect 477242 163144 477902 163946
rect 478070 163144 478822 163946
rect 478990 163144 479650 163946
rect 479818 163144 480478 163946
rect 480646 163144 481398 163946
rect 481566 163144 482226 163946
rect 482394 163144 483146 163946
rect 483314 163144 483974 163946
rect 484142 163144 484802 163946
rect 484970 163144 485722 163946
rect 485890 163144 486550 163946
rect 486718 163144 487470 163946
rect 487638 163144 488298 163946
rect 488466 163144 489218 163946
rect 489386 163144 490046 163946
rect 490214 163144 490874 163946
rect 491042 163144 491794 163946
rect 491962 163144 492622 163946
rect 492790 163144 493542 163946
rect 493710 163144 494370 163946
rect 494538 163144 495290 163946
rect 495458 163144 496118 163946
rect 496286 163144 496946 163946
rect 497114 163144 497866 163946
rect 498034 163144 498694 163946
rect 498862 163144 499614 163946
rect 499782 163144 500442 163946
rect 500610 163144 501362 163946
rect 501530 163144 502190 163946
rect 502358 163144 503018 163946
rect 503186 163144 503938 163946
rect 504106 163144 504766 163946
rect 504934 163144 505686 163946
rect 505854 163144 506514 163946
rect 506682 163144 507342 163946
rect 507510 163144 508262 163946
rect 508430 163144 509090 163946
rect 509258 163144 510010 163946
rect 510178 163144 510838 163946
rect 511006 163144 511758 163946
rect 511926 163144 512586 163946
rect 512754 163144 513414 163946
rect 513582 163144 514334 163946
rect 514502 163144 515162 163946
rect 515330 163144 516082 163946
rect 516250 163144 516910 163946
rect 517078 163144 517830 163946
rect 517998 163144 518658 163946
rect 518826 163144 519486 163946
rect 519654 163144 520406 163946
rect 520574 163144 521234 163946
rect 521402 163144 522154 163946
rect 522322 163144 522982 163946
rect 523150 163144 523810 163946
rect 523978 163144 524730 163946
rect 524898 163144 525558 163946
rect 525726 163144 526478 163946
rect 526646 163144 527306 163946
rect 527474 163144 528226 163946
rect 528394 163144 529054 163946
rect 529222 163144 529882 163946
rect 530050 163144 530802 163946
rect 530970 163144 531630 163946
rect 531798 163144 532550 163946
rect 532718 163144 533378 163946
rect 533546 163144 534298 163946
rect 534466 163144 535126 163946
rect 535294 163144 535954 163946
rect 536122 163144 536874 163946
rect 537042 163144 537702 163946
rect 537870 163144 538622 163946
rect 538790 163144 539450 163946
rect 388 856 539560 163144
rect 388 711 33634 856
rect 33802 711 101070 856
rect 101238 711 168598 856
rect 168766 711 236126 856
rect 236294 711 303654 856
rect 303822 711 371090 856
rect 371258 711 438618 856
rect 438786 711 506146 856
rect 506314 711 539560 856
<< metal3 >>
rect 539200 163072 540000 163192
rect 539200 161576 540000 161696
rect 539200 160080 540000 160200
rect 539200 158584 540000 158704
rect 539200 157088 540000 157208
rect 539200 155592 540000 155712
rect 539200 153960 540000 154080
rect 539200 152464 540000 152584
rect 539200 150968 540000 151088
rect 539200 149472 540000 149592
rect 539200 147976 540000 148096
rect 539200 146480 540000 146600
rect 539200 144848 540000 144968
rect 539200 143352 540000 143472
rect 539200 141856 540000 141976
rect 539200 140360 540000 140480
rect 539200 138864 540000 138984
rect 539200 137368 540000 137488
rect 539200 135736 540000 135856
rect 539200 134240 540000 134360
rect 539200 132744 540000 132864
rect 539200 131248 540000 131368
rect 539200 129752 540000 129872
rect 539200 128256 540000 128376
rect 539200 126624 540000 126744
rect 539200 125128 540000 125248
rect 539200 123632 540000 123752
rect 539200 122136 540000 122256
rect 539200 120640 540000 120760
rect 539200 119144 540000 119264
rect 539200 117512 540000 117632
rect 539200 116016 540000 116136
rect 539200 114520 540000 114640
rect 539200 113024 540000 113144
rect 539200 111528 540000 111648
rect 539200 110032 540000 110152
rect 539200 108400 540000 108520
rect 539200 106904 540000 107024
rect 539200 105408 540000 105528
rect 539200 103912 540000 104032
rect 539200 102416 540000 102536
rect 539200 100920 540000 101040
rect 539200 99288 540000 99408
rect 539200 97792 540000 97912
rect 539200 96296 540000 96416
rect 539200 94800 540000 94920
rect 539200 93304 540000 93424
rect 539200 91808 540000 91928
rect 539200 90176 540000 90296
rect 539200 88680 540000 88800
rect 539200 87184 540000 87304
rect 539200 85688 540000 85808
rect 539200 84192 540000 84312
rect 539200 82696 540000 82816
rect 539200 81064 540000 81184
rect 539200 79568 540000 79688
rect 539200 78072 540000 78192
rect 539200 76576 540000 76696
rect 539200 75080 540000 75200
rect 539200 73584 540000 73704
rect 539200 71952 540000 72072
rect 539200 70456 540000 70576
rect 539200 68960 540000 69080
rect 539200 67464 540000 67584
rect 539200 65968 540000 66088
rect 539200 64472 540000 64592
rect 539200 62840 540000 62960
rect 539200 61344 540000 61464
rect 539200 59848 540000 59968
rect 539200 58352 540000 58472
rect 539200 56856 540000 56976
rect 539200 55360 540000 55480
rect 539200 53728 540000 53848
rect 539200 52232 540000 52352
rect 539200 50736 540000 50856
rect 539200 49240 540000 49360
rect 539200 47744 540000 47864
rect 539200 46248 540000 46368
rect 539200 44616 540000 44736
rect 539200 43120 540000 43240
rect 539200 41624 540000 41744
rect 539200 40128 540000 40248
rect 539200 38632 540000 38752
rect 539200 37136 540000 37256
rect 539200 35504 540000 35624
rect 539200 34008 540000 34128
rect 539200 32512 540000 32632
rect 539200 31016 540000 31136
rect 539200 29520 540000 29640
rect 539200 28024 540000 28144
rect 539200 26392 540000 26512
rect 539200 24896 540000 25016
rect 539200 23400 540000 23520
rect 539200 21904 540000 22024
rect 539200 20408 540000 20528
rect 539200 18912 540000 19032
rect 539200 17280 540000 17400
rect 539200 15784 540000 15904
rect 539200 14288 540000 14408
rect 539200 12792 540000 12912
rect 539200 11296 540000 11416
rect 539200 9800 540000 9920
rect 539200 8168 540000 8288
rect 539200 6672 540000 6792
rect 539200 5176 540000 5296
rect 539200 3680 540000 3800
rect 539200 2184 540000 2304
rect 539200 688 540000 808
<< obsm3 >>
rect 5993 162992 539120 163165
rect 5993 161776 539200 162992
rect 5993 161496 539120 161776
rect 5993 160280 539200 161496
rect 5993 160000 539120 160280
rect 5993 158784 539200 160000
rect 5993 158504 539120 158784
rect 5993 157288 539200 158504
rect 5993 157008 539120 157288
rect 5993 155792 539200 157008
rect 5993 155512 539120 155792
rect 5993 154160 539200 155512
rect 5993 153880 539120 154160
rect 5993 152664 539200 153880
rect 5993 152384 539120 152664
rect 5993 151168 539200 152384
rect 5993 150888 539120 151168
rect 5993 149672 539200 150888
rect 5993 149392 539120 149672
rect 5993 148176 539200 149392
rect 5993 147896 539120 148176
rect 5993 146680 539200 147896
rect 5993 146400 539120 146680
rect 5993 145048 539200 146400
rect 5993 144768 539120 145048
rect 5993 143552 539200 144768
rect 5993 143272 539120 143552
rect 5993 142056 539200 143272
rect 5993 141776 539120 142056
rect 5993 140560 539200 141776
rect 5993 140280 539120 140560
rect 5993 139064 539200 140280
rect 5993 138784 539120 139064
rect 5993 137568 539200 138784
rect 5993 137288 539120 137568
rect 5993 135936 539200 137288
rect 5993 135656 539120 135936
rect 5993 134440 539200 135656
rect 5993 134160 539120 134440
rect 5993 132944 539200 134160
rect 5993 132664 539120 132944
rect 5993 131448 539200 132664
rect 5993 131168 539120 131448
rect 5993 129952 539200 131168
rect 5993 129672 539120 129952
rect 5993 128456 539200 129672
rect 5993 128176 539120 128456
rect 5993 126824 539200 128176
rect 5993 126544 539120 126824
rect 5993 125328 539200 126544
rect 5993 125048 539120 125328
rect 5993 123832 539200 125048
rect 5993 123552 539120 123832
rect 5993 122336 539200 123552
rect 5993 122056 539120 122336
rect 5993 120840 539200 122056
rect 5993 120560 539120 120840
rect 5993 119344 539200 120560
rect 5993 119064 539120 119344
rect 5993 117712 539200 119064
rect 5993 117432 539120 117712
rect 5993 116216 539200 117432
rect 5993 115936 539120 116216
rect 5993 114720 539200 115936
rect 5993 114440 539120 114720
rect 5993 113224 539200 114440
rect 5993 112944 539120 113224
rect 5993 111728 539200 112944
rect 5993 111448 539120 111728
rect 5993 110232 539200 111448
rect 5993 109952 539120 110232
rect 5993 108600 539200 109952
rect 5993 108320 539120 108600
rect 5993 107104 539200 108320
rect 5993 106824 539120 107104
rect 5993 105608 539200 106824
rect 5993 105328 539120 105608
rect 5993 104112 539200 105328
rect 5993 103832 539120 104112
rect 5993 102616 539200 103832
rect 5993 102336 539120 102616
rect 5993 101120 539200 102336
rect 5993 100840 539120 101120
rect 5993 99488 539200 100840
rect 5993 99208 539120 99488
rect 5993 97992 539200 99208
rect 5993 97712 539120 97992
rect 5993 96496 539200 97712
rect 5993 96216 539120 96496
rect 5993 95000 539200 96216
rect 5993 94720 539120 95000
rect 5993 93504 539200 94720
rect 5993 93224 539120 93504
rect 5993 92008 539200 93224
rect 5993 91728 539120 92008
rect 5993 90376 539200 91728
rect 5993 90096 539120 90376
rect 5993 88880 539200 90096
rect 5993 88600 539120 88880
rect 5993 87384 539200 88600
rect 5993 87104 539120 87384
rect 5993 85888 539200 87104
rect 5993 85608 539120 85888
rect 5993 84392 539200 85608
rect 5993 84112 539120 84392
rect 5993 82896 539200 84112
rect 5993 82616 539120 82896
rect 5993 81264 539200 82616
rect 5993 80984 539120 81264
rect 5993 79768 539200 80984
rect 5993 79488 539120 79768
rect 5993 78272 539200 79488
rect 5993 77992 539120 78272
rect 5993 76776 539200 77992
rect 5993 76496 539120 76776
rect 5993 75280 539200 76496
rect 5993 75000 539120 75280
rect 5993 73784 539200 75000
rect 5993 73504 539120 73784
rect 5993 72152 539200 73504
rect 5993 71872 539120 72152
rect 5993 70656 539200 71872
rect 5993 70376 539120 70656
rect 5993 69160 539200 70376
rect 5993 68880 539120 69160
rect 5993 67664 539200 68880
rect 5993 67384 539120 67664
rect 5993 66168 539200 67384
rect 5993 65888 539120 66168
rect 5993 64672 539200 65888
rect 5993 64392 539120 64672
rect 5993 63040 539200 64392
rect 5993 62760 539120 63040
rect 5993 61544 539200 62760
rect 5993 61264 539120 61544
rect 5993 60048 539200 61264
rect 5993 59768 539120 60048
rect 5993 58552 539200 59768
rect 5993 58272 539120 58552
rect 5993 57056 539200 58272
rect 5993 56776 539120 57056
rect 5993 55560 539200 56776
rect 5993 55280 539120 55560
rect 5993 53928 539200 55280
rect 5993 53648 539120 53928
rect 5993 52432 539200 53648
rect 5993 52152 539120 52432
rect 5993 50936 539200 52152
rect 5993 50656 539120 50936
rect 5993 49440 539200 50656
rect 5993 49160 539120 49440
rect 5993 47944 539200 49160
rect 5993 47664 539120 47944
rect 5993 46448 539200 47664
rect 5993 46168 539120 46448
rect 5993 44816 539200 46168
rect 5993 44536 539120 44816
rect 5993 43320 539200 44536
rect 5993 43040 539120 43320
rect 5993 41824 539200 43040
rect 5993 41544 539120 41824
rect 5993 40328 539200 41544
rect 5993 40048 539120 40328
rect 5993 38832 539200 40048
rect 5993 38552 539120 38832
rect 5993 37336 539200 38552
rect 5993 37056 539120 37336
rect 5993 35704 539200 37056
rect 5993 35424 539120 35704
rect 5993 34208 539200 35424
rect 5993 33928 539120 34208
rect 5993 32712 539200 33928
rect 5993 32432 539120 32712
rect 5993 31216 539200 32432
rect 5993 30936 539120 31216
rect 5993 29720 539200 30936
rect 5993 29440 539120 29720
rect 5993 28224 539200 29440
rect 5993 27944 539120 28224
rect 5993 26592 539200 27944
rect 5993 26312 539120 26592
rect 5993 25096 539200 26312
rect 5993 24816 539120 25096
rect 5993 23600 539200 24816
rect 5993 23320 539120 23600
rect 5993 22104 539200 23320
rect 5993 21824 539120 22104
rect 5993 20608 539200 21824
rect 5993 20328 539120 20608
rect 5993 19112 539200 20328
rect 5993 18832 539120 19112
rect 5993 17480 539200 18832
rect 5993 17200 539120 17480
rect 5993 15984 539200 17200
rect 5993 15704 539120 15984
rect 5993 14488 539200 15704
rect 5993 14208 539120 14488
rect 5993 12992 539200 14208
rect 5993 12712 539120 12992
rect 5993 11496 539200 12712
rect 5993 11216 539120 11496
rect 5993 10000 539200 11216
rect 5993 9720 539120 10000
rect 5993 8368 539200 9720
rect 5993 8088 539120 8368
rect 5993 6872 539200 8088
rect 5993 6592 539120 6872
rect 5993 5376 539200 6592
rect 5993 5096 539120 5376
rect 5993 3880 539200 5096
rect 5993 3600 539120 3880
rect 5993 2384 539200 3600
rect 5993 2104 539120 2384
rect 5993 888 539200 2104
rect 5993 715 539120 888
<< obsm4 >>
rect 4004 4156 528018 158898
<< metal5 >>
rect 1104 148346 2000 148666
rect 116000 148346 128000 148666
rect 532000 148346 538844 148666
rect 1104 135346 2000 135666
rect 116000 135346 128000 135666
rect 532000 135346 538844 135666
rect 1104 122346 2000 122666
rect 116000 122346 128000 122666
rect 532000 122346 538844 122666
rect 1104 109346 2000 109666
rect 116000 109346 128000 109666
rect 532000 109346 538844 109666
rect 1104 96346 2000 96666
rect 116000 96346 128000 96666
rect 532000 96346 538844 96666
rect 1104 83346 2000 83666
rect 116000 83346 128000 83666
rect 532000 83346 538844 83666
rect 1104 70346 2000 70666
rect 116000 70346 128000 70666
rect 532000 70346 538844 70666
rect 1104 57346 2000 57666
rect 116000 57346 128000 57666
rect 532000 57346 538844 57666
rect 1104 44346 2000 44666
rect 116000 44346 128000 44666
rect 532000 44346 538844 44666
rect 1104 31346 2000 31666
rect 116000 31346 128000 31666
rect 532000 31346 538844 31666
rect 1104 18346 2000 18666
rect 116000 18346 128000 18666
rect 532000 18346 538844 18666
rect 1104 5346 2000 5666
rect 116000 5346 128000 5666
rect 532000 5346 538844 5666
<< obsm5 >>
rect 4004 148986 528820 158940
rect 4004 148026 115680 148986
rect 128320 148026 528820 148986
rect 4004 135986 528820 148026
rect 4004 135026 115680 135986
rect 128320 135026 528820 135986
rect 4004 122986 528820 135026
rect 4004 122026 115680 122986
rect 128320 122026 528820 122986
rect 4004 109986 528820 122026
rect 4004 109026 115680 109986
rect 128320 109026 528820 109986
rect 4004 96986 528820 109026
rect 4004 96026 115680 96986
rect 128320 96026 528820 96986
rect 4004 83986 528820 96026
rect 4004 83026 115680 83986
rect 128320 83026 528820 83986
rect 4004 70986 528820 83026
rect 4004 70026 115680 70986
rect 128320 70026 528820 70986
rect 4004 57986 528820 70026
rect 4004 57026 115680 57986
rect 128320 57026 528820 57986
rect 4004 44986 528820 57026
rect 4004 44026 115680 44986
rect 128320 44026 528820 44986
rect 4004 31986 528820 44026
rect 4004 31026 115680 31986
rect 128320 31026 528820 31986
rect 4004 18986 528820 31026
rect 4004 18026 115680 18986
rect 128320 18026 528820 18986
rect 4004 5986 528820 18026
rect 4004 5026 115680 5986
rect 128320 5026 528820 5986
rect 4004 4156 528820 5026
<< labels >>
rlabel metal5 s 1104 18346 2000 18666 6 VGND
port 1 nsew ground input
rlabel metal5 s 116000 18346 128000 18666 6 VGND
port 1 nsew ground input
rlabel metal5 s 532000 18346 538844 18666 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 44346 2000 44666 6 VGND
port 1 nsew ground input
rlabel metal5 s 116000 44346 128000 44666 6 VGND
port 1 nsew ground input
rlabel metal5 s 532000 44346 538844 44666 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 70346 2000 70666 6 VGND
port 1 nsew ground input
rlabel metal5 s 116000 70346 128000 70666 6 VGND
port 1 nsew ground input
rlabel metal5 s 532000 70346 538844 70666 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 96346 2000 96666 6 VGND
port 1 nsew ground input
rlabel metal5 s 116000 96346 128000 96666 6 VGND
port 1 nsew ground input
rlabel metal5 s 532000 96346 538844 96666 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 122346 2000 122666 6 VGND
port 1 nsew ground input
rlabel metal5 s 116000 122346 128000 122666 6 VGND
port 1 nsew ground input
rlabel metal5 s 532000 122346 538844 122666 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 148346 2000 148666 6 VGND
port 1 nsew ground input
rlabel metal5 s 116000 148346 128000 148666 6 VGND
port 1 nsew ground input
rlabel metal5 s 532000 148346 538844 148666 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 5346 2000 5666 6 VPWR
port 2 nsew power input
rlabel metal5 s 116000 5346 128000 5666 6 VPWR
port 2 nsew power input
rlabel metal5 s 532000 5346 538844 5666 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 31346 2000 31666 6 VPWR
port 2 nsew power input
rlabel metal5 s 116000 31346 128000 31666 6 VPWR
port 2 nsew power input
rlabel metal5 s 532000 31346 538844 31666 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 57346 2000 57666 6 VPWR
port 2 nsew power input
rlabel metal5 s 116000 57346 128000 57666 6 VPWR
port 2 nsew power input
rlabel metal5 s 532000 57346 538844 57666 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 83346 2000 83666 6 VPWR
port 2 nsew power input
rlabel metal5 s 116000 83346 128000 83666 6 VPWR
port 2 nsew power input
rlabel metal5 s 532000 83346 538844 83666 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 109346 2000 109666 6 VPWR
port 2 nsew power input
rlabel metal5 s 116000 109346 128000 109666 6 VPWR
port 2 nsew power input
rlabel metal5 s 532000 109346 538844 109666 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 135346 2000 135666 6 VPWR
port 2 nsew power input
rlabel metal5 s 116000 135346 128000 135666 6 VPWR
port 2 nsew power input
rlabel metal5 s 532000 135346 538844 135666 6 VPWR
port 2 nsew power input
rlabel metal2 s 506202 0 506258 800 6 core_clk
port 3 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 core_rstn
port 4 nsew signal input
rlabel metal3 s 539200 64472 540000 64592 6 debug_in
port 5 nsew signal input
rlabel metal3 s 539200 65968 540000 66088 6 debug_mode
port 6 nsew signal output
rlabel metal3 s 539200 67464 540000 67584 6 debug_oeb
port 7 nsew signal output
rlabel metal3 s 539200 68960 540000 69080 6 debug_out
port 8 nsew signal output
rlabel metal3 s 539200 144848 540000 144968 6 flash_clk
port 9 nsew signal output
rlabel metal3 s 539200 143352 540000 143472 6 flash_csb
port 10 nsew signal output
rlabel metal3 s 539200 146480 540000 146600 6 flash_io0_di
port 11 nsew signal input
rlabel metal3 s 539200 147976 540000 148096 6 flash_io0_do
port 12 nsew signal output
rlabel metal3 s 539200 149472 540000 149592 6 flash_io0_oeb
port 13 nsew signal output
rlabel metal3 s 539200 150968 540000 151088 6 flash_io1_di
port 14 nsew signal input
rlabel metal3 s 539200 152464 540000 152584 6 flash_io1_do
port 15 nsew signal output
rlabel metal3 s 539200 153960 540000 154080 6 flash_io1_oeb
port 16 nsew signal output
rlabel metal3 s 539200 155592 540000 155712 6 flash_io2_di
port 17 nsew signal input
rlabel metal3 s 539200 157088 540000 157208 6 flash_io2_do
port 18 nsew signal output
rlabel metal3 s 539200 158584 540000 158704 6 flash_io2_oeb
port 19 nsew signal output
rlabel metal3 s 539200 160080 540000 160200 6 flash_io3_di
port 20 nsew signal input
rlabel metal3 s 539200 161576 540000 161696 6 flash_io3_do
port 21 nsew signal output
rlabel metal3 s 539200 163072 540000 163192 6 flash_io3_oeb
port 22 nsew signal output
rlabel metal2 s 101126 0 101182 800 6 gpio_in_pad
port 23 nsew signal input
rlabel metal2 s 168654 0 168710 800 6 gpio_inenb_pad
port 24 nsew signal output
rlabel metal2 s 236182 0 236238 800 6 gpio_mode0_pad
port 25 nsew signal output
rlabel metal2 s 303710 0 303766 800 6 gpio_mode1_pad
port 26 nsew signal output
rlabel metal2 s 371146 0 371202 800 6 gpio_out_pad
port 27 nsew signal output
rlabel metal2 s 438674 0 438730 800 6 gpio_outenb_pad
port 28 nsew signal output
rlabel metal3 s 539200 91808 540000 91928 6 hk_ack_i
port 29 nsew signal input
rlabel metal3 s 539200 94800 540000 94920 6 hk_dat_i[0]
port 30 nsew signal input
rlabel metal3 s 539200 110032 540000 110152 6 hk_dat_i[10]
port 31 nsew signal input
rlabel metal3 s 539200 111528 540000 111648 6 hk_dat_i[11]
port 32 nsew signal input
rlabel metal3 s 539200 113024 540000 113144 6 hk_dat_i[12]
port 33 nsew signal input
rlabel metal3 s 539200 114520 540000 114640 6 hk_dat_i[13]
port 34 nsew signal input
rlabel metal3 s 539200 116016 540000 116136 6 hk_dat_i[14]
port 35 nsew signal input
rlabel metal3 s 539200 117512 540000 117632 6 hk_dat_i[15]
port 36 nsew signal input
rlabel metal3 s 539200 119144 540000 119264 6 hk_dat_i[16]
port 37 nsew signal input
rlabel metal3 s 539200 120640 540000 120760 6 hk_dat_i[17]
port 38 nsew signal input
rlabel metal3 s 539200 122136 540000 122256 6 hk_dat_i[18]
port 39 nsew signal input
rlabel metal3 s 539200 123632 540000 123752 6 hk_dat_i[19]
port 40 nsew signal input
rlabel metal3 s 539200 96296 540000 96416 6 hk_dat_i[1]
port 41 nsew signal input
rlabel metal3 s 539200 125128 540000 125248 6 hk_dat_i[20]
port 42 nsew signal input
rlabel metal3 s 539200 126624 540000 126744 6 hk_dat_i[21]
port 43 nsew signal input
rlabel metal3 s 539200 128256 540000 128376 6 hk_dat_i[22]
port 44 nsew signal input
rlabel metal3 s 539200 129752 540000 129872 6 hk_dat_i[23]
port 45 nsew signal input
rlabel metal3 s 539200 131248 540000 131368 6 hk_dat_i[24]
port 46 nsew signal input
rlabel metal3 s 539200 132744 540000 132864 6 hk_dat_i[25]
port 47 nsew signal input
rlabel metal3 s 539200 134240 540000 134360 6 hk_dat_i[26]
port 48 nsew signal input
rlabel metal3 s 539200 135736 540000 135856 6 hk_dat_i[27]
port 49 nsew signal input
rlabel metal3 s 539200 137368 540000 137488 6 hk_dat_i[28]
port 50 nsew signal input
rlabel metal3 s 539200 138864 540000 138984 6 hk_dat_i[29]
port 51 nsew signal input
rlabel metal3 s 539200 97792 540000 97912 6 hk_dat_i[2]
port 52 nsew signal input
rlabel metal3 s 539200 140360 540000 140480 6 hk_dat_i[30]
port 53 nsew signal input
rlabel metal3 s 539200 141856 540000 141976 6 hk_dat_i[31]
port 54 nsew signal input
rlabel metal3 s 539200 99288 540000 99408 6 hk_dat_i[3]
port 55 nsew signal input
rlabel metal3 s 539200 100920 540000 101040 6 hk_dat_i[4]
port 56 nsew signal input
rlabel metal3 s 539200 102416 540000 102536 6 hk_dat_i[5]
port 57 nsew signal input
rlabel metal3 s 539200 103912 540000 104032 6 hk_dat_i[6]
port 58 nsew signal input
rlabel metal3 s 539200 105408 540000 105528 6 hk_dat_i[7]
port 59 nsew signal input
rlabel metal3 s 539200 106904 540000 107024 6 hk_dat_i[8]
port 60 nsew signal input
rlabel metal3 s 539200 108400 540000 108520 6 hk_dat_i[9]
port 61 nsew signal input
rlabel metal3 s 539200 93304 540000 93424 6 hk_stb_o
port 62 nsew signal output
rlabel metal2 s 537758 163200 537814 164000 6 irq[0]
port 63 nsew signal input
rlabel metal2 s 538678 163200 538734 164000 6 irq[1]
port 64 nsew signal input
rlabel metal2 s 539506 163200 539562 164000 6 irq[2]
port 65 nsew signal input
rlabel metal3 s 539200 75080 540000 75200 6 irq[3]
port 66 nsew signal input
rlabel metal3 s 539200 73584 540000 73704 6 irq[4]
port 67 nsew signal input
rlabel metal3 s 539200 71952 540000 72072 6 irq[5]
port 68 nsew signal input
rlabel metal2 s 386 163200 442 164000 6 la_iena[0]
port 69 nsew signal output
rlabel metal2 s 347042 163200 347098 164000 6 la_iena[100]
port 70 nsew signal output
rlabel metal2 s 350538 163200 350594 164000 6 la_iena[101]
port 71 nsew signal output
rlabel metal2 s 354034 163200 354090 164000 6 la_iena[102]
port 72 nsew signal output
rlabel metal2 s 357438 163200 357494 164000 6 la_iena[103]
port 73 nsew signal output
rlabel metal2 s 360934 163200 360990 164000 6 la_iena[104]
port 74 nsew signal output
rlabel metal2 s 364430 163200 364486 164000 6 la_iena[105]
port 75 nsew signal output
rlabel metal2 s 367834 163200 367890 164000 6 la_iena[106]
port 76 nsew signal output
rlabel metal2 s 371330 163200 371386 164000 6 la_iena[107]
port 77 nsew signal output
rlabel metal2 s 374826 163200 374882 164000 6 la_iena[108]
port 78 nsew signal output
rlabel metal2 s 378322 163200 378378 164000 6 la_iena[109]
port 79 nsew signal output
rlabel metal2 s 34978 163200 35034 164000 6 la_iena[10]
port 80 nsew signal output
rlabel metal2 s 381726 163200 381782 164000 6 la_iena[110]
port 81 nsew signal output
rlabel metal2 s 385222 163200 385278 164000 6 la_iena[111]
port 82 nsew signal output
rlabel metal2 s 388718 163200 388774 164000 6 la_iena[112]
port 83 nsew signal output
rlabel metal2 s 392122 163200 392178 164000 6 la_iena[113]
port 84 nsew signal output
rlabel metal2 s 395618 163200 395674 164000 6 la_iena[114]
port 85 nsew signal output
rlabel metal2 s 399114 163200 399170 164000 6 la_iena[115]
port 86 nsew signal output
rlabel metal2 s 402518 163200 402574 164000 6 la_iena[116]
port 87 nsew signal output
rlabel metal2 s 406014 163200 406070 164000 6 la_iena[117]
port 88 nsew signal output
rlabel metal2 s 409510 163200 409566 164000 6 la_iena[118]
port 89 nsew signal output
rlabel metal2 s 412914 163200 412970 164000 6 la_iena[119]
port 90 nsew signal output
rlabel metal2 s 38474 163200 38530 164000 6 la_iena[11]
port 91 nsew signal output
rlabel metal2 s 416410 163200 416466 164000 6 la_iena[120]
port 92 nsew signal output
rlabel metal2 s 419906 163200 419962 164000 6 la_iena[121]
port 93 nsew signal output
rlabel metal2 s 423402 163200 423458 164000 6 la_iena[122]
port 94 nsew signal output
rlabel metal2 s 426806 163200 426862 164000 6 la_iena[123]
port 95 nsew signal output
rlabel metal2 s 430302 163200 430358 164000 6 la_iena[124]
port 96 nsew signal output
rlabel metal2 s 433798 163200 433854 164000 6 la_iena[125]
port 97 nsew signal output
rlabel metal2 s 437202 163200 437258 164000 6 la_iena[126]
port 98 nsew signal output
rlabel metal2 s 440698 163200 440754 164000 6 la_iena[127]
port 99 nsew signal output
rlabel metal2 s 41970 163200 42026 164000 6 la_iena[12]
port 100 nsew signal output
rlabel metal2 s 45374 163200 45430 164000 6 la_iena[13]
port 101 nsew signal output
rlabel metal2 s 48870 163200 48926 164000 6 la_iena[14]
port 102 nsew signal output
rlabel metal2 s 52366 163200 52422 164000 6 la_iena[15]
port 103 nsew signal output
rlabel metal2 s 55862 163200 55918 164000 6 la_iena[16]
port 104 nsew signal output
rlabel metal2 s 59266 163200 59322 164000 6 la_iena[17]
port 105 nsew signal output
rlabel metal2 s 62762 163200 62818 164000 6 la_iena[18]
port 106 nsew signal output
rlabel metal2 s 66258 163200 66314 164000 6 la_iena[19]
port 107 nsew signal output
rlabel metal2 s 3790 163200 3846 164000 6 la_iena[1]
port 108 nsew signal output
rlabel metal2 s 69662 163200 69718 164000 6 la_iena[20]
port 109 nsew signal output
rlabel metal2 s 73158 163200 73214 164000 6 la_iena[21]
port 110 nsew signal output
rlabel metal2 s 76654 163200 76710 164000 6 la_iena[22]
port 111 nsew signal output
rlabel metal2 s 80058 163200 80114 164000 6 la_iena[23]
port 112 nsew signal output
rlabel metal2 s 83554 163200 83610 164000 6 la_iena[24]
port 113 nsew signal output
rlabel metal2 s 87050 163200 87106 164000 6 la_iena[25]
port 114 nsew signal output
rlabel metal2 s 90454 163200 90510 164000 6 la_iena[26]
port 115 nsew signal output
rlabel metal2 s 93950 163200 94006 164000 6 la_iena[27]
port 116 nsew signal output
rlabel metal2 s 97446 163200 97502 164000 6 la_iena[28]
port 117 nsew signal output
rlabel metal2 s 100850 163200 100906 164000 6 la_iena[29]
port 118 nsew signal output
rlabel metal2 s 7286 163200 7342 164000 6 la_iena[2]
port 119 nsew signal output
rlabel metal2 s 104346 163200 104402 164000 6 la_iena[30]
port 120 nsew signal output
rlabel metal2 s 107842 163200 107898 164000 6 la_iena[31]
port 121 nsew signal output
rlabel metal2 s 111338 163200 111394 164000 6 la_iena[32]
port 122 nsew signal output
rlabel metal2 s 114742 163200 114798 164000 6 la_iena[33]
port 123 nsew signal output
rlabel metal2 s 118238 163200 118294 164000 6 la_iena[34]
port 124 nsew signal output
rlabel metal2 s 121734 163200 121790 164000 6 la_iena[35]
port 125 nsew signal output
rlabel metal2 s 125138 163200 125194 164000 6 la_iena[36]
port 126 nsew signal output
rlabel metal2 s 128634 163200 128690 164000 6 la_iena[37]
port 127 nsew signal output
rlabel metal2 s 132130 163200 132186 164000 6 la_iena[38]
port 128 nsew signal output
rlabel metal2 s 135534 163200 135590 164000 6 la_iena[39]
port 129 nsew signal output
rlabel metal2 s 10782 163200 10838 164000 6 la_iena[3]
port 130 nsew signal output
rlabel metal2 s 139030 163200 139086 164000 6 la_iena[40]
port 131 nsew signal output
rlabel metal2 s 142526 163200 142582 164000 6 la_iena[41]
port 132 nsew signal output
rlabel metal2 s 145930 163200 145986 164000 6 la_iena[42]
port 133 nsew signal output
rlabel metal2 s 149426 163200 149482 164000 6 la_iena[43]
port 134 nsew signal output
rlabel metal2 s 152922 163200 152978 164000 6 la_iena[44]
port 135 nsew signal output
rlabel metal2 s 156326 163200 156382 164000 6 la_iena[45]
port 136 nsew signal output
rlabel metal2 s 159822 163200 159878 164000 6 la_iena[46]
port 137 nsew signal output
rlabel metal2 s 163318 163200 163374 164000 6 la_iena[47]
port 138 nsew signal output
rlabel metal2 s 166814 163200 166870 164000 6 la_iena[48]
port 139 nsew signal output
rlabel metal2 s 170218 163200 170274 164000 6 la_iena[49]
port 140 nsew signal output
rlabel metal2 s 14186 163200 14242 164000 6 la_iena[4]
port 141 nsew signal output
rlabel metal2 s 173714 163200 173770 164000 6 la_iena[50]
port 142 nsew signal output
rlabel metal2 s 177210 163200 177266 164000 6 la_iena[51]
port 143 nsew signal output
rlabel metal2 s 180614 163200 180670 164000 6 la_iena[52]
port 144 nsew signal output
rlabel metal2 s 184110 163200 184166 164000 6 la_iena[53]
port 145 nsew signal output
rlabel metal2 s 187606 163200 187662 164000 6 la_iena[54]
port 146 nsew signal output
rlabel metal2 s 191010 163200 191066 164000 6 la_iena[55]
port 147 nsew signal output
rlabel metal2 s 194506 163200 194562 164000 6 la_iena[56]
port 148 nsew signal output
rlabel metal2 s 198002 163200 198058 164000 6 la_iena[57]
port 149 nsew signal output
rlabel metal2 s 201406 163200 201462 164000 6 la_iena[58]
port 150 nsew signal output
rlabel metal2 s 204902 163200 204958 164000 6 la_iena[59]
port 151 nsew signal output
rlabel metal2 s 17682 163200 17738 164000 6 la_iena[5]
port 152 nsew signal output
rlabel metal2 s 208398 163200 208454 164000 6 la_iena[60]
port 153 nsew signal output
rlabel metal2 s 211894 163200 211950 164000 6 la_iena[61]
port 154 nsew signal output
rlabel metal2 s 215298 163200 215354 164000 6 la_iena[62]
port 155 nsew signal output
rlabel metal2 s 218794 163200 218850 164000 6 la_iena[63]
port 156 nsew signal output
rlabel metal2 s 222290 163200 222346 164000 6 la_iena[64]
port 157 nsew signal output
rlabel metal2 s 225694 163200 225750 164000 6 la_iena[65]
port 158 nsew signal output
rlabel metal2 s 229190 163200 229246 164000 6 la_iena[66]
port 159 nsew signal output
rlabel metal2 s 232686 163200 232742 164000 6 la_iena[67]
port 160 nsew signal output
rlabel metal2 s 236090 163200 236146 164000 6 la_iena[68]
port 161 nsew signal output
rlabel metal2 s 239586 163200 239642 164000 6 la_iena[69]
port 162 nsew signal output
rlabel metal2 s 21178 163200 21234 164000 6 la_iena[6]
port 163 nsew signal output
rlabel metal2 s 243082 163200 243138 164000 6 la_iena[70]
port 164 nsew signal output
rlabel metal2 s 246486 163200 246542 164000 6 la_iena[71]
port 165 nsew signal output
rlabel metal2 s 249982 163200 250038 164000 6 la_iena[72]
port 166 nsew signal output
rlabel metal2 s 253478 163200 253534 164000 6 la_iena[73]
port 167 nsew signal output
rlabel metal2 s 256882 163200 256938 164000 6 la_iena[74]
port 168 nsew signal output
rlabel metal2 s 260378 163200 260434 164000 6 la_iena[75]
port 169 nsew signal output
rlabel metal2 s 263874 163200 263930 164000 6 la_iena[76]
port 170 nsew signal output
rlabel metal2 s 267370 163200 267426 164000 6 la_iena[77]
port 171 nsew signal output
rlabel metal2 s 270774 163200 270830 164000 6 la_iena[78]
port 172 nsew signal output
rlabel metal2 s 274270 163200 274326 164000 6 la_iena[79]
port 173 nsew signal output
rlabel metal2 s 24582 163200 24638 164000 6 la_iena[7]
port 174 nsew signal output
rlabel metal2 s 277766 163200 277822 164000 6 la_iena[80]
port 175 nsew signal output
rlabel metal2 s 281170 163200 281226 164000 6 la_iena[81]
port 176 nsew signal output
rlabel metal2 s 284666 163200 284722 164000 6 la_iena[82]
port 177 nsew signal output
rlabel metal2 s 288162 163200 288218 164000 6 la_iena[83]
port 178 nsew signal output
rlabel metal2 s 291566 163200 291622 164000 6 la_iena[84]
port 179 nsew signal output
rlabel metal2 s 295062 163200 295118 164000 6 la_iena[85]
port 180 nsew signal output
rlabel metal2 s 298558 163200 298614 164000 6 la_iena[86]
port 181 nsew signal output
rlabel metal2 s 301962 163200 302018 164000 6 la_iena[87]
port 182 nsew signal output
rlabel metal2 s 305458 163200 305514 164000 6 la_iena[88]
port 183 nsew signal output
rlabel metal2 s 308954 163200 309010 164000 6 la_iena[89]
port 184 nsew signal output
rlabel metal2 s 28078 163200 28134 164000 6 la_iena[8]
port 185 nsew signal output
rlabel metal2 s 312358 163200 312414 164000 6 la_iena[90]
port 186 nsew signal output
rlabel metal2 s 315854 163200 315910 164000 6 la_iena[91]
port 187 nsew signal output
rlabel metal2 s 319350 163200 319406 164000 6 la_iena[92]
port 188 nsew signal output
rlabel metal2 s 322846 163200 322902 164000 6 la_iena[93]
port 189 nsew signal output
rlabel metal2 s 326250 163200 326306 164000 6 la_iena[94]
port 190 nsew signal output
rlabel metal2 s 329746 163200 329802 164000 6 la_iena[95]
port 191 nsew signal output
rlabel metal2 s 333242 163200 333298 164000 6 la_iena[96]
port 192 nsew signal output
rlabel metal2 s 336646 163200 336702 164000 6 la_iena[97]
port 193 nsew signal output
rlabel metal2 s 340142 163200 340198 164000 6 la_iena[98]
port 194 nsew signal output
rlabel metal2 s 343638 163200 343694 164000 6 la_iena[99]
port 195 nsew signal output
rlabel metal2 s 31574 163200 31630 164000 6 la_iena[9]
port 196 nsew signal output
rlabel metal2 s 1214 163200 1270 164000 6 la_input[0]
port 197 nsew signal input
rlabel metal2 s 347962 163200 348018 164000 6 la_input[100]
port 198 nsew signal input
rlabel metal2 s 351366 163200 351422 164000 6 la_input[101]
port 199 nsew signal input
rlabel metal2 s 354862 163200 354918 164000 6 la_input[102]
port 200 nsew signal input
rlabel metal2 s 358358 163200 358414 164000 6 la_input[103]
port 201 nsew signal input
rlabel metal2 s 361854 163200 361910 164000 6 la_input[104]
port 202 nsew signal input
rlabel metal2 s 365258 163200 365314 164000 6 la_input[105]
port 203 nsew signal input
rlabel metal2 s 368754 163200 368810 164000 6 la_input[106]
port 204 nsew signal input
rlabel metal2 s 372250 163200 372306 164000 6 la_input[107]
port 205 nsew signal input
rlabel metal2 s 375654 163200 375710 164000 6 la_input[108]
port 206 nsew signal input
rlabel metal2 s 379150 163200 379206 164000 6 la_input[109]
port 207 nsew signal input
rlabel metal2 s 35898 163200 35954 164000 6 la_input[10]
port 208 nsew signal input
rlabel metal2 s 382646 163200 382702 164000 6 la_input[110]
port 209 nsew signal input
rlabel metal2 s 386050 163200 386106 164000 6 la_input[111]
port 210 nsew signal input
rlabel metal2 s 389546 163200 389602 164000 6 la_input[112]
port 211 nsew signal input
rlabel metal2 s 393042 163200 393098 164000 6 la_input[113]
port 212 nsew signal input
rlabel metal2 s 396446 163200 396502 164000 6 la_input[114]
port 213 nsew signal input
rlabel metal2 s 399942 163200 399998 164000 6 la_input[115]
port 214 nsew signal input
rlabel metal2 s 403438 163200 403494 164000 6 la_input[116]
port 215 nsew signal input
rlabel metal2 s 406842 163200 406898 164000 6 la_input[117]
port 216 nsew signal input
rlabel metal2 s 410338 163200 410394 164000 6 la_input[118]
port 217 nsew signal input
rlabel metal2 s 413834 163200 413890 164000 6 la_input[119]
port 218 nsew signal input
rlabel metal2 s 39302 163200 39358 164000 6 la_input[11]
port 219 nsew signal input
rlabel metal2 s 417330 163200 417386 164000 6 la_input[120]
port 220 nsew signal input
rlabel metal2 s 420734 163200 420790 164000 6 la_input[121]
port 221 nsew signal input
rlabel metal2 s 424230 163200 424286 164000 6 la_input[122]
port 222 nsew signal input
rlabel metal2 s 427726 163200 427782 164000 6 la_input[123]
port 223 nsew signal input
rlabel metal2 s 431130 163200 431186 164000 6 la_input[124]
port 224 nsew signal input
rlabel metal2 s 434626 163200 434682 164000 6 la_input[125]
port 225 nsew signal input
rlabel metal2 s 438122 163200 438178 164000 6 la_input[126]
port 226 nsew signal input
rlabel metal2 s 441526 163200 441582 164000 6 la_input[127]
port 227 nsew signal input
rlabel metal2 s 42798 163200 42854 164000 6 la_input[12]
port 228 nsew signal input
rlabel metal2 s 46294 163200 46350 164000 6 la_input[13]
port 229 nsew signal input
rlabel metal2 s 49790 163200 49846 164000 6 la_input[14]
port 230 nsew signal input
rlabel metal2 s 53194 163200 53250 164000 6 la_input[15]
port 231 nsew signal input
rlabel metal2 s 56690 163200 56746 164000 6 la_input[16]
port 232 nsew signal input
rlabel metal2 s 60186 163200 60242 164000 6 la_input[17]
port 233 nsew signal input
rlabel metal2 s 63590 163200 63646 164000 6 la_input[18]
port 234 nsew signal input
rlabel metal2 s 67086 163200 67142 164000 6 la_input[19]
port 235 nsew signal input
rlabel metal2 s 4710 163200 4766 164000 6 la_input[1]
port 236 nsew signal input
rlabel metal2 s 70582 163200 70638 164000 6 la_input[20]
port 237 nsew signal input
rlabel metal2 s 73986 163200 74042 164000 6 la_input[21]
port 238 nsew signal input
rlabel metal2 s 77482 163200 77538 164000 6 la_input[22]
port 239 nsew signal input
rlabel metal2 s 80978 163200 81034 164000 6 la_input[23]
port 240 nsew signal input
rlabel metal2 s 84382 163200 84438 164000 6 la_input[24]
port 241 nsew signal input
rlabel metal2 s 87878 163200 87934 164000 6 la_input[25]
port 242 nsew signal input
rlabel metal2 s 91374 163200 91430 164000 6 la_input[26]
port 243 nsew signal input
rlabel metal2 s 94870 163200 94926 164000 6 la_input[27]
port 244 nsew signal input
rlabel metal2 s 98274 163200 98330 164000 6 la_input[28]
port 245 nsew signal input
rlabel metal2 s 101770 163200 101826 164000 6 la_input[29]
port 246 nsew signal input
rlabel metal2 s 8114 163200 8170 164000 6 la_input[2]
port 247 nsew signal input
rlabel metal2 s 105266 163200 105322 164000 6 la_input[30]
port 248 nsew signal input
rlabel metal2 s 108670 163200 108726 164000 6 la_input[31]
port 249 nsew signal input
rlabel metal2 s 112166 163200 112222 164000 6 la_input[32]
port 250 nsew signal input
rlabel metal2 s 115662 163200 115718 164000 6 la_input[33]
port 251 nsew signal input
rlabel metal2 s 119066 163200 119122 164000 6 la_input[34]
port 252 nsew signal input
rlabel metal2 s 122562 163200 122618 164000 6 la_input[35]
port 253 nsew signal input
rlabel metal2 s 126058 163200 126114 164000 6 la_input[36]
port 254 nsew signal input
rlabel metal2 s 129462 163200 129518 164000 6 la_input[37]
port 255 nsew signal input
rlabel metal2 s 132958 163200 133014 164000 6 la_input[38]
port 256 nsew signal input
rlabel metal2 s 136454 163200 136510 164000 6 la_input[39]
port 257 nsew signal input
rlabel metal2 s 11610 163200 11666 164000 6 la_input[3]
port 258 nsew signal input
rlabel metal2 s 139858 163200 139914 164000 6 la_input[40]
port 259 nsew signal input
rlabel metal2 s 143354 163200 143410 164000 6 la_input[41]
port 260 nsew signal input
rlabel metal2 s 146850 163200 146906 164000 6 la_input[42]
port 261 nsew signal input
rlabel metal2 s 150346 163200 150402 164000 6 la_input[43]
port 262 nsew signal input
rlabel metal2 s 153750 163200 153806 164000 6 la_input[44]
port 263 nsew signal input
rlabel metal2 s 157246 163200 157302 164000 6 la_input[45]
port 264 nsew signal input
rlabel metal2 s 160742 163200 160798 164000 6 la_input[46]
port 265 nsew signal input
rlabel metal2 s 164146 163200 164202 164000 6 la_input[47]
port 266 nsew signal input
rlabel metal2 s 167642 163200 167698 164000 6 la_input[48]
port 267 nsew signal input
rlabel metal2 s 171138 163200 171194 164000 6 la_input[49]
port 268 nsew signal input
rlabel metal2 s 15106 163200 15162 164000 6 la_input[4]
port 269 nsew signal input
rlabel metal2 s 174542 163200 174598 164000 6 la_input[50]
port 270 nsew signal input
rlabel metal2 s 178038 163200 178094 164000 6 la_input[51]
port 271 nsew signal input
rlabel metal2 s 181534 163200 181590 164000 6 la_input[52]
port 272 nsew signal input
rlabel metal2 s 184938 163200 184994 164000 6 la_input[53]
port 273 nsew signal input
rlabel metal2 s 188434 163200 188490 164000 6 la_input[54]
port 274 nsew signal input
rlabel metal2 s 191930 163200 191986 164000 6 la_input[55]
port 275 nsew signal input
rlabel metal2 s 195334 163200 195390 164000 6 la_input[56]
port 276 nsew signal input
rlabel metal2 s 198830 163200 198886 164000 6 la_input[57]
port 277 nsew signal input
rlabel metal2 s 202326 163200 202382 164000 6 la_input[58]
port 278 nsew signal input
rlabel metal2 s 205822 163200 205878 164000 6 la_input[59]
port 279 nsew signal input
rlabel metal2 s 18510 163200 18566 164000 6 la_input[5]
port 280 nsew signal input
rlabel metal2 s 209226 163200 209282 164000 6 la_input[60]
port 281 nsew signal input
rlabel metal2 s 212722 163200 212778 164000 6 la_input[61]
port 282 nsew signal input
rlabel metal2 s 216218 163200 216274 164000 6 la_input[62]
port 283 nsew signal input
rlabel metal2 s 219622 163200 219678 164000 6 la_input[63]
port 284 nsew signal input
rlabel metal2 s 223118 163200 223174 164000 6 la_input[64]
port 285 nsew signal input
rlabel metal2 s 226614 163200 226670 164000 6 la_input[65]
port 286 nsew signal input
rlabel metal2 s 230018 163200 230074 164000 6 la_input[66]
port 287 nsew signal input
rlabel metal2 s 233514 163200 233570 164000 6 la_input[67]
port 288 nsew signal input
rlabel metal2 s 237010 163200 237066 164000 6 la_input[68]
port 289 nsew signal input
rlabel metal2 s 240414 163200 240470 164000 6 la_input[69]
port 290 nsew signal input
rlabel metal2 s 22006 163200 22062 164000 6 la_input[6]
port 291 nsew signal input
rlabel metal2 s 243910 163200 243966 164000 6 la_input[70]
port 292 nsew signal input
rlabel metal2 s 247406 163200 247462 164000 6 la_input[71]
port 293 nsew signal input
rlabel metal2 s 250902 163200 250958 164000 6 la_input[72]
port 294 nsew signal input
rlabel metal2 s 254306 163200 254362 164000 6 la_input[73]
port 295 nsew signal input
rlabel metal2 s 257802 163200 257858 164000 6 la_input[74]
port 296 nsew signal input
rlabel metal2 s 261298 163200 261354 164000 6 la_input[75]
port 297 nsew signal input
rlabel metal2 s 264702 163200 264758 164000 6 la_input[76]
port 298 nsew signal input
rlabel metal2 s 268198 163200 268254 164000 6 la_input[77]
port 299 nsew signal input
rlabel metal2 s 271694 163200 271750 164000 6 la_input[78]
port 300 nsew signal input
rlabel metal2 s 275098 163200 275154 164000 6 la_input[79]
port 301 nsew signal input
rlabel metal2 s 25502 163200 25558 164000 6 la_input[7]
port 302 nsew signal input
rlabel metal2 s 278594 163200 278650 164000 6 la_input[80]
port 303 nsew signal input
rlabel metal2 s 282090 163200 282146 164000 6 la_input[81]
port 304 nsew signal input
rlabel metal2 s 285494 163200 285550 164000 6 la_input[82]
port 305 nsew signal input
rlabel metal2 s 288990 163200 289046 164000 6 la_input[83]
port 306 nsew signal input
rlabel metal2 s 292486 163200 292542 164000 6 la_input[84]
port 307 nsew signal input
rlabel metal2 s 295890 163200 295946 164000 6 la_input[85]
port 308 nsew signal input
rlabel metal2 s 299386 163200 299442 164000 6 la_input[86]
port 309 nsew signal input
rlabel metal2 s 302882 163200 302938 164000 6 la_input[87]
port 310 nsew signal input
rlabel metal2 s 306378 163200 306434 164000 6 la_input[88]
port 311 nsew signal input
rlabel metal2 s 309782 163200 309838 164000 6 la_input[89]
port 312 nsew signal input
rlabel metal2 s 28906 163200 28962 164000 6 la_input[8]
port 313 nsew signal input
rlabel metal2 s 313278 163200 313334 164000 6 la_input[90]
port 314 nsew signal input
rlabel metal2 s 316774 163200 316830 164000 6 la_input[91]
port 315 nsew signal input
rlabel metal2 s 320178 163200 320234 164000 6 la_input[92]
port 316 nsew signal input
rlabel metal2 s 323674 163200 323730 164000 6 la_input[93]
port 317 nsew signal input
rlabel metal2 s 327170 163200 327226 164000 6 la_input[94]
port 318 nsew signal input
rlabel metal2 s 330574 163200 330630 164000 6 la_input[95]
port 319 nsew signal input
rlabel metal2 s 334070 163200 334126 164000 6 la_input[96]
port 320 nsew signal input
rlabel metal2 s 337566 163200 337622 164000 6 la_input[97]
port 321 nsew signal input
rlabel metal2 s 340970 163200 341026 164000 6 la_input[98]
port 322 nsew signal input
rlabel metal2 s 344466 163200 344522 164000 6 la_input[99]
port 323 nsew signal input
rlabel metal2 s 32402 163200 32458 164000 6 la_input[9]
port 324 nsew signal input
rlabel metal2 s 2042 163200 2098 164000 6 la_oenb[0]
port 325 nsew signal output
rlabel metal2 s 348790 163200 348846 164000 6 la_oenb[100]
port 326 nsew signal output
rlabel metal2 s 352286 163200 352342 164000 6 la_oenb[101]
port 327 nsew signal output
rlabel metal2 s 355782 163200 355838 164000 6 la_oenb[102]
port 328 nsew signal output
rlabel metal2 s 359186 163200 359242 164000 6 la_oenb[103]
port 329 nsew signal output
rlabel metal2 s 362682 163200 362738 164000 6 la_oenb[104]
port 330 nsew signal output
rlabel metal2 s 366178 163200 366234 164000 6 la_oenb[105]
port 331 nsew signal output
rlabel metal2 s 369582 163200 369638 164000 6 la_oenb[106]
port 332 nsew signal output
rlabel metal2 s 373078 163200 373134 164000 6 la_oenb[107]
port 333 nsew signal output
rlabel metal2 s 376574 163200 376630 164000 6 la_oenb[108]
port 334 nsew signal output
rlabel metal2 s 379978 163200 380034 164000 6 la_oenb[109]
port 335 nsew signal output
rlabel metal2 s 36726 163200 36782 164000 6 la_oenb[10]
port 336 nsew signal output
rlabel metal2 s 383474 163200 383530 164000 6 la_oenb[110]
port 337 nsew signal output
rlabel metal2 s 386970 163200 387026 164000 6 la_oenb[111]
port 338 nsew signal output
rlabel metal2 s 390374 163200 390430 164000 6 la_oenb[112]
port 339 nsew signal output
rlabel metal2 s 393870 163200 393926 164000 6 la_oenb[113]
port 340 nsew signal output
rlabel metal2 s 397366 163200 397422 164000 6 la_oenb[114]
port 341 nsew signal output
rlabel metal2 s 400862 163200 400918 164000 6 la_oenb[115]
port 342 nsew signal output
rlabel metal2 s 404266 163200 404322 164000 6 la_oenb[116]
port 343 nsew signal output
rlabel metal2 s 407762 163200 407818 164000 6 la_oenb[117]
port 344 nsew signal output
rlabel metal2 s 411258 163200 411314 164000 6 la_oenb[118]
port 345 nsew signal output
rlabel metal2 s 414662 163200 414718 164000 6 la_oenb[119]
port 346 nsew signal output
rlabel metal2 s 40222 163200 40278 164000 6 la_oenb[11]
port 347 nsew signal output
rlabel metal2 s 418158 163200 418214 164000 6 la_oenb[120]
port 348 nsew signal output
rlabel metal2 s 421654 163200 421710 164000 6 la_oenb[121]
port 349 nsew signal output
rlabel metal2 s 425058 163200 425114 164000 6 la_oenb[122]
port 350 nsew signal output
rlabel metal2 s 428554 163200 428610 164000 6 la_oenb[123]
port 351 nsew signal output
rlabel metal2 s 432050 163200 432106 164000 6 la_oenb[124]
port 352 nsew signal output
rlabel metal2 s 435454 163200 435510 164000 6 la_oenb[125]
port 353 nsew signal output
rlabel metal2 s 438950 163200 439006 164000 6 la_oenb[126]
port 354 nsew signal output
rlabel metal2 s 442446 163200 442502 164000 6 la_oenb[127]
port 355 nsew signal output
rlabel metal2 s 43718 163200 43774 164000 6 la_oenb[12]
port 356 nsew signal output
rlabel metal2 s 47122 163200 47178 164000 6 la_oenb[13]
port 357 nsew signal output
rlabel metal2 s 50618 163200 50674 164000 6 la_oenb[14]
port 358 nsew signal output
rlabel metal2 s 54114 163200 54170 164000 6 la_oenb[15]
port 359 nsew signal output
rlabel metal2 s 57518 163200 57574 164000 6 la_oenb[16]
port 360 nsew signal output
rlabel metal2 s 61014 163200 61070 164000 6 la_oenb[17]
port 361 nsew signal output
rlabel metal2 s 64510 163200 64566 164000 6 la_oenb[18]
port 362 nsew signal output
rlabel metal2 s 67914 163200 67970 164000 6 la_oenb[19]
port 363 nsew signal output
rlabel metal2 s 5538 163200 5594 164000 6 la_oenb[1]
port 364 nsew signal output
rlabel metal2 s 71410 163200 71466 164000 6 la_oenb[20]
port 365 nsew signal output
rlabel metal2 s 74906 163200 74962 164000 6 la_oenb[21]
port 366 nsew signal output
rlabel metal2 s 78310 163200 78366 164000 6 la_oenb[22]
port 367 nsew signal output
rlabel metal2 s 81806 163200 81862 164000 6 la_oenb[23]
port 368 nsew signal output
rlabel metal2 s 85302 163200 85358 164000 6 la_oenb[24]
port 369 nsew signal output
rlabel metal2 s 88798 163200 88854 164000 6 la_oenb[25]
port 370 nsew signal output
rlabel metal2 s 92202 163200 92258 164000 6 la_oenb[26]
port 371 nsew signal output
rlabel metal2 s 95698 163200 95754 164000 6 la_oenb[27]
port 372 nsew signal output
rlabel metal2 s 99194 163200 99250 164000 6 la_oenb[28]
port 373 nsew signal output
rlabel metal2 s 102598 163200 102654 164000 6 la_oenb[29]
port 374 nsew signal output
rlabel metal2 s 9034 163200 9090 164000 6 la_oenb[2]
port 375 nsew signal output
rlabel metal2 s 106094 163200 106150 164000 6 la_oenb[30]
port 376 nsew signal output
rlabel metal2 s 109590 163200 109646 164000 6 la_oenb[31]
port 377 nsew signal output
rlabel metal2 s 112994 163200 113050 164000 6 la_oenb[32]
port 378 nsew signal output
rlabel metal2 s 116490 163200 116546 164000 6 la_oenb[33]
port 379 nsew signal output
rlabel metal2 s 119986 163200 120042 164000 6 la_oenb[34]
port 380 nsew signal output
rlabel metal2 s 123390 163200 123446 164000 6 la_oenb[35]
port 381 nsew signal output
rlabel metal2 s 126886 163200 126942 164000 6 la_oenb[36]
port 382 nsew signal output
rlabel metal2 s 130382 163200 130438 164000 6 la_oenb[37]
port 383 nsew signal output
rlabel metal2 s 133878 163200 133934 164000 6 la_oenb[38]
port 384 nsew signal output
rlabel metal2 s 137282 163200 137338 164000 6 la_oenb[39]
port 385 nsew signal output
rlabel metal2 s 12438 163200 12494 164000 6 la_oenb[3]
port 386 nsew signal output
rlabel metal2 s 140778 163200 140834 164000 6 la_oenb[40]
port 387 nsew signal output
rlabel metal2 s 144274 163200 144330 164000 6 la_oenb[41]
port 388 nsew signal output
rlabel metal2 s 147678 163200 147734 164000 6 la_oenb[42]
port 389 nsew signal output
rlabel metal2 s 151174 163200 151230 164000 6 la_oenb[43]
port 390 nsew signal output
rlabel metal2 s 154670 163200 154726 164000 6 la_oenb[44]
port 391 nsew signal output
rlabel metal2 s 158074 163200 158130 164000 6 la_oenb[45]
port 392 nsew signal output
rlabel metal2 s 161570 163200 161626 164000 6 la_oenb[46]
port 393 nsew signal output
rlabel metal2 s 165066 163200 165122 164000 6 la_oenb[47]
port 394 nsew signal output
rlabel metal2 s 168470 163200 168526 164000 6 la_oenb[48]
port 395 nsew signal output
rlabel metal2 s 171966 163200 172022 164000 6 la_oenb[49]
port 396 nsew signal output
rlabel metal2 s 15934 163200 15990 164000 6 la_oenb[4]
port 397 nsew signal output
rlabel metal2 s 175462 163200 175518 164000 6 la_oenb[50]
port 398 nsew signal output
rlabel metal2 s 178866 163200 178922 164000 6 la_oenb[51]
port 399 nsew signal output
rlabel metal2 s 182362 163200 182418 164000 6 la_oenb[52]
port 400 nsew signal output
rlabel metal2 s 185858 163200 185914 164000 6 la_oenb[53]
port 401 nsew signal output
rlabel metal2 s 189354 163200 189410 164000 6 la_oenb[54]
port 402 nsew signal output
rlabel metal2 s 192758 163200 192814 164000 6 la_oenb[55]
port 403 nsew signal output
rlabel metal2 s 196254 163200 196310 164000 6 la_oenb[56]
port 404 nsew signal output
rlabel metal2 s 199750 163200 199806 164000 6 la_oenb[57]
port 405 nsew signal output
rlabel metal2 s 203154 163200 203210 164000 6 la_oenb[58]
port 406 nsew signal output
rlabel metal2 s 206650 163200 206706 164000 6 la_oenb[59]
port 407 nsew signal output
rlabel metal2 s 19430 163200 19486 164000 6 la_oenb[5]
port 408 nsew signal output
rlabel metal2 s 210146 163200 210202 164000 6 la_oenb[60]
port 409 nsew signal output
rlabel metal2 s 213550 163200 213606 164000 6 la_oenb[61]
port 410 nsew signal output
rlabel metal2 s 217046 163200 217102 164000 6 la_oenb[62]
port 411 nsew signal output
rlabel metal2 s 220542 163200 220598 164000 6 la_oenb[63]
port 412 nsew signal output
rlabel metal2 s 223946 163200 224002 164000 6 la_oenb[64]
port 413 nsew signal output
rlabel metal2 s 227442 163200 227498 164000 6 la_oenb[65]
port 414 nsew signal output
rlabel metal2 s 230938 163200 230994 164000 6 la_oenb[66]
port 415 nsew signal output
rlabel metal2 s 234342 163200 234398 164000 6 la_oenb[67]
port 416 nsew signal output
rlabel metal2 s 237838 163200 237894 164000 6 la_oenb[68]
port 417 nsew signal output
rlabel metal2 s 241334 163200 241390 164000 6 la_oenb[69]
port 418 nsew signal output
rlabel metal2 s 22834 163200 22890 164000 6 la_oenb[6]
port 419 nsew signal output
rlabel metal2 s 244830 163200 244886 164000 6 la_oenb[70]
port 420 nsew signal output
rlabel metal2 s 248234 163200 248290 164000 6 la_oenb[71]
port 421 nsew signal output
rlabel metal2 s 251730 163200 251786 164000 6 la_oenb[72]
port 422 nsew signal output
rlabel metal2 s 255226 163200 255282 164000 6 la_oenb[73]
port 423 nsew signal output
rlabel metal2 s 258630 163200 258686 164000 6 la_oenb[74]
port 424 nsew signal output
rlabel metal2 s 262126 163200 262182 164000 6 la_oenb[75]
port 425 nsew signal output
rlabel metal2 s 265622 163200 265678 164000 6 la_oenb[76]
port 426 nsew signal output
rlabel metal2 s 269026 163200 269082 164000 6 la_oenb[77]
port 427 nsew signal output
rlabel metal2 s 272522 163200 272578 164000 6 la_oenb[78]
port 428 nsew signal output
rlabel metal2 s 276018 163200 276074 164000 6 la_oenb[79]
port 429 nsew signal output
rlabel metal2 s 26330 163200 26386 164000 6 la_oenb[7]
port 430 nsew signal output
rlabel metal2 s 279422 163200 279478 164000 6 la_oenb[80]
port 431 nsew signal output
rlabel metal2 s 282918 163200 282974 164000 6 la_oenb[81]
port 432 nsew signal output
rlabel metal2 s 286414 163200 286470 164000 6 la_oenb[82]
port 433 nsew signal output
rlabel metal2 s 289818 163200 289874 164000 6 la_oenb[83]
port 434 nsew signal output
rlabel metal2 s 293314 163200 293370 164000 6 la_oenb[84]
port 435 nsew signal output
rlabel metal2 s 296810 163200 296866 164000 6 la_oenb[85]
port 436 nsew signal output
rlabel metal2 s 300306 163200 300362 164000 6 la_oenb[86]
port 437 nsew signal output
rlabel metal2 s 303710 163200 303766 164000 6 la_oenb[87]
port 438 nsew signal output
rlabel metal2 s 307206 163200 307262 164000 6 la_oenb[88]
port 439 nsew signal output
rlabel metal2 s 310702 163200 310758 164000 6 la_oenb[89]
port 440 nsew signal output
rlabel metal2 s 29826 163200 29882 164000 6 la_oenb[8]
port 441 nsew signal output
rlabel metal2 s 314106 163200 314162 164000 6 la_oenb[90]
port 442 nsew signal output
rlabel metal2 s 317602 163200 317658 164000 6 la_oenb[91]
port 443 nsew signal output
rlabel metal2 s 321098 163200 321154 164000 6 la_oenb[92]
port 444 nsew signal output
rlabel metal2 s 324502 163200 324558 164000 6 la_oenb[93]
port 445 nsew signal output
rlabel metal2 s 327998 163200 328054 164000 6 la_oenb[94]
port 446 nsew signal output
rlabel metal2 s 331494 163200 331550 164000 6 la_oenb[95]
port 447 nsew signal output
rlabel metal2 s 334898 163200 334954 164000 6 la_oenb[96]
port 448 nsew signal output
rlabel metal2 s 338394 163200 338450 164000 6 la_oenb[97]
port 449 nsew signal output
rlabel metal2 s 341890 163200 341946 164000 6 la_oenb[98]
port 450 nsew signal output
rlabel metal2 s 345386 163200 345442 164000 6 la_oenb[99]
port 451 nsew signal output
rlabel metal2 s 33322 163200 33378 164000 6 la_oenb[9]
port 452 nsew signal output
rlabel metal2 s 2962 163200 3018 164000 6 la_output[0]
port 453 nsew signal output
rlabel metal2 s 349710 163200 349766 164000 6 la_output[100]
port 454 nsew signal output
rlabel metal2 s 353114 163200 353170 164000 6 la_output[101]
port 455 nsew signal output
rlabel metal2 s 356610 163200 356666 164000 6 la_output[102]
port 456 nsew signal output
rlabel metal2 s 360106 163200 360162 164000 6 la_output[103]
port 457 nsew signal output
rlabel metal2 s 363510 163200 363566 164000 6 la_output[104]
port 458 nsew signal output
rlabel metal2 s 367006 163200 367062 164000 6 la_output[105]
port 459 nsew signal output
rlabel metal2 s 370502 163200 370558 164000 6 la_output[106]
port 460 nsew signal output
rlabel metal2 s 373906 163200 373962 164000 6 la_output[107]
port 461 nsew signal output
rlabel metal2 s 377402 163200 377458 164000 6 la_output[108]
port 462 nsew signal output
rlabel metal2 s 380898 163200 380954 164000 6 la_output[109]
port 463 nsew signal output
rlabel metal2 s 37646 163200 37702 164000 6 la_output[10]
port 464 nsew signal output
rlabel metal2 s 384394 163200 384450 164000 6 la_output[110]
port 465 nsew signal output
rlabel metal2 s 387798 163200 387854 164000 6 la_output[111]
port 466 nsew signal output
rlabel metal2 s 391294 163200 391350 164000 6 la_output[112]
port 467 nsew signal output
rlabel metal2 s 394790 163200 394846 164000 6 la_output[113]
port 468 nsew signal output
rlabel metal2 s 398194 163200 398250 164000 6 la_output[114]
port 469 nsew signal output
rlabel metal2 s 401690 163200 401746 164000 6 la_output[115]
port 470 nsew signal output
rlabel metal2 s 405186 163200 405242 164000 6 la_output[116]
port 471 nsew signal output
rlabel metal2 s 408590 163200 408646 164000 6 la_output[117]
port 472 nsew signal output
rlabel metal2 s 412086 163200 412142 164000 6 la_output[118]
port 473 nsew signal output
rlabel metal2 s 415582 163200 415638 164000 6 la_output[119]
port 474 nsew signal output
rlabel metal2 s 41050 163200 41106 164000 6 la_output[11]
port 475 nsew signal output
rlabel metal2 s 418986 163200 419042 164000 6 la_output[120]
port 476 nsew signal output
rlabel metal2 s 422482 163200 422538 164000 6 la_output[121]
port 477 nsew signal output
rlabel metal2 s 425978 163200 426034 164000 6 la_output[122]
port 478 nsew signal output
rlabel metal2 s 429382 163200 429438 164000 6 la_output[123]
port 479 nsew signal output
rlabel metal2 s 432878 163200 432934 164000 6 la_output[124]
port 480 nsew signal output
rlabel metal2 s 436374 163200 436430 164000 6 la_output[125]
port 481 nsew signal output
rlabel metal2 s 439870 163200 439926 164000 6 la_output[126]
port 482 nsew signal output
rlabel metal2 s 443274 163200 443330 164000 6 la_output[127]
port 483 nsew signal output
rlabel metal2 s 44546 163200 44602 164000 6 la_output[12]
port 484 nsew signal output
rlabel metal2 s 48042 163200 48098 164000 6 la_output[13]
port 485 nsew signal output
rlabel metal2 s 51446 163200 51502 164000 6 la_output[14]
port 486 nsew signal output
rlabel metal2 s 54942 163200 54998 164000 6 la_output[15]
port 487 nsew signal output
rlabel metal2 s 58438 163200 58494 164000 6 la_output[16]
port 488 nsew signal output
rlabel metal2 s 61842 163200 61898 164000 6 la_output[17]
port 489 nsew signal output
rlabel metal2 s 65338 163200 65394 164000 6 la_output[18]
port 490 nsew signal output
rlabel metal2 s 68834 163200 68890 164000 6 la_output[19]
port 491 nsew signal output
rlabel metal2 s 6366 163200 6422 164000 6 la_output[1]
port 492 nsew signal output
rlabel metal2 s 72330 163200 72386 164000 6 la_output[20]
port 493 nsew signal output
rlabel metal2 s 75734 163200 75790 164000 6 la_output[21]
port 494 nsew signal output
rlabel metal2 s 79230 163200 79286 164000 6 la_output[22]
port 495 nsew signal output
rlabel metal2 s 82726 163200 82782 164000 6 la_output[23]
port 496 nsew signal output
rlabel metal2 s 86130 163200 86186 164000 6 la_output[24]
port 497 nsew signal output
rlabel metal2 s 89626 163200 89682 164000 6 la_output[25]
port 498 nsew signal output
rlabel metal2 s 93122 163200 93178 164000 6 la_output[26]
port 499 nsew signal output
rlabel metal2 s 96526 163200 96582 164000 6 la_output[27]
port 500 nsew signal output
rlabel metal2 s 100022 163200 100078 164000 6 la_output[28]
port 501 nsew signal output
rlabel metal2 s 103518 163200 103574 164000 6 la_output[29]
port 502 nsew signal output
rlabel metal2 s 9862 163200 9918 164000 6 la_output[2]
port 503 nsew signal output
rlabel metal2 s 106922 163200 106978 164000 6 la_output[30]
port 504 nsew signal output
rlabel metal2 s 110418 163200 110474 164000 6 la_output[31]
port 505 nsew signal output
rlabel metal2 s 113914 163200 113970 164000 6 la_output[32]
port 506 nsew signal output
rlabel metal2 s 117318 163200 117374 164000 6 la_output[33]
port 507 nsew signal output
rlabel metal2 s 120814 163200 120870 164000 6 la_output[34]
port 508 nsew signal output
rlabel metal2 s 124310 163200 124366 164000 6 la_output[35]
port 509 nsew signal output
rlabel metal2 s 127806 163200 127862 164000 6 la_output[36]
port 510 nsew signal output
rlabel metal2 s 131210 163200 131266 164000 6 la_output[37]
port 511 nsew signal output
rlabel metal2 s 134706 163200 134762 164000 6 la_output[38]
port 512 nsew signal output
rlabel metal2 s 138202 163200 138258 164000 6 la_output[39]
port 513 nsew signal output
rlabel metal2 s 13358 163200 13414 164000 6 la_output[3]
port 514 nsew signal output
rlabel metal2 s 141606 163200 141662 164000 6 la_output[40]
port 515 nsew signal output
rlabel metal2 s 145102 163200 145158 164000 6 la_output[41]
port 516 nsew signal output
rlabel metal2 s 148598 163200 148654 164000 6 la_output[42]
port 517 nsew signal output
rlabel metal2 s 152002 163200 152058 164000 6 la_output[43]
port 518 nsew signal output
rlabel metal2 s 155498 163200 155554 164000 6 la_output[44]
port 519 nsew signal output
rlabel metal2 s 158994 163200 159050 164000 6 la_output[45]
port 520 nsew signal output
rlabel metal2 s 162398 163200 162454 164000 6 la_output[46]
port 521 nsew signal output
rlabel metal2 s 165894 163200 165950 164000 6 la_output[47]
port 522 nsew signal output
rlabel metal2 s 169390 163200 169446 164000 6 la_output[48]
port 523 nsew signal output
rlabel metal2 s 172886 163200 172942 164000 6 la_output[49]
port 524 nsew signal output
rlabel metal2 s 16854 163200 16910 164000 6 la_output[4]
port 525 nsew signal output
rlabel metal2 s 176290 163200 176346 164000 6 la_output[50]
port 526 nsew signal output
rlabel metal2 s 179786 163200 179842 164000 6 la_output[51]
port 527 nsew signal output
rlabel metal2 s 183282 163200 183338 164000 6 la_output[52]
port 528 nsew signal output
rlabel metal2 s 186686 163200 186742 164000 6 la_output[53]
port 529 nsew signal output
rlabel metal2 s 190182 163200 190238 164000 6 la_output[54]
port 530 nsew signal output
rlabel metal2 s 193678 163200 193734 164000 6 la_output[55]
port 531 nsew signal output
rlabel metal2 s 197082 163200 197138 164000 6 la_output[56]
port 532 nsew signal output
rlabel metal2 s 200578 163200 200634 164000 6 la_output[57]
port 533 nsew signal output
rlabel metal2 s 204074 163200 204130 164000 6 la_output[58]
port 534 nsew signal output
rlabel metal2 s 207478 163200 207534 164000 6 la_output[59]
port 535 nsew signal output
rlabel metal2 s 20258 163200 20314 164000 6 la_output[5]
port 536 nsew signal output
rlabel metal2 s 210974 163200 211030 164000 6 la_output[60]
port 537 nsew signal output
rlabel metal2 s 214470 163200 214526 164000 6 la_output[61]
port 538 nsew signal output
rlabel metal2 s 217874 163200 217930 164000 6 la_output[62]
port 539 nsew signal output
rlabel metal2 s 221370 163200 221426 164000 6 la_output[63]
port 540 nsew signal output
rlabel metal2 s 224866 163200 224922 164000 6 la_output[64]
port 541 nsew signal output
rlabel metal2 s 228362 163200 228418 164000 6 la_output[65]
port 542 nsew signal output
rlabel metal2 s 231766 163200 231822 164000 6 la_output[66]
port 543 nsew signal output
rlabel metal2 s 235262 163200 235318 164000 6 la_output[67]
port 544 nsew signal output
rlabel metal2 s 238758 163200 238814 164000 6 la_output[68]
port 545 nsew signal output
rlabel metal2 s 242162 163200 242218 164000 6 la_output[69]
port 546 nsew signal output
rlabel metal2 s 23754 163200 23810 164000 6 la_output[6]
port 547 nsew signal output
rlabel metal2 s 245658 163200 245714 164000 6 la_output[70]
port 548 nsew signal output
rlabel metal2 s 249154 163200 249210 164000 6 la_output[71]
port 549 nsew signal output
rlabel metal2 s 252558 163200 252614 164000 6 la_output[72]
port 550 nsew signal output
rlabel metal2 s 256054 163200 256110 164000 6 la_output[73]
port 551 nsew signal output
rlabel metal2 s 259550 163200 259606 164000 6 la_output[74]
port 552 nsew signal output
rlabel metal2 s 262954 163200 263010 164000 6 la_output[75]
port 553 nsew signal output
rlabel metal2 s 266450 163200 266506 164000 6 la_output[76]
port 554 nsew signal output
rlabel metal2 s 269946 163200 270002 164000 6 la_output[77]
port 555 nsew signal output
rlabel metal2 s 273350 163200 273406 164000 6 la_output[78]
port 556 nsew signal output
rlabel metal2 s 276846 163200 276902 164000 6 la_output[79]
port 557 nsew signal output
rlabel metal2 s 27250 163200 27306 164000 6 la_output[7]
port 558 nsew signal output
rlabel metal2 s 280342 163200 280398 164000 6 la_output[80]
port 559 nsew signal output
rlabel metal2 s 283838 163200 283894 164000 6 la_output[81]
port 560 nsew signal output
rlabel metal2 s 287242 163200 287298 164000 6 la_output[82]
port 561 nsew signal output
rlabel metal2 s 290738 163200 290794 164000 6 la_output[83]
port 562 nsew signal output
rlabel metal2 s 294234 163200 294290 164000 6 la_output[84]
port 563 nsew signal output
rlabel metal2 s 297638 163200 297694 164000 6 la_output[85]
port 564 nsew signal output
rlabel metal2 s 301134 163200 301190 164000 6 la_output[86]
port 565 nsew signal output
rlabel metal2 s 304630 163200 304686 164000 6 la_output[87]
port 566 nsew signal output
rlabel metal2 s 308034 163200 308090 164000 6 la_output[88]
port 567 nsew signal output
rlabel metal2 s 311530 163200 311586 164000 6 la_output[89]
port 568 nsew signal output
rlabel metal2 s 30654 163200 30710 164000 6 la_output[8]
port 569 nsew signal output
rlabel metal2 s 315026 163200 315082 164000 6 la_output[90]
port 570 nsew signal output
rlabel metal2 s 318430 163200 318486 164000 6 la_output[91]
port 571 nsew signal output
rlabel metal2 s 321926 163200 321982 164000 6 la_output[92]
port 572 nsew signal output
rlabel metal2 s 325422 163200 325478 164000 6 la_output[93]
port 573 nsew signal output
rlabel metal2 s 328826 163200 328882 164000 6 la_output[94]
port 574 nsew signal output
rlabel metal2 s 332322 163200 332378 164000 6 la_output[95]
port 575 nsew signal output
rlabel metal2 s 335818 163200 335874 164000 6 la_output[96]
port 576 nsew signal output
rlabel metal2 s 339314 163200 339370 164000 6 la_output[97]
port 577 nsew signal output
rlabel metal2 s 342718 163200 342774 164000 6 la_output[98]
port 578 nsew signal output
rlabel metal2 s 346214 163200 346270 164000 6 la_output[99]
port 579 nsew signal output
rlabel metal2 s 34150 163200 34206 164000 6 la_output[9]
port 580 nsew signal output
rlabel metal2 s 444194 163200 444250 164000 6 mprj_ack_i
port 581 nsew signal input
rlabel metal2 s 448518 163200 448574 164000 6 mprj_adr_o[0]
port 582 nsew signal output
rlabel metal2 s 477958 163200 478014 164000 6 mprj_adr_o[10]
port 583 nsew signal output
rlabel metal2 s 480534 163200 480590 164000 6 mprj_adr_o[11]
port 584 nsew signal output
rlabel metal2 s 483202 163200 483258 164000 6 mprj_adr_o[12]
port 585 nsew signal output
rlabel metal2 s 485778 163200 485834 164000 6 mprj_adr_o[13]
port 586 nsew signal output
rlabel metal2 s 488354 163200 488410 164000 6 mprj_adr_o[14]
port 587 nsew signal output
rlabel metal2 s 490930 163200 490986 164000 6 mprj_adr_o[15]
port 588 nsew signal output
rlabel metal2 s 493598 163200 493654 164000 6 mprj_adr_o[16]
port 589 nsew signal output
rlabel metal2 s 496174 163200 496230 164000 6 mprj_adr_o[17]
port 590 nsew signal output
rlabel metal2 s 498750 163200 498806 164000 6 mprj_adr_o[18]
port 591 nsew signal output
rlabel metal2 s 501418 163200 501474 164000 6 mprj_adr_o[19]
port 592 nsew signal output
rlabel metal2 s 451922 163200 451978 164000 6 mprj_adr_o[1]
port 593 nsew signal output
rlabel metal2 s 503994 163200 504050 164000 6 mprj_adr_o[20]
port 594 nsew signal output
rlabel metal2 s 506570 163200 506626 164000 6 mprj_adr_o[21]
port 595 nsew signal output
rlabel metal2 s 509146 163200 509202 164000 6 mprj_adr_o[22]
port 596 nsew signal output
rlabel metal2 s 511814 163200 511870 164000 6 mprj_adr_o[23]
port 597 nsew signal output
rlabel metal2 s 514390 163200 514446 164000 6 mprj_adr_o[24]
port 598 nsew signal output
rlabel metal2 s 516966 163200 517022 164000 6 mprj_adr_o[25]
port 599 nsew signal output
rlabel metal2 s 519542 163200 519598 164000 6 mprj_adr_o[26]
port 600 nsew signal output
rlabel metal2 s 522210 163200 522266 164000 6 mprj_adr_o[27]
port 601 nsew signal output
rlabel metal2 s 524786 163200 524842 164000 6 mprj_adr_o[28]
port 602 nsew signal output
rlabel metal2 s 527362 163200 527418 164000 6 mprj_adr_o[29]
port 603 nsew signal output
rlabel metal2 s 455418 163200 455474 164000 6 mprj_adr_o[2]
port 604 nsew signal output
rlabel metal2 s 529938 163200 529994 164000 6 mprj_adr_o[30]
port 605 nsew signal output
rlabel metal2 s 532606 163200 532662 164000 6 mprj_adr_o[31]
port 606 nsew signal output
rlabel metal2 s 458914 163200 458970 164000 6 mprj_adr_o[3]
port 607 nsew signal output
rlabel metal2 s 462410 163200 462466 164000 6 mprj_adr_o[4]
port 608 nsew signal output
rlabel metal2 s 464986 163200 465042 164000 6 mprj_adr_o[5]
port 609 nsew signal output
rlabel metal2 s 467562 163200 467618 164000 6 mprj_adr_o[6]
port 610 nsew signal output
rlabel metal2 s 470138 163200 470194 164000 6 mprj_adr_o[7]
port 611 nsew signal output
rlabel metal2 s 472806 163200 472862 164000 6 mprj_adr_o[8]
port 612 nsew signal output
rlabel metal2 s 475382 163200 475438 164000 6 mprj_adr_o[9]
port 613 nsew signal output
rlabel metal2 s 445022 163200 445078 164000 6 mprj_cyc_o
port 614 nsew signal output
rlabel metal2 s 449346 163200 449402 164000 6 mprj_dat_i[0]
port 615 nsew signal input
rlabel metal2 s 478878 163200 478934 164000 6 mprj_dat_i[10]
port 616 nsew signal input
rlabel metal2 s 481454 163200 481510 164000 6 mprj_dat_i[11]
port 617 nsew signal input
rlabel metal2 s 484030 163200 484086 164000 6 mprj_dat_i[12]
port 618 nsew signal input
rlabel metal2 s 486606 163200 486662 164000 6 mprj_dat_i[13]
port 619 nsew signal input
rlabel metal2 s 489274 163200 489330 164000 6 mprj_dat_i[14]
port 620 nsew signal input
rlabel metal2 s 491850 163200 491906 164000 6 mprj_dat_i[15]
port 621 nsew signal input
rlabel metal2 s 494426 163200 494482 164000 6 mprj_dat_i[16]
port 622 nsew signal input
rlabel metal2 s 497002 163200 497058 164000 6 mprj_dat_i[17]
port 623 nsew signal input
rlabel metal2 s 499670 163200 499726 164000 6 mprj_dat_i[18]
port 624 nsew signal input
rlabel metal2 s 502246 163200 502302 164000 6 mprj_dat_i[19]
port 625 nsew signal input
rlabel metal2 s 452842 163200 452898 164000 6 mprj_dat_i[1]
port 626 nsew signal input
rlabel metal2 s 504822 163200 504878 164000 6 mprj_dat_i[20]
port 627 nsew signal input
rlabel metal2 s 507398 163200 507454 164000 6 mprj_dat_i[21]
port 628 nsew signal input
rlabel metal2 s 510066 163200 510122 164000 6 mprj_dat_i[22]
port 629 nsew signal input
rlabel metal2 s 512642 163200 512698 164000 6 mprj_dat_i[23]
port 630 nsew signal input
rlabel metal2 s 515218 163200 515274 164000 6 mprj_dat_i[24]
port 631 nsew signal input
rlabel metal2 s 517886 163200 517942 164000 6 mprj_dat_i[25]
port 632 nsew signal input
rlabel metal2 s 520462 163200 520518 164000 6 mprj_dat_i[26]
port 633 nsew signal input
rlabel metal2 s 523038 163200 523094 164000 6 mprj_dat_i[27]
port 634 nsew signal input
rlabel metal2 s 525614 163200 525670 164000 6 mprj_dat_i[28]
port 635 nsew signal input
rlabel metal2 s 528282 163200 528338 164000 6 mprj_dat_i[29]
port 636 nsew signal input
rlabel metal2 s 456338 163200 456394 164000 6 mprj_dat_i[2]
port 637 nsew signal input
rlabel metal2 s 530858 163200 530914 164000 6 mprj_dat_i[30]
port 638 nsew signal input
rlabel metal2 s 533434 163200 533490 164000 6 mprj_dat_i[31]
port 639 nsew signal input
rlabel metal2 s 459742 163200 459798 164000 6 mprj_dat_i[3]
port 640 nsew signal input
rlabel metal2 s 463238 163200 463294 164000 6 mprj_dat_i[4]
port 641 nsew signal input
rlabel metal2 s 465814 163200 465870 164000 6 mprj_dat_i[5]
port 642 nsew signal input
rlabel metal2 s 468390 163200 468446 164000 6 mprj_dat_i[6]
port 643 nsew signal input
rlabel metal2 s 471058 163200 471114 164000 6 mprj_dat_i[7]
port 644 nsew signal input
rlabel metal2 s 473634 163200 473690 164000 6 mprj_dat_i[8]
port 645 nsew signal input
rlabel metal2 s 476210 163200 476266 164000 6 mprj_dat_i[9]
port 646 nsew signal input
rlabel metal2 s 450266 163200 450322 164000 6 mprj_dat_o[0]
port 647 nsew signal output
rlabel metal2 s 479706 163200 479762 164000 6 mprj_dat_o[10]
port 648 nsew signal output
rlabel metal2 s 482282 163200 482338 164000 6 mprj_dat_o[11]
port 649 nsew signal output
rlabel metal2 s 484858 163200 484914 164000 6 mprj_dat_o[12]
port 650 nsew signal output
rlabel metal2 s 487526 163200 487582 164000 6 mprj_dat_o[13]
port 651 nsew signal output
rlabel metal2 s 490102 163200 490158 164000 6 mprj_dat_o[14]
port 652 nsew signal output
rlabel metal2 s 492678 163200 492734 164000 6 mprj_dat_o[15]
port 653 nsew signal output
rlabel metal2 s 495346 163200 495402 164000 6 mprj_dat_o[16]
port 654 nsew signal output
rlabel metal2 s 497922 163200 497978 164000 6 mprj_dat_o[17]
port 655 nsew signal output
rlabel metal2 s 500498 163200 500554 164000 6 mprj_dat_o[18]
port 656 nsew signal output
rlabel metal2 s 503074 163200 503130 164000 6 mprj_dat_o[19]
port 657 nsew signal output
rlabel metal2 s 453670 163200 453726 164000 6 mprj_dat_o[1]
port 658 nsew signal output
rlabel metal2 s 505742 163200 505798 164000 6 mprj_dat_o[20]
port 659 nsew signal output
rlabel metal2 s 508318 163200 508374 164000 6 mprj_dat_o[21]
port 660 nsew signal output
rlabel metal2 s 510894 163200 510950 164000 6 mprj_dat_o[22]
port 661 nsew signal output
rlabel metal2 s 513470 163200 513526 164000 6 mprj_dat_o[23]
port 662 nsew signal output
rlabel metal2 s 516138 163200 516194 164000 6 mprj_dat_o[24]
port 663 nsew signal output
rlabel metal2 s 518714 163200 518770 164000 6 mprj_dat_o[25]
port 664 nsew signal output
rlabel metal2 s 521290 163200 521346 164000 6 mprj_dat_o[26]
port 665 nsew signal output
rlabel metal2 s 523866 163200 523922 164000 6 mprj_dat_o[27]
port 666 nsew signal output
rlabel metal2 s 526534 163200 526590 164000 6 mprj_dat_o[28]
port 667 nsew signal output
rlabel metal2 s 529110 163200 529166 164000 6 mprj_dat_o[29]
port 668 nsew signal output
rlabel metal2 s 457166 163200 457222 164000 6 mprj_dat_o[2]
port 669 nsew signal output
rlabel metal2 s 531686 163200 531742 164000 6 mprj_dat_o[30]
port 670 nsew signal output
rlabel metal2 s 534354 163200 534410 164000 6 mprj_dat_o[31]
port 671 nsew signal output
rlabel metal2 s 460662 163200 460718 164000 6 mprj_dat_o[3]
port 672 nsew signal output
rlabel metal2 s 464066 163200 464122 164000 6 mprj_dat_o[4]
port 673 nsew signal output
rlabel metal2 s 466734 163200 466790 164000 6 mprj_dat_o[5]
port 674 nsew signal output
rlabel metal2 s 469310 163200 469366 164000 6 mprj_dat_o[6]
port 675 nsew signal output
rlabel metal2 s 471886 163200 471942 164000 6 mprj_dat_o[7]
port 676 nsew signal output
rlabel metal2 s 474462 163200 474518 164000 6 mprj_dat_o[8]
port 677 nsew signal output
rlabel metal2 s 477130 163200 477186 164000 6 mprj_dat_o[9]
port 678 nsew signal output
rlabel metal2 s 451094 163200 451150 164000 6 mprj_sel_o[0]
port 679 nsew signal output
rlabel metal2 s 454590 163200 454646 164000 6 mprj_sel_o[1]
port 680 nsew signal output
rlabel metal2 s 457994 163200 458050 164000 6 mprj_sel_o[2]
port 681 nsew signal output
rlabel metal2 s 461490 163200 461546 164000 6 mprj_sel_o[3]
port 682 nsew signal output
rlabel metal2 s 445850 163200 445906 164000 6 mprj_stb_o
port 683 nsew signal output
rlabel metal2 s 446770 163200 446826 164000 6 mprj_wb_iena
port 684 nsew signal output
rlabel metal2 s 447598 163200 447654 164000 6 mprj_we_o
port 685 nsew signal output
rlabel metal3 s 539200 90176 540000 90296 6 qspi_enabled
port 686 nsew signal output
rlabel metal3 s 539200 84192 540000 84312 6 ser_rx
port 687 nsew signal input
rlabel metal3 s 539200 85688 540000 85808 6 ser_tx
port 688 nsew signal output
rlabel metal3 s 539200 81064 540000 81184 6 spi_csb
port 689 nsew signal output
rlabel metal3 s 539200 87184 540000 87304 6 spi_enabled
port 690 nsew signal output
rlabel metal3 s 539200 79568 540000 79688 6 spi_sck
port 691 nsew signal output
rlabel metal3 s 539200 82696 540000 82816 6 spi_sdi
port 692 nsew signal input
rlabel metal3 s 539200 78072 540000 78192 6 spi_sdo
port 693 nsew signal output
rlabel metal3 s 539200 76576 540000 76696 6 spi_sdoenb
port 694 nsew signal output
rlabel metal3 s 539200 2184 540000 2304 6 sram_ro_addr[0]
port 695 nsew signal input
rlabel metal3 s 539200 3680 540000 3800 6 sram_ro_addr[1]
port 696 nsew signal input
rlabel metal3 s 539200 5176 540000 5296 6 sram_ro_addr[2]
port 697 nsew signal input
rlabel metal3 s 539200 6672 540000 6792 6 sram_ro_addr[3]
port 698 nsew signal input
rlabel metal3 s 539200 8168 540000 8288 6 sram_ro_addr[4]
port 699 nsew signal input
rlabel metal3 s 539200 9800 540000 9920 6 sram_ro_addr[5]
port 700 nsew signal input
rlabel metal3 s 539200 11296 540000 11416 6 sram_ro_addr[6]
port 701 nsew signal input
rlabel metal3 s 539200 12792 540000 12912 6 sram_ro_addr[7]
port 702 nsew signal input
rlabel metal3 s 539200 14288 540000 14408 6 sram_ro_clk
port 703 nsew signal input
rlabel metal3 s 539200 688 540000 808 6 sram_ro_csb
port 704 nsew signal input
rlabel metal3 s 539200 15784 540000 15904 6 sram_ro_data[0]
port 705 nsew signal output
rlabel metal3 s 539200 31016 540000 31136 6 sram_ro_data[10]
port 706 nsew signal output
rlabel metal3 s 539200 32512 540000 32632 6 sram_ro_data[11]
port 707 nsew signal output
rlabel metal3 s 539200 34008 540000 34128 6 sram_ro_data[12]
port 708 nsew signal output
rlabel metal3 s 539200 35504 540000 35624 6 sram_ro_data[13]
port 709 nsew signal output
rlabel metal3 s 539200 37136 540000 37256 6 sram_ro_data[14]
port 710 nsew signal output
rlabel metal3 s 539200 38632 540000 38752 6 sram_ro_data[15]
port 711 nsew signal output
rlabel metal3 s 539200 40128 540000 40248 6 sram_ro_data[16]
port 712 nsew signal output
rlabel metal3 s 539200 41624 540000 41744 6 sram_ro_data[17]
port 713 nsew signal output
rlabel metal3 s 539200 43120 540000 43240 6 sram_ro_data[18]
port 714 nsew signal output
rlabel metal3 s 539200 44616 540000 44736 6 sram_ro_data[19]
port 715 nsew signal output
rlabel metal3 s 539200 17280 540000 17400 6 sram_ro_data[1]
port 716 nsew signal output
rlabel metal3 s 539200 46248 540000 46368 6 sram_ro_data[20]
port 717 nsew signal output
rlabel metal3 s 539200 47744 540000 47864 6 sram_ro_data[21]
port 718 nsew signal output
rlabel metal3 s 539200 49240 540000 49360 6 sram_ro_data[22]
port 719 nsew signal output
rlabel metal3 s 539200 50736 540000 50856 6 sram_ro_data[23]
port 720 nsew signal output
rlabel metal3 s 539200 52232 540000 52352 6 sram_ro_data[24]
port 721 nsew signal output
rlabel metal3 s 539200 53728 540000 53848 6 sram_ro_data[25]
port 722 nsew signal output
rlabel metal3 s 539200 55360 540000 55480 6 sram_ro_data[26]
port 723 nsew signal output
rlabel metal3 s 539200 56856 540000 56976 6 sram_ro_data[27]
port 724 nsew signal output
rlabel metal3 s 539200 58352 540000 58472 6 sram_ro_data[28]
port 725 nsew signal output
rlabel metal3 s 539200 59848 540000 59968 6 sram_ro_data[29]
port 726 nsew signal output
rlabel metal3 s 539200 18912 540000 19032 6 sram_ro_data[2]
port 727 nsew signal output
rlabel metal3 s 539200 61344 540000 61464 6 sram_ro_data[30]
port 728 nsew signal output
rlabel metal3 s 539200 62840 540000 62960 6 sram_ro_data[31]
port 729 nsew signal output
rlabel metal3 s 539200 20408 540000 20528 6 sram_ro_data[3]
port 730 nsew signal output
rlabel metal3 s 539200 21904 540000 22024 6 sram_ro_data[4]
port 731 nsew signal output
rlabel metal3 s 539200 23400 540000 23520 6 sram_ro_data[5]
port 732 nsew signal output
rlabel metal3 s 539200 24896 540000 25016 6 sram_ro_data[6]
port 733 nsew signal output
rlabel metal3 s 539200 26392 540000 26512 6 sram_ro_data[7]
port 734 nsew signal output
rlabel metal3 s 539200 28024 540000 28144 6 sram_ro_data[8]
port 735 nsew signal output
rlabel metal3 s 539200 29520 540000 29640 6 sram_ro_data[9]
port 736 nsew signal output
rlabel metal3 s 539200 70456 540000 70576 6 trap
port 737 nsew signal output
rlabel metal3 s 539200 88680 540000 88800 6 uart_enabled
port 738 nsew signal output
rlabel metal2 s 535182 163200 535238 164000 6 user_irq_ena[0]
port 739 nsew signal output
rlabel metal2 s 536010 163200 536066 164000 6 user_irq_ena[1]
port 740 nsew signal output
rlabel metal2 s 536930 163200 536986 164000 6 user_irq_ena[2]
port 741 nsew signal output
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 540000 164000
string LEFview TRUE
string GDS_FILE /project/openlane/mgmt_core_wrapper/runs/mgmt_core_wrapper/results/magic/mgmt_core_wrapper.gds
string GDS_END 179937298
string GDS_START 178930976
<< end >>

