magic
tech sky130A
magscale 1 2
timestamp 1640295518
<< metal1 >>
rect 146662 161372 146668 161424
rect 146720 161412 146726 161424
rect 153746 161412 153752 161424
rect 146720 161384 153752 161412
rect 146720 161372 146726 161384
rect 153746 161372 153752 161384
rect 153804 161372 153810 161424
rect 136634 160080 136640 160132
rect 136692 160120 136698 160132
rect 144270 160120 144276 160132
rect 136692 160092 144276 160120
rect 136692 160080 136698 160092
rect 144270 160080 144276 160092
rect 144328 160080 144334 160132
rect 83642 160012 83648 160064
rect 83700 160052 83706 160064
rect 166994 160052 167000 160064
rect 83700 160024 167000 160052
rect 83700 160012 83706 160024
rect 166994 160012 167000 160024
rect 167052 160012 167058 160064
rect 170214 160012 170220 160064
rect 170272 160052 170278 160064
rect 198918 160052 198924 160064
rect 170272 160024 198924 160052
rect 170272 160012 170278 160024
rect 198918 160012 198924 160024
rect 198976 160012 198982 160064
rect 203058 160012 203064 160064
rect 203116 160052 203122 160064
rect 211062 160052 211068 160064
rect 203116 160024 211068 160052
rect 203116 160012 203122 160024
rect 211062 160012 211068 160024
rect 211120 160012 211126 160064
rect 211430 160012 211436 160064
rect 211488 160052 211494 160064
rect 280338 160052 280344 160064
rect 211488 160024 280344 160052
rect 211488 160012 211494 160024
rect 280338 160012 280344 160024
rect 280396 160012 280402 160064
rect 281258 160012 281264 160064
rect 281316 160052 281322 160064
rect 332686 160052 332692 160064
rect 281316 160024 332692 160052
rect 281316 160012 281322 160024
rect 332686 160012 332692 160024
rect 332744 160012 332750 160064
rect 335078 160012 335084 160064
rect 335136 160052 335142 160064
rect 373994 160052 374000 160064
rect 335136 160024 374000 160052
rect 335136 160012 335142 160024
rect 373994 160012 374000 160024
rect 374052 160012 374058 160064
rect 378870 160012 378876 160064
rect 378928 160052 378934 160064
rect 398558 160052 398564 160064
rect 378928 160024 398564 160052
rect 378928 160012 378934 160024
rect 398558 160012 398564 160024
rect 398616 160012 398622 160064
rect 25590 159944 25596 159996
rect 25648 159984 25654 159996
rect 109862 159984 109868 159996
rect 25648 159956 109868 159984
rect 25648 159944 25654 159956
rect 109862 159944 109868 159956
rect 109920 159944 109926 159996
rect 117222 159944 117228 159996
rect 117280 159984 117286 159996
rect 191742 159984 191748 159996
rect 117280 159956 191748 159984
rect 117280 159944 117286 159956
rect 191742 159944 191748 159956
rect 191800 159944 191806 159996
rect 197998 159944 198004 159996
rect 198056 159984 198062 159996
rect 269114 159984 269120 159996
rect 198056 159956 269120 159984
rect 198056 159944 198062 159956
rect 269114 159944 269120 159956
rect 269172 159944 269178 159996
rect 271230 159944 271236 159996
rect 271288 159984 271294 159996
rect 272794 159984 272800 159996
rect 271288 159956 272800 159984
rect 271288 159944 271294 159956
rect 272794 159944 272800 159956
rect 272852 159944 272858 159996
rect 275370 159944 275376 159996
rect 275428 159984 275434 159996
rect 329098 159984 329104 159996
rect 275428 159956 329104 159984
rect 275428 159944 275434 159956
rect 329098 159944 329104 159956
rect 329156 159944 329162 159996
rect 329190 159944 329196 159996
rect 329248 159984 329254 159996
rect 369854 159984 369860 159996
rect 329248 159956 369860 159984
rect 329248 159944 329254 159956
rect 369854 159944 369860 159956
rect 369912 159944 369918 159996
rect 372154 159944 372160 159996
rect 372212 159984 372218 159996
rect 396166 159984 396172 159996
rect 372212 159956 396172 159984
rect 372212 159944 372218 159956
rect 396166 159944 396172 159956
rect 396224 159944 396230 159996
rect 399018 159944 399024 159996
rect 399076 159984 399082 159996
rect 408494 159984 408500 159996
rect 399076 159956 408500 159984
rect 399076 159944 399082 159956
rect 408494 159944 408500 159956
rect 408552 159944 408558 159996
rect 476114 159984 476120 159996
rect 470566 159956 476120 159984
rect 470566 159928 470594 159956
rect 476114 159944 476120 159956
rect 476172 159944 476178 159996
rect 70118 159876 70124 159928
rect 70176 159916 70182 159928
rect 148686 159916 148692 159928
rect 70176 159888 148692 159916
rect 70176 159876 70182 159888
rect 148686 159876 148692 159888
rect 148744 159876 148750 159928
rect 152458 159876 152464 159928
rect 152516 159916 152522 159928
rect 160094 159916 160100 159928
rect 152516 159888 160100 159916
rect 152516 159876 152522 159888
rect 160094 159876 160100 159888
rect 160152 159876 160158 159928
rect 160186 159876 160192 159928
rect 160244 159916 160250 159928
rect 188246 159916 188252 159928
rect 160244 159888 188252 159916
rect 160244 159876 160250 159888
rect 188246 159876 188252 159888
rect 188304 159876 188310 159928
rect 191282 159876 191288 159928
rect 191340 159916 191346 159928
rect 264882 159916 264888 159928
rect 191340 159888 264888 159916
rect 191340 159876 191346 159888
rect 264882 159876 264888 159888
rect 264940 159876 264946 159928
rect 268654 159876 268660 159928
rect 268712 159916 268718 159928
rect 324038 159916 324044 159928
rect 268712 159888 324044 159916
rect 268712 159876 268718 159888
rect 324038 159876 324044 159888
rect 324096 159876 324102 159928
rect 328362 159876 328368 159928
rect 328420 159916 328426 159928
rect 369486 159916 369492 159928
rect 328420 159888 369492 159916
rect 328420 159876 328426 159888
rect 369486 159876 369492 159888
rect 369544 159876 369550 159928
rect 379698 159876 379704 159928
rect 379756 159916 379762 159928
rect 405826 159916 405832 159928
rect 379756 159888 405832 159916
rect 379756 159876 379762 159888
rect 405826 159876 405832 159888
rect 405884 159876 405890 159928
rect 470502 159876 470508 159928
rect 470560 159888 470594 159928
rect 470560 159876 470566 159888
rect 471422 159876 471428 159928
rect 471480 159916 471486 159928
rect 477678 159916 477684 159928
rect 471480 159888 477684 159916
rect 471480 159876 471486 159888
rect 477678 159876 477684 159888
rect 477736 159876 477742 159928
rect 480622 159876 480628 159928
rect 480680 159916 480686 159928
rect 485958 159916 485964 159928
rect 480680 159888 485964 159916
rect 480680 159876 480686 159888
rect 485958 159876 485964 159888
rect 486016 159876 486022 159928
rect 56686 159808 56692 159860
rect 56744 159848 56750 159860
rect 136542 159848 136548 159860
rect 56744 159820 136548 159848
rect 56744 159808 56750 159820
rect 136542 159808 136548 159820
rect 136600 159808 136606 159860
rect 142614 159808 142620 159860
rect 142672 159848 142678 159860
rect 146294 159848 146300 159860
rect 142672 159820 146300 159848
rect 142672 159808 142678 159820
rect 146294 159808 146300 159820
rect 146352 159808 146358 159860
rect 153746 159808 153752 159860
rect 153804 159848 153810 159860
rect 174998 159848 175004 159860
rect 153804 159820 175004 159848
rect 153804 159808 153810 159820
rect 174998 159808 175004 159820
rect 175056 159808 175062 159860
rect 180702 159848 180708 159860
rect 175936 159820 180708 159848
rect 63402 159740 63408 159792
rect 63460 159780 63466 159792
rect 146846 159780 146852 159792
rect 63460 159752 139900 159780
rect 63460 159740 63466 159752
rect 18874 159672 18880 159724
rect 18932 159712 18938 159724
rect 107286 159712 107292 159724
rect 18932 159684 107292 159712
rect 18932 159672 18938 159684
rect 107286 159672 107292 159684
rect 107344 159672 107350 159724
rect 109678 159672 109684 159724
rect 109736 159712 109742 159724
rect 137646 159712 137652 159724
rect 109736 159684 137652 159712
rect 109736 159672 109742 159684
rect 137646 159672 137652 159684
rect 137704 159672 137710 159724
rect 139872 159712 139900 159752
rect 140056 159752 146852 159780
rect 140056 159712 140084 159752
rect 146846 159740 146852 159752
rect 146904 159740 146910 159792
rect 148594 159740 148600 159792
rect 148652 159780 148658 159792
rect 148652 159752 149100 159780
rect 148652 159740 148658 159752
rect 139872 159684 140084 159712
rect 144270 159672 144276 159724
rect 144328 159712 144334 159724
rect 148778 159712 148784 159724
rect 144328 159684 148784 159712
rect 144328 159672 144334 159684
rect 148778 159672 148784 159684
rect 148836 159672 148842 159724
rect 148962 159672 148968 159724
rect 149020 159672 149026 159724
rect 149072 159712 149100 159752
rect 150802 159740 150808 159792
rect 150860 159780 150866 159792
rect 152550 159780 152556 159792
rect 150860 159752 152556 159780
rect 150860 159740 150866 159752
rect 152550 159740 152556 159752
rect 152608 159740 152614 159792
rect 153470 159740 153476 159792
rect 153528 159780 153534 159792
rect 175936 159780 175964 159820
rect 180702 159808 180708 159820
rect 180760 159808 180766 159860
rect 184566 159808 184572 159860
rect 184624 159848 184630 159860
rect 259546 159848 259552 159860
rect 184624 159820 259552 159848
rect 184624 159808 184630 159820
rect 259546 159808 259552 159820
rect 259604 159808 259610 159860
rect 261938 159808 261944 159860
rect 261996 159848 262002 159860
rect 318794 159848 318800 159860
rect 261996 159820 318800 159848
rect 261996 159808 262002 159820
rect 318794 159808 318800 159820
rect 318852 159808 318858 159860
rect 320818 159808 320824 159860
rect 320876 159848 320882 159860
rect 362954 159848 362960 159860
rect 320876 159820 362960 159848
rect 320876 159808 320882 159820
rect 362954 159808 362960 159820
rect 363012 159808 363018 159860
rect 376294 159808 376300 159860
rect 376352 159848 376358 159860
rect 406194 159848 406200 159860
rect 376352 159820 406200 159848
rect 376352 159808 376358 159820
rect 406194 159808 406200 159820
rect 406252 159808 406258 159860
rect 409966 159808 409972 159860
rect 410024 159848 410030 159860
rect 417418 159848 417424 159860
rect 410024 159820 417424 159848
rect 410024 159808 410030 159820
rect 417418 159808 417424 159820
rect 417476 159808 417482 159860
rect 467190 159808 467196 159860
rect 467248 159848 467254 159860
rect 473354 159848 473360 159860
rect 467248 159820 473360 159848
rect 467248 159808 467254 159820
rect 473354 159808 473360 159820
rect 473412 159808 473418 159860
rect 153528 159752 175964 159780
rect 153528 159740 153534 159752
rect 177850 159740 177856 159792
rect 177908 159780 177914 159792
rect 253934 159780 253940 159792
rect 177908 159752 253940 159780
rect 177908 159740 177914 159752
rect 253934 159740 253940 159752
rect 253992 159740 253998 159792
rect 255222 159740 255228 159792
rect 255280 159780 255286 159792
rect 313366 159780 313372 159792
rect 255280 159752 313372 159780
rect 255280 159740 255286 159752
rect 313366 159740 313372 159752
rect 313424 159740 313430 159792
rect 314102 159740 314108 159792
rect 314160 159780 314166 159792
rect 357986 159780 357992 159792
rect 314160 159752 357992 159780
rect 314160 159740 314166 159752
rect 357986 159740 357992 159752
rect 358044 159740 358050 159792
rect 365438 159740 365444 159792
rect 365496 159780 365502 159792
rect 395522 159780 395528 159792
rect 365496 159752 395528 159780
rect 365496 159740 365502 159752
rect 395522 159740 395528 159752
rect 395580 159740 395586 159792
rect 396534 159740 396540 159792
rect 396592 159780 396598 159792
rect 413186 159780 413192 159792
rect 396592 159752 413192 159780
rect 396592 159740 396598 159752
rect 413186 159740 413192 159752
rect 413244 159740 413250 159792
rect 424318 159740 424324 159792
rect 424376 159780 424382 159792
rect 442810 159780 442816 159792
rect 424376 159752 442816 159780
rect 424376 159740 424382 159752
rect 442810 159740 442816 159752
rect 442868 159740 442874 159792
rect 472250 159740 472256 159792
rect 472308 159780 472314 159792
rect 479426 159780 479432 159792
rect 472308 159752 479432 159780
rect 472308 159740 472314 159752
rect 479426 159740 479432 159752
rect 479484 159740 479490 159792
rect 479794 159740 479800 159792
rect 479852 159780 479858 159792
rect 485222 159780 485228 159792
rect 479852 159752 485228 159780
rect 479852 159740 479858 159752
rect 485222 159740 485228 159752
rect 485280 159740 485286 159792
rect 164142 159712 164148 159724
rect 149072 159684 164148 159712
rect 164142 159672 164148 159684
rect 164200 159672 164206 159724
rect 167730 159672 167736 159724
rect 167788 159712 167794 159724
rect 246942 159712 246948 159724
rect 167788 159684 246948 159712
rect 167788 159672 167794 159684
rect 246942 159672 246948 159684
rect 247000 159672 247006 159724
rect 248506 159672 248512 159724
rect 248564 159712 248570 159724
rect 301406 159712 301412 159724
rect 248564 159684 301412 159712
rect 248564 159672 248570 159684
rect 301406 159672 301412 159684
rect 301464 159672 301470 159724
rect 303522 159712 303528 159724
rect 301516 159684 303528 159712
rect 49970 159604 49976 159656
rect 50028 159644 50034 159656
rect 142246 159644 142252 159656
rect 50028 159616 142252 159644
rect 50028 159604 50034 159616
rect 142246 159604 142252 159616
rect 142304 159604 142310 159656
rect 143350 159604 143356 159656
rect 143408 159644 143414 159656
rect 148594 159644 148600 159656
rect 143408 159616 148600 159644
rect 143408 159604 143414 159616
rect 148594 159604 148600 159616
rect 148652 159604 148658 159656
rect 148980 159644 149008 159672
rect 160094 159644 160100 159656
rect 148980 159616 160100 159644
rect 160094 159604 160100 159616
rect 160152 159604 160158 159656
rect 161014 159604 161020 159656
rect 161072 159644 161078 159656
rect 240318 159644 240324 159656
rect 161072 159616 240324 159644
rect 161072 159604 161078 159616
rect 240318 159604 240324 159616
rect 240376 159604 240382 159656
rect 241790 159604 241796 159656
rect 241848 159644 241854 159656
rect 301516 159644 301544 159684
rect 303522 159672 303528 159684
rect 303580 159672 303586 159724
rect 309042 159672 309048 159724
rect 309100 159712 309106 159724
rect 354858 159712 354864 159724
rect 309100 159684 354864 159712
rect 309100 159672 309106 159684
rect 354858 159672 354864 159684
rect 354916 159672 354922 159724
rect 357802 159672 357808 159724
rect 357860 159712 357866 159724
rect 369210 159712 369216 159724
rect 357860 159684 369216 159712
rect 357860 159672 357866 159684
rect 369210 159672 369216 159684
rect 369268 159672 369274 159724
rect 369578 159672 369584 159724
rect 369636 159712 369642 159724
rect 401042 159712 401048 159724
rect 369636 159684 401048 159712
rect 369636 159672 369642 159684
rect 401042 159672 401048 159684
rect 401100 159672 401106 159724
rect 403250 159672 403256 159724
rect 403308 159712 403314 159724
rect 416590 159712 416596 159724
rect 403308 159684 416596 159712
rect 403308 159672 403314 159684
rect 416590 159672 416596 159684
rect 416648 159672 416654 159724
rect 420914 159672 420920 159724
rect 420972 159712 420978 159724
rect 440418 159712 440424 159724
rect 420972 159684 440424 159712
rect 420972 159672 420978 159684
rect 440418 159672 440424 159684
rect 440476 159672 440482 159724
rect 241848 159616 301544 159644
rect 241848 159604 241854 159616
rect 302326 159604 302332 159656
rect 302384 159644 302390 159656
rect 349246 159644 349252 159656
rect 302384 159616 349252 159644
rect 302384 159604 302390 159616
rect 349246 159604 349252 159616
rect 349304 159604 349310 159656
rect 351914 159604 351920 159656
rect 351972 159644 351978 159656
rect 385310 159644 385316 159656
rect 351972 159616 385316 159644
rect 351972 159604 351978 159616
rect 385310 159604 385316 159616
rect 385368 159604 385374 159656
rect 389818 159604 389824 159656
rect 389876 159644 389882 159656
rect 413830 159644 413836 159656
rect 389876 159616 413836 159644
rect 389876 159604 389882 159616
rect 413830 159604 413836 159616
rect 413888 159604 413894 159656
rect 417510 159604 417516 159656
rect 417568 159644 417574 159656
rect 437658 159644 437664 159656
rect 417568 159616 437664 159644
rect 417568 159604 417574 159616
rect 437658 159604 437664 159616
rect 437716 159604 437722 159656
rect 448698 159604 448704 159656
rect 448756 159644 448762 159656
rect 455874 159644 455880 159656
rect 448756 159616 455880 159644
rect 448756 159604 448762 159616
rect 455874 159604 455880 159616
rect 455932 159604 455938 159656
rect 32306 159536 32312 159588
rect 32364 159576 32370 159588
rect 126238 159576 126244 159588
rect 32364 159548 126244 159576
rect 32364 159536 32370 159548
rect 126238 159536 126244 159548
rect 126296 159536 126302 159588
rect 127618 159536 127624 159588
rect 127676 159576 127682 159588
rect 139854 159576 139860 159588
rect 127676 159548 139860 159576
rect 127676 159536 127682 159548
rect 139854 159536 139860 159548
rect 139912 159536 139918 159588
rect 139946 159536 139952 159588
rect 140004 159576 140010 159588
rect 157242 159576 157248 159588
rect 140004 159548 157248 159576
rect 140004 159536 140010 159548
rect 157242 159536 157248 159548
rect 157300 159536 157306 159588
rect 157610 159536 157616 159588
rect 157668 159576 157674 159588
rect 239306 159576 239312 159588
rect 157668 159548 239312 159576
rect 157668 159536 157674 159548
rect 239306 159536 239312 159548
rect 239364 159536 239370 159588
rect 250990 159536 250996 159588
rect 251048 159576 251054 159588
rect 310606 159576 310612 159588
rect 251048 159548 310612 159576
rect 251048 159536 251054 159548
rect 310606 159536 310612 159548
rect 310664 159536 310670 159588
rect 315758 159536 315764 159588
rect 315816 159576 315822 159588
rect 358906 159576 358912 159588
rect 315816 159548 358912 159576
rect 315816 159536 315822 159548
rect 358906 159536 358912 159548
rect 358964 159536 358970 159588
rect 362862 159536 362868 159588
rect 362920 159576 362926 159588
rect 395982 159576 395988 159588
rect 362920 159548 395988 159576
rect 362920 159536 362926 159548
rect 395982 159536 395988 159548
rect 396040 159536 396046 159588
rect 407482 159536 407488 159588
rect 407540 159576 407546 159588
rect 429930 159576 429936 159588
rect 407540 159548 429936 159576
rect 407540 159536 407546 159548
rect 429930 159536 429936 159548
rect 429988 159536 429994 159588
rect 450354 159536 450360 159588
rect 450412 159576 450418 159588
rect 457162 159576 457168 159588
rect 450412 159548 457168 159576
rect 450412 159536 450418 159548
rect 457162 159536 457168 159548
rect 457220 159536 457226 159588
rect 458726 159536 458732 159588
rect 458784 159576 458790 159588
rect 465074 159576 465080 159588
rect 458784 159548 465080 159576
rect 458784 159536 458790 159548
rect 465074 159536 465080 159548
rect 465132 159536 465138 159588
rect 468018 159536 468024 159588
rect 468076 159576 468082 159588
rect 476022 159576 476028 159588
rect 468076 159548 476028 159576
rect 468076 159536 468082 159548
rect 476022 159536 476028 159548
rect 476080 159536 476086 159588
rect 478966 159536 478972 159588
rect 479024 159576 479030 159588
rect 484578 159576 484584 159588
rect 479024 159548 484584 159576
rect 479024 159536 479030 159548
rect 484578 159536 484584 159548
rect 484636 159536 484642 159588
rect 43254 159468 43260 159520
rect 43312 159508 43318 159520
rect 43312 159480 136496 159508
rect 43312 159468 43318 159480
rect 36538 159400 36544 159452
rect 36596 159440 36602 159452
rect 135162 159440 135168 159452
rect 36596 159412 135168 159440
rect 36596 159400 36602 159412
rect 135162 159400 135168 159412
rect 135220 159400 135226 159452
rect 136468 159440 136496 159480
rect 136542 159468 136548 159520
rect 136600 159508 136606 159520
rect 136600 159480 142936 159508
rect 136600 159468 136606 159480
rect 137370 159440 137376 159452
rect 136468 159412 137376 159440
rect 137370 159400 137376 159412
rect 137428 159400 137434 159452
rect 137462 159400 137468 159452
rect 137520 159440 137526 159452
rect 142908 159440 142936 159480
rect 144178 159468 144184 159520
rect 144236 159508 144242 159520
rect 225230 159508 225236 159520
rect 144236 159480 225236 159508
rect 144236 159468 144242 159480
rect 225230 159468 225236 159480
rect 225288 159468 225294 159520
rect 231670 159468 231676 159520
rect 231728 159508 231734 159520
rect 295518 159508 295524 159520
rect 231728 159480 295524 159508
rect 231728 159468 231734 159480
rect 295518 159468 295524 159480
rect 295576 159468 295582 159520
rect 295610 159468 295616 159520
rect 295668 159508 295674 159520
rect 342438 159508 342444 159520
rect 295668 159480 342444 159508
rect 295668 159468 295674 159480
rect 342438 159468 342444 159480
rect 342496 159468 342502 159520
rect 347682 159468 347688 159520
rect 347740 159508 347746 159520
rect 354214 159508 354220 159520
rect 347740 159480 354220 159508
rect 347740 159468 347746 159480
rect 354214 159468 354220 159480
rect 354272 159468 354278 159520
rect 356146 159468 356152 159520
rect 356204 159508 356210 159520
rect 390554 159508 390560 159520
rect 356204 159480 390560 159508
rect 356204 159468 356210 159480
rect 390554 159468 390560 159480
rect 390612 159468 390618 159520
rect 392302 159468 392308 159520
rect 392360 159508 392366 159520
rect 404262 159508 404268 159520
rect 392360 159480 404268 159508
rect 392360 159468 392366 159480
rect 404262 159468 404268 159480
rect 404320 159468 404326 159520
rect 410794 159468 410800 159520
rect 410852 159508 410858 159520
rect 432506 159508 432512 159520
rect 410852 159480 432512 159508
rect 410852 159468 410858 159480
rect 432506 159468 432512 159480
rect 432564 159468 432570 159520
rect 449526 159468 449532 159520
rect 449584 159508 449590 159520
rect 455506 159508 455512 159520
rect 449584 159480 455512 159508
rect 449584 159468 449590 159480
rect 455506 159468 455512 159480
rect 455564 159468 455570 159520
rect 457070 159468 457076 159520
rect 457128 159508 457134 159520
rect 464338 159508 464344 159520
rect 457128 159480 464344 159508
rect 457128 159468 457134 159480
rect 464338 159468 464344 159480
rect 464396 159468 464402 159520
rect 144822 159440 144828 159452
rect 137520 159412 142844 159440
rect 142908 159412 144828 159440
rect 137520 159400 137526 159412
rect 6270 159332 6276 159384
rect 6328 159372 6334 159384
rect 122834 159372 122840 159384
rect 6328 159344 122840 159372
rect 6328 159332 6334 159344
rect 122834 159332 122840 159344
rect 122892 159332 122898 159384
rect 123110 159332 123116 159384
rect 123168 159372 123174 159384
rect 142614 159372 142620 159384
rect 123168 159344 142620 159372
rect 123168 159332 123174 159344
rect 142614 159332 142620 159344
rect 142672 159332 142678 159384
rect 142816 159372 142844 159412
rect 144822 159400 144828 159412
rect 144880 159400 144886 159452
rect 144914 159400 144920 159452
rect 144972 159440 144978 159452
rect 146202 159440 146208 159452
rect 144972 159412 146208 159440
rect 144972 159400 144978 159412
rect 146202 159400 146208 159412
rect 146260 159400 146266 159452
rect 146294 159400 146300 159452
rect 146352 159440 146358 159452
rect 147122 159440 147128 159452
rect 146352 159412 147128 159440
rect 146352 159400 146358 159412
rect 147122 159400 147128 159412
rect 147180 159400 147186 159452
rect 147582 159400 147588 159452
rect 147640 159440 147646 159452
rect 149054 159440 149060 159452
rect 147640 159412 149060 159440
rect 147640 159400 147646 159412
rect 149054 159400 149060 159412
rect 149112 159400 149118 159452
rect 149146 159400 149152 159452
rect 149204 159440 149210 159452
rect 150802 159440 150808 159452
rect 149204 159412 150808 159440
rect 149204 159400 149210 159412
rect 150802 159400 150808 159412
rect 150860 159400 150866 159452
rect 150894 159400 150900 159452
rect 150952 159440 150958 159452
rect 234062 159440 234068 159452
rect 150952 159412 234068 159440
rect 150952 159400 150958 159412
rect 234062 159400 234068 159412
rect 234120 159400 234126 159452
rect 234982 159400 234988 159452
rect 235040 159440 235046 159452
rect 298002 159440 298008 159452
rect 235040 159412 298008 159440
rect 235040 159400 235046 159412
rect 298002 159400 298008 159412
rect 298060 159400 298066 159452
rect 301498 159400 301504 159452
rect 301556 159440 301562 159452
rect 349062 159440 349068 159452
rect 301556 159412 349068 159440
rect 301556 159400 301562 159412
rect 349062 159400 349068 159412
rect 349120 159400 349126 159452
rect 349338 159400 349344 159452
rect 349396 159440 349402 159452
rect 353202 159440 353208 159452
rect 349396 159412 353208 159440
rect 349396 159400 349402 159412
rect 353202 159400 353208 159412
rect 353260 159400 353266 159452
rect 358630 159400 358636 159452
rect 358688 159440 358694 159452
rect 392762 159440 392768 159452
rect 358688 159412 392768 159440
rect 358688 159400 358694 159412
rect 392762 159400 392768 159412
rect 392820 159400 392826 159452
rect 404078 159400 404084 159452
rect 404136 159440 404142 159452
rect 427354 159440 427360 159452
rect 404136 159412 427360 159440
rect 404136 159400 404142 159412
rect 427354 159400 427360 159412
rect 427412 159400 427418 159452
rect 427630 159400 427636 159452
rect 427688 159440 427694 159452
rect 445386 159440 445392 159452
rect 427688 159412 445392 159440
rect 427688 159400 427694 159412
rect 445386 159400 445392 159412
rect 445444 159400 445450 159452
rect 451182 159400 451188 159452
rect 451240 159440 451246 159452
rect 456794 159440 456800 159452
rect 451240 159412 456800 159440
rect 451240 159400 451246 159412
rect 456794 159400 456800 159412
rect 456852 159400 456858 159452
rect 459646 159400 459652 159452
rect 459704 159440 459710 159452
rect 466454 159440 466460 159452
rect 459704 159412 466460 159440
rect 459704 159400 459710 159412
rect 466454 159400 466460 159412
rect 466512 159400 466518 159452
rect 468846 159400 468852 159452
rect 468904 159440 468910 159452
rect 474826 159440 474832 159452
rect 468904 159412 474832 159440
rect 468904 159400 468910 159412
rect 474826 159400 474832 159412
rect 474884 159400 474890 159452
rect 477310 159400 477316 159452
rect 477368 159440 477374 159452
rect 483290 159440 483296 159452
rect 477368 159412 483296 159440
rect 477368 159400 477374 159412
rect 483290 159400 483296 159412
rect 483348 159400 483354 159452
rect 518802 159400 518808 159452
rect 518860 159440 518866 159452
rect 522666 159440 522672 159452
rect 518860 159412 522672 159440
rect 518860 159400 518866 159412
rect 522666 159400 522672 159412
rect 522724 159400 522730 159452
rect 223666 159372 223672 159384
rect 142816 159344 223672 159372
rect 223666 159332 223672 159344
rect 223724 159332 223730 159384
rect 224954 159332 224960 159384
rect 225012 159372 225018 159384
rect 290642 159372 290648 159384
rect 225012 159344 290648 159372
rect 225012 159332 225018 159344
rect 290642 159332 290648 159344
rect 290700 159332 290706 159384
rect 294782 159332 294788 159384
rect 294840 159372 294846 159384
rect 342254 159372 342260 159384
rect 294840 159344 342260 159372
rect 294840 159332 294846 159344
rect 342254 159332 342260 159344
rect 342312 159332 342318 159384
rect 342714 159332 342720 159384
rect 342772 159372 342778 159384
rect 343634 159372 343640 159384
rect 342772 159344 343640 159372
rect 342772 159332 342778 159344
rect 343634 159332 343640 159344
rect 343692 159332 343698 159384
rect 346026 159332 346032 159384
rect 346084 159372 346090 159384
rect 382826 159372 382832 159384
rect 346084 159344 382832 159372
rect 346084 159332 346090 159344
rect 382826 159332 382832 159344
rect 382884 159332 382890 159384
rect 383102 159332 383108 159384
rect 383160 159372 383166 159384
rect 411346 159372 411352 159384
rect 383160 159344 411352 159372
rect 383160 159332 383166 159344
rect 411346 159332 411352 159344
rect 411404 159332 411410 159384
rect 414198 159332 414204 159384
rect 414256 159372 414262 159384
rect 435082 159372 435088 159384
rect 414256 159344 435088 159372
rect 414256 159332 414262 159344
rect 435082 159332 435088 159344
rect 435140 159332 435146 159384
rect 447870 159332 447876 159384
rect 447928 159372 447934 159384
rect 456886 159372 456892 159384
rect 447928 159344 456892 159372
rect 447928 159332 447934 159344
rect 456886 159332 456892 159344
rect 456944 159332 456950 159384
rect 469674 159332 469680 159384
rect 469732 159372 469738 159384
rect 477402 159372 477408 159384
rect 469732 159344 477408 159372
rect 469732 159332 469738 159344
rect 477402 159332 477408 159344
rect 477460 159332 477466 159384
rect 478138 159332 478144 159384
rect 478196 159372 478202 159384
rect 483198 159372 483204 159384
rect 478196 159344 483204 159372
rect 478196 159332 478202 159344
rect 483198 159332 483204 159344
rect 483256 159332 483262 159384
rect 518710 159332 518716 159384
rect 518768 159372 518774 159384
rect 523494 159372 523500 159384
rect 518768 159344 523500 159372
rect 518768 159332 518774 159344
rect 523494 159332 523500 159344
rect 523552 159332 523558 159384
rect 76926 159264 76932 159316
rect 76984 159304 76990 159316
rect 152458 159304 152464 159316
rect 76984 159276 152464 159304
rect 76984 159264 76990 159276
rect 152458 159264 152464 159276
rect 152516 159264 152522 159316
rect 152550 159264 152556 159316
rect 152608 159304 152614 159316
rect 156046 159304 156052 159316
rect 152608 159276 156052 159304
rect 152608 159264 152614 159276
rect 156046 159264 156052 159276
rect 156104 159264 156110 159316
rect 163498 159264 163504 159316
rect 163556 159304 163562 159316
rect 193582 159304 193588 159316
rect 163556 159276 193588 159304
rect 163556 159264 163562 159276
rect 193582 159264 193588 159276
rect 193640 159264 193646 159316
rect 193674 159264 193680 159316
rect 193732 159304 193738 159316
rect 197354 159304 197360 159316
rect 193732 159276 197360 159304
rect 193732 159264 193738 159276
rect 197354 159264 197360 159276
rect 197412 159264 197418 159316
rect 201402 159264 201408 159316
rect 201460 159304 201466 159316
rect 207382 159304 207388 159316
rect 201460 159276 207388 159304
rect 201460 159264 201466 159276
rect 207382 159264 207388 159276
rect 207440 159264 207446 159316
rect 208118 159264 208124 159316
rect 208176 159304 208182 159316
rect 212442 159304 212448 159316
rect 208176 159276 212448 159304
rect 208176 159264 208182 159276
rect 212442 159264 212448 159276
rect 212500 159264 212506 159316
rect 214006 159264 214012 159316
rect 214064 159304 214070 159316
rect 281534 159304 281540 159316
rect 214064 159276 281540 159304
rect 214064 159264 214070 159276
rect 281534 159264 281540 159276
rect 281592 159264 281598 159316
rect 282086 159264 282092 159316
rect 282144 159304 282150 159316
rect 334158 159304 334164 159316
rect 282144 159276 334164 159304
rect 282144 159264 282150 159276
rect 334158 159264 334164 159276
rect 334216 159264 334222 159316
rect 334250 159264 334256 159316
rect 334308 159304 334314 159316
rect 374086 159304 374092 159316
rect 334308 159276 374092 159304
rect 334308 159264 334314 159276
rect 374086 159264 374092 159276
rect 374144 159264 374150 159316
rect 378042 159264 378048 159316
rect 378100 159304 378106 159316
rect 388346 159304 388352 159316
rect 378100 159276 388352 159304
rect 378100 159264 378106 159276
rect 388346 159264 388352 159276
rect 388404 159264 388410 159316
rect 395706 159264 395712 159316
rect 395764 159304 395770 159316
rect 404722 159304 404728 159316
rect 395764 159276 404728 159304
rect 395764 159264 395770 159276
rect 404722 159264 404728 159276
rect 404780 159264 404786 159316
rect 460474 159264 460480 159316
rect 460532 159304 460538 159316
rect 466638 159304 466644 159316
rect 460532 159276 466644 159304
rect 460532 159264 460538 159276
rect 466638 159264 466644 159276
rect 466696 159264 466702 159316
rect 93670 159196 93676 159248
rect 93728 159236 93734 159248
rect 175826 159236 175832 159248
rect 93728 159208 175832 159236
rect 93728 159196 93734 159208
rect 175826 159196 175832 159208
rect 175884 159196 175890 159248
rect 183094 159236 183100 159248
rect 176028 159208 183100 159236
rect 86954 159128 86960 159180
rect 87012 159168 87018 159180
rect 169754 159168 169760 159180
rect 87012 159140 169760 159168
rect 87012 159128 87018 159140
rect 169754 159128 169760 159140
rect 169812 159128 169818 159180
rect 173618 159128 173624 159180
rect 173676 159168 173682 159180
rect 175918 159168 175924 159180
rect 173676 159140 175924 159168
rect 173676 159128 173682 159140
rect 175918 159128 175924 159140
rect 175976 159128 175982 159180
rect 100478 159060 100484 159112
rect 100536 159100 100542 159112
rect 176028 159100 176056 159208
rect 183094 159196 183100 159208
rect 183152 159196 183158 159248
rect 187050 159196 187056 159248
rect 187108 159236 187114 159248
rect 216766 159236 216772 159248
rect 187108 159208 216772 159236
rect 187108 159196 187114 159208
rect 216766 159196 216772 159208
rect 216824 159196 216830 159248
rect 218238 159196 218244 159248
rect 218296 159236 218302 159248
rect 284386 159236 284392 159248
rect 218296 159208 284392 159236
rect 218296 159196 218302 159208
rect 284386 159196 284392 159208
rect 284444 159196 284450 159248
rect 287974 159196 287980 159248
rect 288032 159236 288038 159248
rect 338758 159236 338764 159248
rect 288032 159208 338764 159236
rect 288032 159196 288038 159208
rect 338758 159196 338764 159208
rect 338816 159196 338822 159248
rect 339310 159196 339316 159248
rect 339368 159236 339374 159248
rect 377950 159236 377956 159248
rect 339368 159208 377956 159236
rect 339368 159196 339374 159208
rect 377950 159196 377956 159208
rect 378008 159196 378014 159248
rect 385586 159196 385592 159248
rect 385644 159236 385650 159248
rect 398834 159236 398840 159248
rect 385644 159208 398840 159236
rect 385644 159196 385650 159208
rect 398834 159196 398840 159208
rect 398892 159196 398898 159248
rect 453758 159196 453764 159248
rect 453816 159236 453822 159248
rect 459554 159236 459560 159248
rect 453816 159208 459560 159236
rect 453816 159196 453822 159208
rect 459554 159196 459560 159208
rect 459612 159196 459618 159248
rect 462958 159196 462964 159248
rect 463016 159236 463022 159248
rect 469214 159236 469220 159248
rect 463016 159208 469220 159236
rect 463016 159196 463022 159208
rect 469214 159196 469220 159208
rect 469272 159196 469278 159248
rect 176102 159128 176108 159180
rect 176160 159168 176166 159180
rect 193674 159168 193680 159180
rect 176160 159140 193680 159168
rect 176160 159128 176166 159140
rect 193674 159128 193680 159140
rect 193732 159128 193738 159180
rect 193766 159128 193772 159180
rect 193824 159168 193830 159180
rect 193824 159140 200114 159168
rect 193824 159128 193830 159140
rect 100536 159072 176056 159100
rect 100536 159060 100542 159072
rect 180334 159060 180340 159112
rect 180392 159100 180398 159112
rect 200086 159100 200114 159140
rect 203886 159128 203892 159180
rect 203944 159168 203950 159180
rect 206922 159168 206928 159180
rect 203944 159140 206928 159168
rect 203944 159128 203950 159140
rect 206922 159128 206928 159140
rect 206980 159128 206986 159180
rect 220630 159168 220636 159180
rect 207032 159140 220636 159168
rect 207032 159100 207060 159140
rect 220630 159128 220636 159140
rect 220688 159128 220694 159180
rect 220722 159128 220728 159180
rect 220780 159168 220786 159180
rect 283190 159168 283196 159180
rect 220780 159140 283196 159168
rect 220780 159128 220786 159140
rect 283190 159128 283196 159140
rect 283248 159128 283254 159180
rect 284662 159128 284668 159180
rect 284720 159168 284726 159180
rect 285766 159168 285772 159180
rect 284720 159140 285772 159168
rect 284720 159128 284726 159140
rect 285766 159128 285772 159140
rect 285824 159128 285830 159180
rect 288250 159168 288256 159180
rect 287026 159140 288256 159168
rect 180392 159072 197124 159100
rect 200086 159072 207060 159100
rect 180392 159060 180398 159072
rect 107194 158992 107200 159044
rect 107252 159032 107258 159044
rect 185578 159032 185584 159044
rect 107252 159004 185584 159032
rect 107252 158992 107258 159004
rect 185578 158992 185584 159004
rect 185636 158992 185642 159044
rect 193582 158992 193588 159044
rect 193640 159032 193646 159044
rect 196986 159032 196992 159044
rect 193640 159004 196992 159032
rect 193640 158992 193646 159004
rect 196986 158992 196992 159004
rect 197044 158992 197050 159044
rect 73522 158924 73528 158976
rect 73580 158964 73586 158976
rect 107562 158964 107568 158976
rect 73580 158936 107568 158964
rect 73580 158924 73586 158936
rect 107562 158924 107568 158936
rect 107620 158924 107626 158976
rect 119798 158924 119804 158976
rect 119856 158964 119862 158976
rect 127618 158964 127624 158976
rect 119856 158936 127624 158964
rect 119856 158924 119862 158936
rect 127618 158924 127624 158936
rect 127676 158924 127682 158976
rect 192662 158964 192668 158976
rect 127728 158936 192668 158964
rect 96246 158856 96252 158908
rect 96304 158896 96310 158908
rect 121822 158896 121828 158908
rect 96304 158868 121828 158896
rect 96304 158856 96310 158868
rect 121822 158856 121828 158868
rect 121880 158856 121886 158908
rect 124030 158856 124036 158908
rect 124088 158896 124094 158908
rect 127728 158896 127756 158936
rect 192662 158924 192668 158936
rect 192720 158924 192726 158976
rect 124088 158868 127756 158896
rect 124088 158856 124094 158868
rect 130746 158856 130752 158908
rect 130804 158896 130810 158908
rect 195146 158896 195152 158908
rect 130804 158868 195152 158896
rect 130804 158856 130810 158868
rect 195146 158856 195152 158868
rect 195204 158856 195210 158908
rect 197096 158896 197124 159072
rect 207382 159060 207388 159112
rect 207440 159100 207446 159112
rect 212718 159100 212724 159112
rect 207440 159072 212724 159100
rect 207440 159060 207446 159072
rect 212718 159060 212724 159072
rect 212776 159060 212782 159112
rect 212810 159060 212816 159112
rect 212868 159100 212874 159112
rect 222102 159100 222108 159112
rect 212868 159072 222108 159100
rect 212868 159060 212874 159072
rect 222102 159060 222108 159072
rect 222160 159060 222166 159112
rect 224126 159060 224132 159112
rect 224184 159100 224190 159112
rect 287026 159100 287054 159140
rect 288250 159128 288256 159140
rect 288308 159128 288314 159180
rect 288894 159128 288900 159180
rect 288952 159168 288958 159180
rect 338390 159168 338396 159180
rect 288952 159140 338396 159168
rect 288952 159128 288958 159140
rect 338390 159128 338396 159140
rect 338448 159128 338454 159180
rect 338482 159128 338488 159180
rect 338540 159168 338546 159180
rect 340782 159168 340788 159180
rect 338540 159140 340788 159168
rect 338540 159128 338546 159140
rect 340782 159128 340788 159140
rect 340840 159128 340846 159180
rect 341886 159128 341892 159180
rect 341944 159168 341950 159180
rect 378226 159168 378232 159180
rect 341944 159140 378232 159168
rect 341944 159128 341950 159140
rect 378226 159128 378232 159140
rect 378284 159128 378290 159180
rect 457898 159128 457904 159180
rect 457956 159168 457962 159180
rect 463878 159168 463884 159180
rect 457956 159140 463884 159168
rect 457956 159128 457962 159140
rect 463878 159128 463884 159140
rect 463936 159128 463942 159180
rect 224184 159072 287054 159100
rect 224184 159060 224190 159072
rect 307386 159060 307392 159112
rect 307444 159100 307450 159112
rect 349338 159100 349344 159112
rect 307444 159072 349344 159100
rect 307444 159060 307450 159072
rect 349338 159060 349344 159072
rect 349396 159060 349402 159112
rect 351086 159060 351092 159112
rect 351144 159100 351150 159112
rect 382274 159100 382280 159112
rect 351144 159072 382280 159100
rect 351144 159060 351150 159072
rect 382274 159060 382280 159072
rect 382332 159060 382338 159112
rect 409138 159060 409144 159112
rect 409196 159100 409202 159112
rect 410886 159100 410892 159112
rect 409196 159072 410892 159100
rect 409196 159060 409202 159072
rect 410886 159060 410892 159072
rect 410944 159060 410950 159112
rect 452838 159060 452844 159112
rect 452896 159100 452902 159112
rect 459646 159100 459652 159112
rect 452896 159072 459652 159100
rect 452896 159060 452902 159072
rect 459646 159060 459652 159072
rect 459704 159060 459710 159112
rect 461302 159060 461308 159112
rect 461360 159100 461366 159112
rect 467834 159100 467840 159112
rect 461360 159072 467840 159100
rect 461360 159060 461366 159072
rect 467834 159060 467840 159072
rect 467892 159060 467898 159112
rect 200574 158992 200580 159044
rect 200632 159032 200638 159044
rect 227714 159032 227720 159044
rect 200632 159004 212764 159032
rect 200632 158992 200638 159004
rect 197170 158924 197176 158976
rect 197228 158964 197234 158976
rect 212626 158964 212632 158976
rect 197228 158936 212632 158964
rect 197228 158924 197234 158936
rect 212626 158924 212632 158936
rect 212684 158924 212690 158976
rect 212736 158964 212764 159004
rect 215266 159004 227720 159032
rect 215266 158964 215294 159004
rect 227714 158992 227720 159004
rect 227772 158992 227778 159044
rect 230842 158992 230848 159044
rect 230900 159032 230906 159044
rect 295150 159032 295156 159044
rect 230900 159004 295156 159032
rect 230900 158992 230906 159004
rect 295150 158992 295156 159004
rect 295208 158992 295214 159044
rect 298094 158992 298100 159044
rect 298152 159032 298158 159044
rect 300762 159032 300768 159044
rect 298152 159004 300768 159032
rect 298152 158992 298158 159004
rect 300762 158992 300768 159004
rect 300820 158992 300826 159044
rect 308214 158992 308220 159044
rect 308272 159032 308278 159044
rect 347682 159032 347688 159044
rect 308272 159004 347688 159032
rect 308272 158992 308278 159004
rect 347682 158992 347688 159004
rect 347740 158992 347746 159044
rect 347774 158992 347780 159044
rect 347832 159032 347838 159044
rect 378778 159032 378784 159044
rect 347832 159004 378784 159032
rect 347832 158992 347838 159004
rect 378778 158992 378784 159004
rect 378836 158992 378842 159044
rect 384666 158992 384672 159044
rect 384724 159032 384730 159044
rect 388438 159032 388444 159044
rect 384724 159004 388444 159032
rect 384724 158992 384730 159004
rect 388438 158992 388444 159004
rect 388496 158992 388502 159044
rect 388990 158992 388996 159044
rect 389048 159032 389054 159044
rect 403250 159032 403256 159044
rect 389048 159004 403256 159032
rect 389048 158992 389054 159004
rect 403250 158992 403256 159004
rect 403308 158992 403314 159044
rect 455414 158992 455420 159044
rect 455472 159032 455478 159044
rect 463510 159032 463516 159044
rect 455472 159004 463516 159032
rect 455472 158992 455478 159004
rect 463510 158992 463516 159004
rect 463568 158992 463574 159044
rect 465534 158992 465540 159044
rect 465592 159032 465598 159044
rect 472434 159032 472440 159044
rect 465592 159004 472440 159032
rect 465592 158992 465598 159004
rect 472434 158992 472440 159004
rect 472492 158992 472498 159044
rect 473906 158992 473912 159044
rect 473964 159032 473970 159044
rect 480254 159032 480260 159044
rect 473964 159004 480260 159032
rect 473964 158992 473970 159004
rect 480254 158992 480260 159004
rect 480312 158992 480318 159044
rect 212736 158936 215294 158964
rect 217318 158924 217324 158976
rect 217376 158964 217382 158976
rect 220446 158964 220452 158976
rect 217376 158936 220452 158964
rect 217376 158924 217382 158936
rect 220446 158924 220452 158936
rect 220504 158924 220510 158976
rect 237558 158924 237564 158976
rect 237616 158964 237622 158976
rect 299474 158964 299480 158976
rect 237616 158936 299480 158964
rect 237616 158924 237622 158936
rect 299474 158924 299480 158936
rect 299532 158924 299538 158976
rect 301406 158924 301412 158976
rect 301464 158964 301470 158976
rect 308582 158964 308588 158976
rect 301464 158936 308588 158964
rect 301464 158924 301470 158936
rect 308582 158924 308588 158936
rect 308640 158924 308646 158976
rect 314930 158924 314936 158976
rect 314988 158964 314994 158976
rect 357434 158964 357440 158976
rect 314988 158936 357440 158964
rect 314988 158924 314994 158936
rect 357434 158924 357440 158936
rect 357492 158924 357498 158976
rect 361206 158924 361212 158976
rect 361264 158964 361270 158976
rect 361264 158936 367876 158964
rect 361264 158924 361270 158936
rect 201402 158896 201408 158908
rect 197096 158868 201408 158896
rect 201402 158856 201408 158868
rect 201460 158856 201466 158908
rect 207290 158856 207296 158908
rect 207348 158896 207354 158908
rect 231762 158896 231768 158908
rect 207348 158868 231768 158896
rect 207348 158856 207354 158868
rect 231762 158856 231768 158868
rect 231820 158856 231826 158908
rect 238386 158856 238392 158908
rect 238444 158896 238450 158908
rect 242802 158896 242808 158908
rect 238444 158868 242808 158896
rect 238444 158856 238450 158868
rect 242802 158856 242808 158868
rect 242860 158856 242866 158908
rect 244274 158856 244280 158908
rect 244332 158896 244338 158908
rect 305362 158896 305368 158908
rect 244332 158868 305368 158896
rect 244332 158856 244338 158868
rect 305362 158856 305368 158868
rect 305420 158856 305426 158908
rect 305638 158856 305644 158908
rect 305696 158896 305702 158908
rect 307662 158896 307668 158908
rect 305696 158868 307668 158896
rect 305696 158856 305702 158868
rect 307662 158856 307668 158868
rect 307720 158856 307726 158908
rect 310698 158856 310704 158908
rect 310756 158896 310762 158908
rect 311986 158896 311992 158908
rect 310756 158868 311992 158896
rect 310756 158856 310762 158868
rect 311986 158856 311992 158868
rect 312044 158856 312050 158908
rect 312446 158856 312452 158908
rect 312504 158896 312510 158908
rect 313458 158896 313464 158908
rect 312504 158868 313464 158896
rect 312504 158856 312510 158868
rect 313458 158856 313464 158868
rect 313516 158856 313522 158908
rect 322474 158856 322480 158908
rect 322532 158896 322538 158908
rect 365162 158896 365168 158908
rect 322532 158868 365168 158896
rect 322532 158856 322538 158868
rect 365162 158856 365168 158868
rect 365220 158856 365226 158908
rect 102962 158788 102968 158840
rect 103020 158828 103026 158840
rect 125502 158828 125508 158840
rect 103020 158800 125508 158828
rect 103020 158788 103026 158800
rect 125502 158788 125508 158800
rect 125560 158788 125566 158840
rect 126514 158788 126520 158840
rect 126572 158828 126578 158840
rect 154482 158828 154488 158840
rect 126572 158800 154488 158828
rect 126572 158788 126578 158800
rect 154482 158788 154488 158800
rect 154540 158788 154546 158840
rect 156782 158788 156788 158840
rect 156840 158828 156846 158840
rect 194502 158828 194508 158840
rect 156840 158800 194508 158828
rect 156840 158788 156846 158800
rect 194502 158788 194508 158800
rect 194560 158788 194566 158840
rect 194686 158788 194692 158840
rect 194744 158828 194750 158840
rect 203702 158828 203708 158840
rect 194744 158800 203708 158828
rect 194744 158788 194750 158800
rect 203702 158788 203708 158800
rect 203760 158788 203766 158840
rect 206922 158788 206928 158840
rect 206980 158828 206986 158840
rect 213822 158828 213828 158840
rect 206980 158800 213828 158828
rect 206980 158788 206986 158800
rect 213822 158788 213828 158800
rect 213880 158788 213886 158840
rect 214834 158788 214840 158840
rect 214892 158828 214898 158840
rect 221734 158828 221740 158840
rect 214892 158800 221740 158828
rect 214892 158788 214898 158800
rect 221734 158788 221740 158800
rect 221792 158788 221798 158840
rect 261110 158788 261116 158840
rect 261168 158828 261174 158840
rect 317046 158828 317052 158840
rect 261168 158800 317052 158828
rect 261168 158788 261174 158800
rect 317046 158788 317052 158800
rect 317104 158788 317110 158840
rect 320266 158828 320272 158840
rect 319088 158800 320272 158828
rect 106366 158720 106372 158772
rect 106424 158760 106430 158772
rect 127250 158760 127256 158772
rect 106424 158732 127256 158760
rect 106424 158720 106430 158732
rect 127250 158720 127256 158732
rect 127308 158720 127314 158772
rect 127342 158720 127348 158772
rect 127400 158760 127406 158772
rect 129734 158760 129740 158772
rect 127400 158732 129740 158760
rect 127400 158720 127406 158732
rect 129734 158720 129740 158732
rect 129792 158720 129798 158772
rect 133230 158720 133236 158772
rect 133288 158760 133294 158772
rect 158714 158760 158720 158772
rect 133288 158732 158720 158760
rect 133288 158720 133294 158732
rect 158714 158720 158720 158732
rect 158772 158720 158778 158772
rect 163148 158732 167776 158760
rect 81066 158652 81072 158704
rect 81124 158692 81130 158704
rect 163038 158692 163044 158704
rect 81124 158664 163044 158692
rect 81124 158652 81130 158664
rect 163038 158652 163044 158664
rect 163096 158652 163102 158704
rect 67634 158584 67640 158636
rect 67692 158624 67698 158636
rect 163148 158624 163176 158732
rect 163222 158652 163228 158704
rect 163280 158692 163286 158704
rect 167638 158692 167644 158704
rect 163280 158664 167644 158692
rect 163280 158652 163286 158664
rect 167638 158652 167644 158664
rect 167696 158652 167702 158704
rect 67692 158596 163176 158624
rect 67692 158584 67698 158596
rect 163314 158584 163320 158636
rect 163372 158624 163378 158636
rect 167546 158624 167552 158636
rect 163372 158596 167552 158624
rect 163372 158584 163378 158596
rect 167546 158584 167552 158596
rect 167604 158584 167610 158636
rect 167748 158624 167776 158732
rect 171134 158720 171140 158772
rect 171192 158760 171198 158772
rect 172606 158760 172612 158772
rect 171192 158732 172612 158760
rect 171192 158720 171198 158732
rect 172606 158720 172612 158732
rect 172664 158720 172670 158772
rect 175826 158720 175832 158772
rect 175884 158760 175890 158772
rect 176654 158760 176660 158772
rect 175884 158732 176660 158760
rect 175884 158720 175890 158732
rect 176654 158720 176660 158732
rect 176712 158720 176718 158772
rect 180702 158720 180708 158772
rect 180760 158760 180766 158772
rect 180760 158732 181024 158760
rect 180760 158720 180766 158732
rect 167822 158652 167828 158704
rect 167880 158692 167886 158704
rect 180886 158692 180892 158704
rect 167880 158664 180892 158692
rect 167880 158652 167886 158664
rect 180886 158652 180892 158664
rect 180944 158652 180950 158704
rect 180996 158692 181024 158732
rect 183738 158720 183744 158772
rect 183796 158760 183802 158772
rect 204898 158760 204904 158772
rect 183796 158732 204904 158760
rect 183796 158720 183802 158732
rect 204898 158720 204904 158732
rect 204956 158720 204962 158772
rect 210602 158720 210608 158772
rect 210660 158760 210666 158772
rect 215386 158760 215392 158772
rect 210660 158732 215392 158760
rect 210660 158720 210666 158732
rect 215386 158720 215392 158732
rect 215444 158720 215450 158772
rect 221550 158720 221556 158772
rect 221608 158760 221614 158772
rect 223850 158760 223856 158772
rect 221608 158732 223856 158760
rect 221608 158720 221614 158732
rect 223850 158720 223856 158732
rect 223908 158720 223914 158772
rect 240870 158720 240876 158772
rect 240928 158760 240934 158772
rect 243354 158760 243360 158772
rect 240928 158732 243360 158760
rect 240928 158720 240934 158732
rect 243354 158720 243360 158732
rect 243412 158720 243418 158772
rect 254394 158720 254400 158772
rect 254452 158760 254458 158772
rect 255498 158760 255504 158772
rect 254452 158732 255504 158760
rect 254452 158720 254458 158732
rect 255498 158720 255504 158732
rect 255556 158720 255562 158772
rect 258534 158720 258540 158772
rect 258592 158760 258598 158772
rect 261018 158760 261024 158772
rect 258592 158732 261024 158760
rect 258592 158720 258598 158732
rect 261018 158720 261024 158732
rect 261076 158720 261082 158772
rect 264422 158720 264428 158772
rect 264480 158760 264486 158772
rect 266354 158760 266360 158772
rect 264480 158732 266360 158760
rect 264480 158720 264486 158732
rect 266354 158720 266360 158732
rect 266412 158720 266418 158772
rect 267826 158720 267832 158772
rect 267884 158760 267890 158772
rect 319088 158760 319116 158800
rect 320266 158788 320272 158800
rect 320324 158788 320330 158840
rect 327534 158788 327540 158840
rect 327592 158828 327598 158840
rect 330478 158828 330484 158840
rect 327592 158800 330484 158828
rect 327592 158788 327598 158800
rect 330478 158788 330484 158800
rect 330536 158788 330542 158840
rect 363138 158828 363144 158840
rect 330588 158800 363144 158828
rect 267884 158732 319116 158760
rect 267884 158720 267890 158732
rect 319162 158720 319168 158772
rect 319220 158760 319226 158772
rect 321554 158760 321560 158772
rect 319220 158732 321560 158760
rect 319220 158720 319226 158732
rect 321554 158720 321560 158732
rect 321612 158720 321618 158772
rect 321646 158720 321652 158772
rect 321704 158760 321710 158772
rect 321704 158732 330432 158760
rect 321704 158720 321710 158732
rect 181714 158692 181720 158704
rect 180996 158664 181720 158692
rect 181714 158652 181720 158664
rect 181772 158652 181778 158704
rect 181990 158652 181996 158704
rect 182048 158692 182054 158704
rect 256786 158692 256792 158704
rect 182048 158664 256792 158692
rect 182048 158652 182054 158664
rect 256786 158652 256792 158664
rect 256844 158652 256850 158704
rect 330404 158692 330432 158732
rect 330588 158692 330616 158800
rect 363138 158788 363144 158800
rect 363196 158788 363202 158840
rect 367848 158828 367876 158936
rect 369210 158924 369216 158976
rect 369268 158964 369274 158976
rect 384942 158964 384948 158976
rect 369268 158936 384948 158964
rect 369268 158924 369274 158936
rect 384942 158924 384948 158936
rect 385000 158924 385006 158976
rect 420086 158924 420092 158976
rect 420144 158964 420150 158976
rect 423582 158964 423588 158976
rect 420144 158936 423588 158964
rect 420144 158924 420150 158936
rect 423582 158924 423588 158936
rect 423640 158924 423646 158976
rect 446122 158924 446128 158976
rect 446180 158964 446186 158976
rect 453850 158964 453856 158976
rect 446180 158936 453856 158964
rect 446180 158924 446186 158936
rect 453850 158924 453856 158936
rect 453908 158924 453914 158976
rect 454586 158924 454592 158976
rect 454644 158964 454650 158976
rect 461854 158964 461860 158976
rect 454644 158936 461860 158964
rect 454644 158924 454650 158936
rect 461854 158924 461860 158936
rect 461912 158924 461918 158976
rect 464614 158924 464620 158976
rect 464672 158964 464678 158976
rect 471238 158964 471244 158976
rect 464672 158936 471244 158964
rect 464672 158924 464678 158936
rect 471238 158924 471244 158936
rect 471296 158924 471302 158976
rect 475562 158924 475568 158976
rect 475620 158964 475626 158976
rect 482002 158964 482008 158976
rect 475620 158936 482008 158964
rect 475620 158924 475626 158936
rect 482002 158924 482008 158936
rect 482060 158924 482066 158976
rect 367922 158856 367928 158908
rect 367980 158896 367986 158908
rect 386230 158896 386236 158908
rect 367980 158868 386236 158896
rect 367980 158856 367986 158868
rect 386230 158856 386236 158868
rect 386288 158856 386294 158908
rect 391474 158856 391480 158908
rect 391532 158896 391538 158908
rect 394326 158896 394332 158908
rect 391532 158868 394332 158896
rect 391532 158856 391538 158868
rect 394326 158856 394332 158868
rect 394384 158856 394390 158908
rect 412542 158856 412548 158908
rect 412600 158896 412606 158908
rect 413094 158896 413100 158908
rect 412600 158868 413100 158896
rect 412600 158856 412606 158868
rect 413094 158856 413100 158868
rect 413152 158856 413158 158908
rect 456242 158856 456248 158908
rect 456300 158896 456306 158908
rect 462958 158896 462964 158908
rect 456300 158868 462964 158896
rect 456300 158856 456306 158868
rect 462958 158856 462964 158868
rect 463016 158856 463022 158908
rect 466362 158856 466368 158908
rect 466420 158896 466426 158908
rect 472342 158896 472348 158908
rect 466420 158868 472348 158896
rect 466420 158856 466426 158868
rect 472342 158856 472348 158868
rect 472400 158856 472406 158908
rect 474734 158856 474740 158908
rect 474792 158896 474798 158908
rect 481358 158896 481364 158908
rect 474792 158868 481364 158896
rect 474792 158856 474798 158868
rect 481358 158856 481364 158868
rect 481416 158856 481422 158908
rect 481450 158856 481456 158908
rect 481508 158896 481514 158908
rect 486510 158896 486516 158908
rect 481508 158868 486516 158896
rect 481508 158856 481514 158868
rect 486510 158856 486516 158868
rect 486568 158856 486574 158908
rect 508314 158856 508320 158908
rect 508372 158896 508378 158908
rect 510062 158896 510068 158908
rect 508372 158868 510068 158896
rect 508372 158856 508378 158868
rect 510062 158856 510068 158868
rect 510120 158856 510126 158908
rect 385770 158828 385776 158840
rect 367848 158800 385776 158828
rect 385770 158788 385776 158800
rect 385828 158788 385834 158840
rect 388070 158788 388076 158840
rect 388128 158828 388134 158840
rect 390370 158828 390376 158840
rect 388128 158800 390376 158828
rect 388128 158788 388134 158800
rect 390370 158788 390376 158800
rect 390428 158788 390434 158840
rect 405734 158788 405740 158840
rect 405792 158828 405798 158840
rect 409230 158828 409236 158840
rect 405792 158800 409236 158828
rect 405792 158788 405798 158800
rect 409230 158788 409236 158800
rect 409288 158788 409294 158840
rect 413370 158788 413376 158840
rect 413428 158828 413434 158840
rect 419626 158828 419632 158840
rect 413428 158800 419632 158828
rect 413428 158788 413434 158800
rect 419626 158788 419632 158800
rect 419684 158788 419690 158840
rect 463786 158788 463792 158840
rect 463844 158828 463850 158840
rect 471422 158828 471428 158840
rect 463844 158800 471428 158828
rect 463844 158788 463850 158800
rect 471422 158788 471428 158800
rect 471480 158788 471486 158840
rect 476390 158788 476396 158840
rect 476448 158828 476454 158840
rect 481634 158828 481640 158840
rect 476448 158800 481640 158828
rect 476448 158788 476454 158800
rect 481634 158788 481640 158800
rect 481692 158788 481698 158840
rect 505278 158788 505284 158840
rect 505336 158828 505342 158840
rect 507578 158828 507584 158840
rect 505336 158800 507584 158828
rect 505336 158788 505342 158800
rect 507578 158788 507584 158800
rect 507636 158788 507642 158840
rect 330662 158720 330668 158772
rect 330720 158760 330726 158772
rect 367186 158760 367192 158772
rect 330720 158732 367192 158760
rect 330720 158720 330726 158732
rect 367186 158720 367192 158732
rect 367244 158720 367250 158772
rect 374638 158720 374644 158772
rect 374696 158760 374702 158772
rect 384666 158760 384672 158772
rect 374696 158732 384672 158760
rect 374696 158720 374702 158732
rect 384666 158720 384672 158732
rect 384724 158720 384730 158772
rect 384758 158720 384764 158772
rect 384816 158760 384822 158772
rect 389174 158760 389180 158772
rect 384816 158732 389180 158760
rect 384816 158720 384822 158732
rect 389174 158720 389180 158732
rect 389232 158720 389238 158772
rect 416682 158720 416688 158772
rect 416740 158760 416746 158772
rect 419534 158760 419540 158772
rect 416740 158732 419540 158760
rect 416740 158720 416746 158732
rect 419534 158720 419540 158732
rect 419592 158720 419598 158772
rect 452010 158720 452016 158772
rect 452068 158760 452074 158772
rect 458174 158760 458180 158772
rect 452068 158732 458180 158760
rect 452068 158720 452074 158732
rect 458174 158720 458180 158732
rect 458232 158720 458238 158772
rect 462130 158720 462136 158772
rect 462188 158760 462194 158772
rect 467926 158760 467932 158772
rect 462188 158732 467932 158760
rect 462188 158720 462194 158732
rect 467926 158720 467932 158732
rect 467984 158720 467990 158772
rect 473078 158720 473084 158772
rect 473136 158760 473142 158772
rect 478966 158760 478972 158772
rect 473136 158732 478972 158760
rect 473136 158720 473142 158732
rect 478966 158720 478972 158732
rect 479024 158720 479030 158772
rect 482278 158720 482284 158772
rect 482336 158760 482342 158772
rect 487246 158760 487252 158772
rect 482336 158732 487252 158760
rect 482336 158720 482342 158732
rect 487246 158720 487252 158732
rect 487304 158720 487310 158772
rect 505738 158720 505744 158772
rect 505796 158760 505802 158772
rect 506750 158760 506756 158772
rect 505796 158732 506756 158760
rect 505796 158720 505802 158732
rect 506750 158720 506756 158732
rect 506808 158720 506814 158772
rect 507026 158720 507032 158772
rect 507084 158760 507090 158772
rect 508406 158760 508412 158772
rect 507084 158732 508412 158760
rect 507084 158720 507090 158732
rect 508406 158720 508412 158732
rect 508464 158720 508470 158772
rect 509418 158720 509424 158772
rect 509476 158760 509482 158772
rect 511718 158760 511724 158772
rect 509476 158732 511724 158760
rect 509476 158720 509482 158732
rect 511718 158720 511724 158732
rect 511776 158720 511782 158772
rect 514938 158720 514944 158772
rect 514996 158760 515002 158772
rect 518526 158760 518532 158772
rect 514996 158732 518532 158760
rect 514996 158720 515002 158732
rect 518526 158720 518532 158732
rect 518584 158720 518590 158772
rect 330404 158664 330616 158692
rect 170306 158624 170312 158636
rect 167748 158596 170312 158624
rect 170306 158584 170312 158596
rect 170364 158584 170370 158636
rect 171962 158584 171968 158636
rect 172020 158624 172026 158636
rect 250070 158624 250076 158636
rect 172020 158596 250076 158624
rect 172020 158584 172026 158596
rect 250070 158584 250076 158596
rect 250128 158584 250134 158636
rect 74350 158516 74356 158568
rect 74408 158556 74414 158568
rect 74408 158528 173296 158556
rect 74408 158516 74414 158528
rect 71038 158448 71044 158500
rect 71096 158488 71102 158500
rect 173066 158488 173072 158500
rect 71096 158460 173072 158488
rect 71096 158448 71102 158460
rect 173066 158448 173072 158460
rect 173124 158448 173130 158500
rect 173268 158488 173296 158528
rect 175274 158516 175280 158568
rect 175332 158556 175338 158568
rect 252738 158556 252744 158568
rect 175332 158528 252744 158556
rect 175332 158516 175338 158528
rect 252738 158516 252744 158528
rect 252796 158516 252802 158568
rect 175366 158488 175372 158500
rect 173268 158460 175372 158488
rect 175366 158448 175372 158460
rect 175424 158448 175430 158500
rect 178678 158448 178684 158500
rect 178736 158488 178742 158500
rect 255406 158488 255412 158500
rect 178736 158460 255412 158488
rect 178736 158448 178742 158460
rect 255406 158448 255412 158460
rect 255464 158448 255470 158500
rect 64230 158380 64236 158432
rect 64288 158420 64294 158432
rect 163314 158420 163320 158432
rect 64288 158392 163320 158420
rect 64288 158380 64294 158392
rect 163314 158380 163320 158392
rect 163372 158380 163378 158432
rect 165430 158420 165436 158432
rect 163424 158392 165436 158420
rect 60918 158312 60924 158364
rect 60976 158352 60982 158364
rect 163424 158352 163452 158392
rect 165430 158380 165436 158392
rect 165488 158380 165494 158432
rect 168558 158380 168564 158432
rect 168616 158420 168622 158432
rect 247126 158420 247132 158432
rect 168616 158392 247132 158420
rect 168616 158380 168622 158392
rect 247126 158380 247132 158392
rect 247184 158380 247190 158432
rect 60976 158324 163452 158352
rect 60976 158312 60982 158324
rect 165246 158312 165252 158364
rect 165304 158352 165310 158364
rect 245010 158352 245016 158364
rect 165304 158324 245016 158352
rect 165304 158312 165310 158324
rect 245010 158312 245016 158324
rect 245068 158312 245074 158364
rect 54202 158244 54208 158296
rect 54260 158284 54266 158296
rect 160278 158284 160284 158296
rect 54260 158256 160284 158284
rect 54260 158244 54266 158256
rect 160278 158244 160284 158256
rect 160336 158244 160342 158296
rect 161842 158244 161848 158296
rect 161900 158284 161906 158296
rect 242066 158284 242072 158296
rect 161900 158256 242072 158284
rect 161900 158244 161906 158256
rect 242066 158244 242072 158256
rect 242124 158244 242130 158296
rect 50798 158176 50804 158228
rect 50856 158216 50862 158228
rect 157702 158216 157708 158228
rect 50856 158188 157708 158216
rect 50856 158176 50862 158188
rect 157702 158176 157708 158188
rect 157760 158176 157766 158228
rect 158438 158176 158444 158228
rect 158496 158216 158502 158228
rect 238938 158216 238944 158228
rect 158496 158188 238944 158216
rect 158496 158176 158502 158188
rect 238938 158176 238944 158188
rect 238996 158176 239002 158228
rect 256878 158176 256884 158228
rect 256936 158216 256942 158228
rect 315022 158216 315028 158228
rect 256936 158188 315028 158216
rect 256936 158176 256942 158188
rect 315022 158176 315028 158188
rect 315080 158176 315086 158228
rect 47486 158108 47492 158160
rect 47544 158148 47550 158160
rect 155034 158148 155040 158160
rect 47544 158120 155040 158148
rect 47544 158108 47550 158120
rect 155034 158108 155040 158120
rect 155092 158108 155098 158160
rect 155126 158108 155132 158160
rect 155184 158148 155190 158160
rect 237374 158148 237380 158160
rect 155184 158120 237380 158148
rect 155184 158108 155190 158120
rect 237374 158108 237380 158120
rect 237432 158108 237438 158160
rect 246758 158108 246764 158160
rect 246816 158148 246822 158160
rect 306926 158148 306932 158160
rect 246816 158120 306932 158148
rect 246816 158108 246822 158120
rect 306926 158108 306932 158120
rect 306984 158108 306990 158160
rect 37366 158040 37372 158092
rect 37424 158080 37430 158092
rect 146386 158080 146392 158092
rect 37424 158052 146392 158080
rect 37424 158040 37430 158052
rect 146386 158040 146392 158052
rect 146444 158040 146450 158092
rect 148410 158040 148416 158092
rect 148468 158080 148474 158092
rect 231946 158080 231952 158092
rect 148468 158052 231952 158080
rect 148468 158040 148474 158052
rect 231946 158040 231952 158052
rect 232004 158040 232010 158092
rect 233326 158040 233332 158092
rect 233384 158080 233390 158092
rect 297082 158080 297088 158092
rect 233384 158052 297088 158080
rect 233384 158040 233390 158052
rect 297082 158040 297088 158052
rect 297140 158040 297146 158092
rect 300670 158040 300676 158092
rect 300728 158080 300734 158092
rect 348050 158080 348056 158092
rect 300728 158052 348056 158080
rect 300728 158040 300734 158052
rect 348050 158040 348056 158052
rect 348108 158040 348114 158092
rect 382 157972 388 158024
rect 440 158012 446 158024
rect 118878 158012 118884 158024
rect 440 157984 118884 158012
rect 440 157972 446 157984
rect 118878 157972 118884 157984
rect 118936 157972 118942 158024
rect 127250 157972 127256 158024
rect 127308 158012 127314 158024
rect 127894 158012 127900 158024
rect 127308 157984 127900 158012
rect 127308 157972 127314 157984
rect 127894 157972 127900 157984
rect 127952 157972 127958 158024
rect 131574 157972 131580 158024
rect 131632 158012 131638 158024
rect 219342 158012 219348 158024
rect 131632 157984 219348 158012
rect 131632 157972 131638 157984
rect 219342 157972 219348 157984
rect 219400 157972 219406 158024
rect 240042 157972 240048 158024
rect 240100 158012 240106 158024
rect 302234 158012 302240 158024
rect 240100 157984 302240 158012
rect 240100 157972 240106 157984
rect 302234 157972 302240 157984
rect 302292 157972 302298 158024
rect 77754 157904 77760 157956
rect 77812 157944 77818 157956
rect 77812 157916 176056 157944
rect 77812 157904 77818 157916
rect 84470 157836 84476 157888
rect 84528 157876 84534 157888
rect 175918 157876 175924 157888
rect 84528 157848 175924 157876
rect 84528 157836 84534 157848
rect 175918 157836 175924 157848
rect 175976 157836 175982 157888
rect 176028 157876 176056 157916
rect 176194 157904 176200 157956
rect 176252 157944 176258 157956
rect 182266 157944 182272 157956
rect 176252 157916 182272 157944
rect 176252 157904 176258 157916
rect 182266 157904 182272 157916
rect 182324 157904 182330 157956
rect 185394 157904 185400 157956
rect 185452 157944 185458 157956
rect 260466 157944 260472 157956
rect 185452 157916 260472 157944
rect 185452 157904 185458 157916
rect 260466 157904 260472 157916
rect 260524 157904 260530 157956
rect 178034 157876 178040 157888
rect 176028 157848 178040 157876
rect 178034 157836 178040 157848
rect 178092 157836 178098 157888
rect 188522 157876 188528 157888
rect 181456 157848 188528 157876
rect 87782 157768 87788 157820
rect 87840 157808 87846 157820
rect 181346 157808 181352 157820
rect 87840 157780 181352 157808
rect 87840 157768 87846 157780
rect 181346 157768 181352 157780
rect 181404 157768 181410 157820
rect 91186 157700 91192 157752
rect 91244 157740 91250 157752
rect 181456 157740 181484 157848
rect 188522 157836 188528 157848
rect 188580 157836 188586 157888
rect 188798 157836 188804 157888
rect 188856 157876 188862 157888
rect 263042 157876 263048 157888
rect 188856 157848 263048 157876
rect 188856 157836 188862 157848
rect 263042 157836 263048 157848
rect 263100 157836 263106 157888
rect 190638 157808 190644 157820
rect 91244 157712 181484 157740
rect 181548 157780 190644 157808
rect 91244 157700 91250 157712
rect 94590 157632 94596 157684
rect 94648 157672 94654 157684
rect 181548 157672 181576 157780
rect 190638 157768 190644 157780
rect 190696 157768 190702 157820
rect 195514 157768 195520 157820
rect 195572 157808 195578 157820
rect 267734 157808 267740 157820
rect 195572 157780 267740 157808
rect 195572 157768 195578 157780
rect 267734 157768 267740 157780
rect 267792 157768 267798 157820
rect 181714 157700 181720 157752
rect 181772 157740 181778 157752
rect 181772 157712 186314 157740
rect 181772 157700 181778 157712
rect 94648 157644 181576 157672
rect 94648 157632 94654 157644
rect 181622 157632 181628 157684
rect 181680 157672 181686 157684
rect 185394 157672 185400 157684
rect 181680 157644 185400 157672
rect 181680 157632 181686 157644
rect 185394 157632 185400 157644
rect 185452 157632 185458 157684
rect 186286 157672 186314 157712
rect 190454 157700 190460 157752
rect 190512 157740 190518 157752
rect 263686 157740 263692 157752
rect 190512 157712 263692 157740
rect 190512 157700 190518 157712
rect 263686 157700 263692 157712
rect 263744 157700 263750 157752
rect 236178 157672 236184 157684
rect 186286 157644 236184 157672
rect 236178 157632 236184 157644
rect 236236 157632 236242 157684
rect 97902 157564 97908 157616
rect 97960 157604 97966 157616
rect 193214 157604 193220 157616
rect 97960 157576 193220 157604
rect 97960 157564 97966 157576
rect 193214 157564 193220 157576
rect 193272 157564 193278 157616
rect 197354 157564 197360 157616
rect 197412 157604 197418 157616
rect 251450 157604 251456 157616
rect 197412 157576 251456 157604
rect 197412 157564 197418 157576
rect 251450 157564 251456 157576
rect 251508 157564 251514 157616
rect 111334 157496 111340 157548
rect 111392 157536 111398 157548
rect 203426 157536 203432 157548
rect 111392 157508 203432 157536
rect 111392 157496 111398 157508
rect 203426 157496 203432 157508
rect 203484 157496 203490 157548
rect 204898 157496 204904 157548
rect 204956 157536 204962 157548
rect 258074 157536 258080 157548
rect 204956 157508 258080 157536
rect 204956 157496 204962 157508
rect 258074 157496 258080 157508
rect 258132 157496 258138 157548
rect 114738 157428 114744 157480
rect 114796 157468 114802 157480
rect 206554 157468 206560 157480
rect 114796 157440 206560 157468
rect 114796 157428 114802 157440
rect 206554 157428 206560 157440
rect 206612 157428 206618 157480
rect 141694 157360 141700 157412
rect 141752 157400 141758 157412
rect 227070 157400 227076 157412
rect 141752 157372 227076 157400
rect 141752 157360 141758 157372
rect 227070 157360 227076 157372
rect 227128 157360 227134 157412
rect 52454 157292 52460 157344
rect 52512 157332 52518 157344
rect 158622 157332 158628 157344
rect 52512 157304 158628 157332
rect 52512 157292 52518 157304
rect 158622 157292 158628 157304
rect 158680 157292 158686 157344
rect 158714 157292 158720 157344
rect 158772 157332 158778 157344
rect 158772 157304 203932 157332
rect 158772 157292 158778 157304
rect 55858 157224 55864 157276
rect 55916 157264 55922 157276
rect 161566 157264 161572 157276
rect 55916 157236 161572 157264
rect 55916 157224 55922 157236
rect 161566 157224 161572 157236
rect 161624 157224 161630 157276
rect 202782 157264 202788 157276
rect 171106 157236 202788 157264
rect 45738 157156 45744 157208
rect 45796 157196 45802 157208
rect 153746 157196 153752 157208
rect 45796 157168 153752 157196
rect 45796 157156 45802 157168
rect 153746 157156 153752 157168
rect 153804 157156 153810 157208
rect 160094 157156 160100 157208
rect 160152 157196 160158 157208
rect 171106 157196 171134 157236
rect 202782 157224 202788 157236
rect 202840 157224 202846 157276
rect 203904 157264 203932 157304
rect 204898 157292 204904 157344
rect 204956 157332 204962 157344
rect 270494 157332 270500 157344
rect 204956 157304 270500 157332
rect 204956 157292 204962 157304
rect 270494 157292 270500 157304
rect 270552 157292 270558 157344
rect 204990 157264 204996 157276
rect 203904 157236 204996 157264
rect 204990 157224 204996 157236
rect 205048 157224 205054 157276
rect 205082 157224 205088 157276
rect 205140 157264 205146 157276
rect 273254 157264 273260 157276
rect 205140 157236 273260 157264
rect 205140 157224 205146 157236
rect 273254 157224 273260 157236
rect 273312 157224 273318 157276
rect 283834 157224 283840 157276
rect 283892 157264 283898 157276
rect 335538 157264 335544 157276
rect 283892 157236 335544 157264
rect 283892 157224 283898 157236
rect 335538 157224 335544 157236
rect 335596 157224 335602 157276
rect 160152 157168 171134 157196
rect 160152 157156 160158 157168
rect 192110 157156 192116 157208
rect 192168 157196 192174 157208
rect 265158 157196 265164 157208
rect 192168 157168 265164 157196
rect 192168 157156 192174 157168
rect 265158 157156 265164 157168
rect 265216 157156 265222 157208
rect 280430 157156 280436 157208
rect 280488 157196 280494 157208
rect 333054 157196 333060 157208
rect 280488 157168 333060 157196
rect 280488 157156 280494 157168
rect 333054 157156 333060 157168
rect 333112 157156 333118 157208
rect 39022 157088 39028 157140
rect 39080 157128 39086 157140
rect 147674 157128 147680 157140
rect 39080 157100 147680 157128
rect 39080 157088 39086 157100
rect 147674 157088 147680 157100
rect 147732 157088 147738 157140
rect 166902 157088 166908 157140
rect 166960 157128 166966 157140
rect 245838 157128 245844 157140
rect 166960 157100 245844 157128
rect 166960 157088 166966 157100
rect 245838 157088 245844 157100
rect 245896 157088 245902 157140
rect 273714 157088 273720 157140
rect 273772 157128 273778 157140
rect 327902 157128 327908 157140
rect 273772 157100 327908 157128
rect 273772 157088 273778 157100
rect 327902 157088 327908 157100
rect 327960 157088 327966 157140
rect 35710 157020 35716 157072
rect 35768 157060 35774 157072
rect 145466 157060 145472 157072
rect 35768 157032 145472 157060
rect 35768 157020 35774 157032
rect 145466 157020 145472 157032
rect 145524 157020 145530 157072
rect 146846 157020 146852 157072
rect 146904 157060 146910 157072
rect 150434 157060 150440 157072
rect 146904 157032 150440 157060
rect 146904 157020 146910 157032
rect 150434 157020 150440 157032
rect 150492 157020 150498 157072
rect 151722 157020 151728 157072
rect 151780 157060 151786 157072
rect 234798 157060 234804 157072
rect 151780 157032 234804 157060
rect 151780 157020 151786 157032
rect 234798 157020 234804 157032
rect 234856 157020 234862 157072
rect 277118 157020 277124 157072
rect 277176 157060 277182 157072
rect 330478 157060 330484 157072
rect 277176 157032 330484 157060
rect 277176 157020 277182 157032
rect 330478 157020 330484 157032
rect 330536 157020 330542 157072
rect 24762 156952 24768 157004
rect 24820 156992 24826 157004
rect 136910 156992 136916 157004
rect 24820 156964 136916 156992
rect 24820 156952 24826 156964
rect 136910 156952 136916 156964
rect 136968 156952 136974 157004
rect 138290 156952 138296 157004
rect 138348 156992 138354 157004
rect 224126 156992 224132 157004
rect 138348 156964 224132 156992
rect 138348 156952 138354 156964
rect 224126 156952 224132 156964
rect 224184 156952 224190 157004
rect 270310 156952 270316 157004
rect 270368 156992 270374 157004
rect 325326 156992 325332 157004
rect 270368 156964 325332 156992
rect 270368 156952 270374 156964
rect 325326 156952 325332 156964
rect 325384 156952 325390 157004
rect 18046 156884 18052 156936
rect 18104 156924 18110 156936
rect 132494 156924 132500 156936
rect 18104 156896 132500 156924
rect 18104 156884 18110 156896
rect 132494 156884 132500 156896
rect 132552 156884 132558 156936
rect 134886 156884 134892 156936
rect 134944 156924 134950 156936
rect 210510 156924 210516 156936
rect 134944 156896 210516 156924
rect 134944 156884 134950 156896
rect 210510 156884 210516 156896
rect 210568 156884 210574 156936
rect 210602 156884 210608 156936
rect 210660 156924 210666 156936
rect 222286 156924 222292 156936
rect 210660 156896 222292 156924
rect 210660 156884 210666 156896
rect 222286 156884 222292 156896
rect 222344 156884 222350 156936
rect 226610 156884 226616 156936
rect 226668 156924 226674 156936
rect 291930 156924 291936 156936
rect 226668 156896 291936 156924
rect 226668 156884 226674 156896
rect 291930 156884 291936 156896
rect 291988 156884 291994 156936
rect 293862 156884 293868 156936
rect 293920 156924 293926 156936
rect 342714 156924 342720 156936
rect 293920 156896 342720 156924
rect 293920 156884 293926 156896
rect 342714 156884 342720 156896
rect 342772 156884 342778 156936
rect 21358 156816 21364 156868
rect 21416 156856 21422 156868
rect 135254 156856 135260 156868
rect 21416 156828 135260 156856
rect 21416 156816 21422 156828
rect 135254 156816 135260 156828
rect 135312 156816 135318 156868
rect 139118 156816 139124 156868
rect 139176 156856 139182 156868
rect 225138 156856 225144 156868
rect 139176 156828 225144 156856
rect 139176 156816 139182 156828
rect 225138 156816 225144 156828
rect 225196 156816 225202 156868
rect 230014 156816 230020 156868
rect 230072 156856 230078 156868
rect 294046 156856 294052 156868
rect 230072 156828 294052 156856
rect 230072 156816 230078 156828
rect 294046 156816 294052 156828
rect 294104 156816 294110 156868
rect 297266 156816 297272 156868
rect 297324 156856 297330 156868
rect 345106 156856 345112 156868
rect 297324 156828 345112 156856
rect 297324 156816 297330 156828
rect 345106 156816 345112 156828
rect 345164 156816 345170 156868
rect 128170 156748 128176 156800
rect 128228 156788 128234 156800
rect 214098 156788 214104 156800
rect 128228 156760 214104 156788
rect 128228 156748 128234 156760
rect 214098 156748 214104 156760
rect 214156 156748 214162 156800
rect 214208 156760 215294 156788
rect 14642 156680 14648 156732
rect 14700 156720 14706 156732
rect 130102 156720 130108 156732
rect 14700 156692 130108 156720
rect 14700 156680 14706 156692
rect 130102 156680 130108 156692
rect 130160 156680 130166 156732
rect 132402 156680 132408 156732
rect 132460 156720 132466 156732
rect 214208 156720 214236 156760
rect 132460 156692 214236 156720
rect 215266 156720 215294 156760
rect 219894 156748 219900 156800
rect 219952 156788 219958 156800
rect 286318 156788 286324 156800
rect 219952 156760 286324 156788
rect 219952 156748 219958 156760
rect 286318 156748 286324 156760
rect 286376 156748 286382 156800
rect 287146 156748 287152 156800
rect 287204 156788 287210 156800
rect 338114 156788 338120 156800
rect 287204 156760 338120 156788
rect 287204 156748 287210 156760
rect 338114 156748 338120 156760
rect 338172 156748 338178 156800
rect 219986 156720 219992 156732
rect 215266 156692 219992 156720
rect 132460 156680 132466 156692
rect 219986 156680 219992 156692
rect 220044 156680 220050 156732
rect 223206 156680 223212 156732
rect 223264 156720 223270 156732
rect 289354 156720 289360 156732
rect 223264 156692 289360 156720
rect 223264 156680 223270 156692
rect 289354 156680 289360 156692
rect 289412 156680 289418 156732
rect 290550 156680 290556 156732
rect 290608 156720 290614 156732
rect 340690 156720 340696 156732
rect 290608 156692 340696 156720
rect 290608 156680 290614 156692
rect 340690 156680 340696 156692
rect 340748 156680 340754 156732
rect 344370 156680 344376 156732
rect 344428 156720 344434 156732
rect 381814 156720 381820 156732
rect 344428 156692 381820 156720
rect 344428 156680 344434 156692
rect 381814 156680 381820 156692
rect 381872 156680 381878 156732
rect 2038 156612 2044 156664
rect 2096 156652 2102 156664
rect 120442 156652 120448 156664
rect 2096 156624 120448 156652
rect 2096 156612 2102 156624
rect 120442 156612 120448 156624
rect 120500 156612 120506 156664
rect 124858 156612 124864 156664
rect 124916 156652 124922 156664
rect 209682 156652 209688 156664
rect 124916 156624 209688 156652
rect 124916 156612 124922 156624
rect 209682 156612 209688 156624
rect 209740 156612 209746 156664
rect 209774 156612 209780 156664
rect 209832 156652 209838 156664
rect 210694 156652 210700 156664
rect 209832 156624 210700 156652
rect 209832 156612 209838 156624
rect 210694 156612 210700 156624
rect 210752 156612 210758 156664
rect 210786 156612 210792 156664
rect 210844 156652 210850 156664
rect 214190 156652 214196 156664
rect 210844 156624 214196 156652
rect 210844 156612 210850 156624
rect 214190 156612 214196 156624
rect 214248 156612 214254 156664
rect 214282 156612 214288 156664
rect 214340 156652 214346 156664
rect 216398 156652 216404 156664
rect 214340 156624 216404 156652
rect 214340 156612 214346 156624
rect 216398 156612 216404 156624
rect 216456 156612 216462 156664
rect 216490 156612 216496 156664
rect 216548 156652 216554 156664
rect 283098 156652 283104 156664
rect 216548 156624 283104 156652
rect 216548 156612 216554 156624
rect 283098 156612 283104 156624
rect 283156 156612 283162 156664
rect 337654 156612 337660 156664
rect 337712 156652 337718 156664
rect 376662 156652 376668 156664
rect 337712 156624 376668 156652
rect 337712 156612 337718 156624
rect 376662 156612 376668 156624
rect 376720 156612 376726 156664
rect 498286 156612 498292 156664
rect 498344 156652 498350 156664
rect 499298 156652 499304 156664
rect 498344 156624 499304 156652
rect 498344 156612 498350 156624
rect 499298 156612 499304 156624
rect 499356 156612 499362 156664
rect 59262 156544 59268 156596
rect 59320 156584 59326 156596
rect 164142 156584 164148 156596
rect 59320 156556 164148 156584
rect 59320 156544 59326 156556
rect 164142 156544 164148 156556
rect 164200 156544 164206 156596
rect 164234 156544 164240 156596
rect 164292 156584 164298 156596
rect 228358 156584 228364 156596
rect 164292 156556 228364 156584
rect 164292 156544 164298 156556
rect 228358 156544 228364 156556
rect 228416 156544 228422 156596
rect 72694 156476 72700 156528
rect 72752 156516 72758 156528
rect 174446 156516 174452 156528
rect 72752 156488 174452 156516
rect 72752 156476 72758 156488
rect 174446 156476 174452 156488
rect 174504 156476 174510 156528
rect 174998 156476 175004 156528
rect 175056 156516 175062 156528
rect 175056 156488 195974 156516
rect 175056 156476 175062 156488
rect 79410 156408 79416 156460
rect 79468 156448 79474 156460
rect 179598 156448 179604 156460
rect 79468 156420 179604 156448
rect 79468 156408 79474 156420
rect 179598 156408 179604 156420
rect 179656 156408 179662 156460
rect 92842 156340 92848 156392
rect 92900 156380 92906 156392
rect 189810 156380 189816 156392
rect 92900 156352 189816 156380
rect 92900 156340 92906 156352
rect 189810 156340 189816 156352
rect 189868 156340 189874 156392
rect 195946 156380 195974 156488
rect 198826 156476 198832 156528
rect 198884 156516 198890 156528
rect 204898 156516 204904 156528
rect 198884 156488 204904 156516
rect 198884 156476 198890 156488
rect 204898 156476 204904 156488
rect 204956 156476 204962 156528
rect 204990 156476 204996 156528
rect 205048 156516 205054 156528
rect 210418 156516 210424 156528
rect 205048 156488 210424 156516
rect 205048 156476 205054 156488
rect 210418 156476 210424 156488
rect 210476 156476 210482 156528
rect 210510 156476 210516 156528
rect 210568 156516 210574 156528
rect 221366 156516 221372 156528
rect 210568 156488 221372 156516
rect 210568 156476 210574 156488
rect 221366 156476 221372 156488
rect 221424 156476 221430 156528
rect 223574 156476 223580 156528
rect 223632 156516 223638 156528
rect 281626 156516 281632 156528
rect 223632 156488 281632 156516
rect 223632 156476 223638 156488
rect 281626 156476 281632 156488
rect 281684 156476 281690 156528
rect 202690 156408 202696 156460
rect 202748 156448 202754 156460
rect 205082 156448 205088 156460
rect 202748 156420 205088 156448
rect 202748 156408 202754 156420
rect 205082 156408 205088 156420
rect 205140 156408 205146 156460
rect 210344 156420 210648 156448
rect 210344 156380 210372 156420
rect 195946 156352 210372 156380
rect 210620 156380 210648 156420
rect 210694 156408 210700 156460
rect 210752 156448 210758 156460
rect 279050 156448 279056 156460
rect 210752 156420 279056 156448
rect 210752 156408 210758 156420
rect 279050 156408 279056 156420
rect 279108 156408 279114 156460
rect 230934 156380 230940 156392
rect 210620 156352 230940 156380
rect 230934 156340 230940 156352
rect 230992 156340 230998 156392
rect 101306 156272 101312 156324
rect 101364 156312 101370 156324
rect 196250 156312 196256 156324
rect 101364 156284 196256 156312
rect 101364 156272 101370 156284
rect 196250 156272 196256 156284
rect 196308 156272 196314 156324
rect 202782 156272 202788 156324
rect 202840 156312 202846 156324
rect 202840 156284 210372 156312
rect 202840 156272 202846 156284
rect 108022 156204 108028 156256
rect 108080 156244 108086 156256
rect 200298 156244 200304 156256
rect 108080 156216 200304 156244
rect 108080 156204 108086 156216
rect 200298 156204 200304 156216
rect 200356 156204 200362 156256
rect 205910 156204 205916 156256
rect 205968 156244 205974 156256
rect 210344 156244 210372 156284
rect 210418 156272 210424 156324
rect 210476 156312 210482 156324
rect 219526 156312 219532 156324
rect 210476 156284 219532 156312
rect 210476 156272 210482 156284
rect 219526 156272 219532 156284
rect 219584 156272 219590 156324
rect 222102 156272 222108 156324
rect 222160 156312 222166 156324
rect 269482 156312 269488 156324
rect 222160 156284 269488 156312
rect 222160 156272 222166 156284
rect 269482 156272 269488 156284
rect 269540 156272 269546 156324
rect 210602 156244 210608 156256
rect 205968 156216 210280 156244
rect 210344 156216 210608 156244
rect 205968 156204 205974 156216
rect 118142 156136 118148 156188
rect 118200 156176 118206 156188
rect 203886 156176 203892 156188
rect 118200 156148 203892 156176
rect 118200 156136 118206 156148
rect 203886 156136 203892 156148
rect 203944 156136 203950 156188
rect 210252 156176 210280 156216
rect 210602 156204 210608 156216
rect 210660 156204 210666 156256
rect 213178 156204 213184 156256
rect 213236 156244 213242 156256
rect 223574 156244 223580 156256
rect 213236 156216 223580 156244
rect 213236 156204 213242 156216
rect 223574 156204 223580 156216
rect 223632 156204 223638 156256
rect 266906 156244 266912 156256
rect 224052 156216 266912 156244
rect 211614 156176 211620 156188
rect 210252 156148 211620 156176
rect 211614 156136 211620 156148
rect 211672 156136 211678 156188
rect 220630 156136 220636 156188
rect 220688 156176 220694 156188
rect 224052 156176 224080 156216
rect 266906 156204 266912 156216
rect 266964 156204 266970 156256
rect 220688 156148 224080 156176
rect 220688 156136 220694 156148
rect 227714 156136 227720 156188
rect 227772 156176 227778 156188
rect 272058 156176 272064 156188
rect 227772 156148 272064 156176
rect 227772 156136 227778 156148
rect 272058 156136 272064 156148
rect 272116 156136 272122 156188
rect 121454 156068 121460 156120
rect 121512 156108 121518 156120
rect 205726 156108 205732 156120
rect 121512 156080 205732 156108
rect 121512 156068 121518 156080
rect 205726 156068 205732 156080
rect 205784 156068 205790 156120
rect 211062 156068 211068 156120
rect 211120 156108 211126 156120
rect 273898 156108 273904 156120
rect 211120 156080 273904 156108
rect 211120 156068 211126 156080
rect 273898 156068 273904 156080
rect 273956 156068 273962 156120
rect 11238 156000 11244 156052
rect 11296 156040 11302 156052
rect 127526 156040 127532 156052
rect 11296 156012 127532 156040
rect 11296 156000 11302 156012
rect 127526 156000 127532 156012
rect 127584 156000 127590 156052
rect 135806 156000 135812 156052
rect 135864 156040 135870 156052
rect 222562 156040 222568 156052
rect 135864 156012 222568 156040
rect 135864 156000 135870 156012
rect 222562 156000 222568 156012
rect 222620 156000 222626 156052
rect 145006 155932 145012 155984
rect 145064 155972 145070 155984
rect 229646 155972 229652 155984
rect 145064 155944 229652 155972
rect 145064 155932 145070 155944
rect 229646 155932 229652 155944
rect 229704 155932 229710 155984
rect 60090 155864 60096 155916
rect 60148 155904 60154 155916
rect 84746 155904 84752 155916
rect 60148 155876 84752 155904
rect 60148 155864 60154 155876
rect 84746 155864 84752 155876
rect 84804 155864 84810 155916
rect 88702 155864 88708 155916
rect 88760 155904 88766 155916
rect 186774 155904 186780 155916
rect 88760 155876 186780 155904
rect 88760 155864 88766 155876
rect 186774 155864 186780 155876
rect 186832 155864 186838 155916
rect 189626 155864 189632 155916
rect 189684 155904 189690 155916
rect 263778 155904 263784 155916
rect 189684 155876 263784 155904
rect 189684 155864 189690 155876
rect 263778 155864 263784 155876
rect 263836 155864 263842 155916
rect 299750 155864 299756 155916
rect 299808 155904 299814 155916
rect 347866 155904 347872 155916
rect 299808 155876 347872 155904
rect 299808 155864 299814 155876
rect 347866 155864 347872 155876
rect 347924 155864 347930 155916
rect 12158 155796 12164 155848
rect 12216 155836 12222 155848
rect 109034 155836 109040 155848
rect 12216 155808 109040 155836
rect 12216 155796 12222 155808
rect 109034 155796 109040 155808
rect 109092 155796 109098 155848
rect 112254 155796 112260 155848
rect 112312 155836 112318 155848
rect 204346 155836 204352 155848
rect 112312 155808 204352 155836
rect 112312 155796 112318 155808
rect 204346 155796 204352 155808
rect 204404 155796 204410 155848
rect 206462 155796 206468 155848
rect 206520 155836 206526 155848
rect 276106 155836 276112 155848
rect 206520 155808 276112 155836
rect 206520 155796 206526 155808
rect 276106 155796 276112 155808
rect 276164 155796 276170 155848
rect 296438 155796 296444 155848
rect 296496 155836 296502 155848
rect 345198 155836 345204 155848
rect 296496 155808 345204 155836
rect 296496 155796 296502 155808
rect 345198 155796 345204 155808
rect 345256 155796 345262 155848
rect 46566 155728 46572 155780
rect 46624 155768 46630 155780
rect 75822 155768 75828 155780
rect 46624 155740 75828 155768
rect 46624 155728 46630 155740
rect 75822 155728 75828 155740
rect 75880 155728 75886 155780
rect 81894 155728 81900 155780
rect 81952 155768 81958 155780
rect 181438 155768 181444 155780
rect 81952 155740 181444 155768
rect 81952 155728 81958 155740
rect 181438 155728 181444 155740
rect 181496 155728 181502 155780
rect 186222 155728 186228 155780
rect 186280 155768 186286 155780
rect 260834 155768 260840 155780
rect 186280 155740 260840 155768
rect 186280 155728 186286 155740
rect 260834 155728 260840 155740
rect 260892 155728 260898 155780
rect 293034 155728 293040 155780
rect 293092 155768 293098 155780
rect 342346 155768 342352 155780
rect 293092 155740 342352 155768
rect 293092 155728 293098 155740
rect 342346 155728 342352 155740
rect 342404 155728 342410 155780
rect 71866 155660 71872 155712
rect 71924 155700 71930 155712
rect 172698 155700 172704 155712
rect 71924 155672 172704 155700
rect 71924 155660 71930 155672
rect 172698 155660 172704 155672
rect 172756 155660 172762 155712
rect 176286 155660 176292 155712
rect 176344 155700 176350 155712
rect 253382 155700 253388 155712
rect 176344 155672 253388 155700
rect 176344 155660 176350 155672
rect 253382 155660 253388 155672
rect 253440 155660 253446 155712
rect 289722 155660 289728 155712
rect 289780 155700 289786 155712
rect 340046 155700 340052 155712
rect 289780 155672 340052 155700
rect 289780 155660 289786 155672
rect 340046 155660 340052 155672
rect 340104 155660 340110 155712
rect 33134 155592 33140 155644
rect 33192 155632 33198 155644
rect 59998 155632 60004 155644
rect 33192 155604 60004 155632
rect 33192 155592 33198 155604
rect 59998 155592 60004 155604
rect 60056 155592 60062 155644
rect 75178 155592 75184 155644
rect 75236 155632 75242 155644
rect 176378 155632 176384 155644
rect 75236 155604 176384 155632
rect 75236 155592 75242 155604
rect 176378 155592 176384 155604
rect 176436 155592 176442 155644
rect 177114 155592 177120 155644
rect 177172 155632 177178 155644
rect 254026 155632 254032 155644
rect 177172 155604 254032 155632
rect 177172 155592 177178 155604
rect 254026 155592 254032 155604
rect 254084 155592 254090 155644
rect 266998 155592 267004 155644
rect 267056 155632 267062 155644
rect 321738 155632 321744 155644
rect 267056 155604 321744 155632
rect 267056 155592 267062 155604
rect 321738 155592 321744 155604
rect 321796 155592 321802 155644
rect 39850 155524 39856 155576
rect 39908 155564 39914 155576
rect 71774 155564 71780 155576
rect 39908 155536 71780 155564
rect 39908 155524 39914 155536
rect 71774 155524 71780 155536
rect 71832 155524 71838 155576
rect 78582 155524 78588 155576
rect 78640 155564 78646 155576
rect 178954 155564 178960 155576
rect 78640 155536 178960 155564
rect 78640 155524 78646 155536
rect 178954 155524 178960 155536
rect 179012 155524 179018 155576
rect 179506 155524 179512 155576
rect 179564 155564 179570 155576
rect 255866 155564 255872 155576
rect 179564 155536 255872 155564
rect 179564 155524 179570 155536
rect 255866 155524 255872 155536
rect 255924 155524 255930 155576
rect 263594 155524 263600 155576
rect 263652 155564 263658 155576
rect 320174 155564 320180 155576
rect 263652 155536 320180 155564
rect 263652 155524 263658 155536
rect 320174 155524 320180 155536
rect 320232 155524 320238 155576
rect 340966 155524 340972 155576
rect 341024 155564 341030 155576
rect 378134 155564 378140 155576
rect 341024 155536 378140 155564
rect 341024 155524 341030 155536
rect 378134 155524 378140 155536
rect 378192 155524 378198 155576
rect 28902 155456 28908 155508
rect 28960 155496 28966 155508
rect 56502 155496 56508 155508
rect 28960 155468 56508 155496
rect 28960 155456 28966 155468
rect 56502 155456 56508 155468
rect 56560 155456 56566 155508
rect 62574 155456 62580 155508
rect 62632 155496 62638 155508
rect 165706 155496 165712 155508
rect 62632 155468 165712 155496
rect 62632 155456 62638 155468
rect 165706 155456 165712 155468
rect 165764 155456 165770 155508
rect 169386 155456 169392 155508
rect 169444 155496 169450 155508
rect 248230 155496 248236 155508
rect 169444 155468 248236 155496
rect 169444 155456 169450 155468
rect 248230 155456 248236 155468
rect 248288 155456 248294 155508
rect 260282 155456 260288 155508
rect 260340 155496 260346 155508
rect 317598 155496 317604 155508
rect 260340 155468 317604 155496
rect 260340 155456 260346 155468
rect 317598 155456 317604 155468
rect 317656 155456 317662 155508
rect 333422 155456 333428 155508
rect 333480 155496 333486 155508
rect 373442 155496 373448 155508
rect 333480 155468 373448 155496
rect 333480 155456 333486 155468
rect 373442 155456 373448 155468
rect 373500 155456 373506 155508
rect 7926 155388 7932 155440
rect 7984 155428 7990 155440
rect 124674 155428 124680 155440
rect 7984 155400 124680 155428
rect 7984 155388 7990 155400
rect 124674 155388 124680 155400
rect 124732 155388 124738 155440
rect 134058 155388 134064 155440
rect 134116 155428 134122 155440
rect 137554 155428 137560 155440
rect 134116 155400 137560 155428
rect 134116 155388 134122 155400
rect 137554 155388 137560 155400
rect 137612 155388 137618 155440
rect 149238 155388 149244 155440
rect 149296 155428 149302 155440
rect 232866 155428 232872 155440
rect 149296 155400 232872 155428
rect 149296 155388 149302 155400
rect 232866 155388 232872 155400
rect 232924 155388 232930 155440
rect 253566 155388 253572 155440
rect 253624 155428 253630 155440
rect 312446 155428 312452 155440
rect 253624 155400 312452 155428
rect 253624 155388 253630 155400
rect 312446 155388 312452 155400
rect 312504 155388 312510 155440
rect 330110 155388 330116 155440
rect 330168 155428 330174 155440
rect 370866 155428 370872 155440
rect 330168 155400 370872 155428
rect 330168 155388 330174 155400
rect 370866 155388 370872 155400
rect 370924 155388 370930 155440
rect 8754 155320 8760 155372
rect 8812 155360 8818 155372
rect 125686 155360 125692 155372
rect 8812 155332 125692 155360
rect 8812 155320 8818 155332
rect 125686 155320 125692 155332
rect 125744 155320 125750 155372
rect 145834 155320 145840 155372
rect 145892 155360 145898 155372
rect 229186 155360 229192 155372
rect 145892 155332 229192 155360
rect 145892 155320 145898 155332
rect 229186 155320 229192 155332
rect 229244 155320 229250 155372
rect 250162 155320 250168 155372
rect 250220 155360 250226 155372
rect 309870 155360 309876 155372
rect 250220 155332 309876 155360
rect 250220 155320 250226 155332
rect 309870 155320 309876 155332
rect 309928 155320 309934 155372
rect 316586 155320 316592 155372
rect 316644 155360 316650 155372
rect 360654 155360 360660 155372
rect 316644 155332 360660 155360
rect 316644 155320 316650 155332
rect 360654 155320 360660 155332
rect 360712 155320 360718 155372
rect 4522 155252 4528 155304
rect 4580 155292 4586 155304
rect 122006 155292 122012 155304
rect 4580 155264 122012 155292
rect 4580 155252 4586 155264
rect 122006 155252 122012 155264
rect 122064 155252 122070 155304
rect 142522 155252 142528 155304
rect 142580 155292 142586 155304
rect 227806 155292 227812 155304
rect 142580 155264 227812 155292
rect 142580 155252 142586 155264
rect 227806 155252 227812 155264
rect 227864 155252 227870 155304
rect 243446 155252 243452 155304
rect 243504 155292 243510 155304
rect 304718 155292 304724 155304
rect 243504 155264 304724 155292
rect 243504 155252 243510 155264
rect 304718 155252 304724 155264
rect 304776 155252 304782 155304
rect 306558 155252 306564 155304
rect 306616 155292 306622 155304
rect 352466 155292 352472 155304
rect 306616 155264 352472 155292
rect 306616 155252 306622 155264
rect 352466 155252 352472 155264
rect 352524 155252 352530 155304
rect 373810 155252 373816 155304
rect 373868 155292 373874 155304
rect 403158 155292 403164 155304
rect 373868 155264 403164 155292
rect 373868 155252 373874 155264
rect 403158 155252 403164 155264
rect 403216 155252 403222 155304
rect 5350 155184 5356 155236
rect 5408 155224 5414 155236
rect 123018 155224 123024 155236
rect 5408 155196 123024 155224
rect 5408 155184 5414 155196
rect 123018 155184 123024 155196
rect 123076 155184 123082 155236
rect 128998 155184 129004 155236
rect 129056 155224 129062 155236
rect 217410 155224 217416 155236
rect 129056 155196 217416 155224
rect 129056 155184 129062 155196
rect 217410 155184 217416 155196
rect 217468 155184 217474 155236
rect 236730 155184 236736 155236
rect 236788 155224 236794 155236
rect 299658 155224 299664 155236
rect 236788 155196 299664 155224
rect 236788 155184 236794 155196
rect 299658 155184 299664 155196
rect 299716 155184 299722 155236
rect 303154 155184 303160 155236
rect 303212 155224 303218 155236
rect 350350 155224 350356 155236
rect 303212 155196 350356 155224
rect 303212 155184 303218 155196
rect 350350 155184 350356 155196
rect 350408 155184 350414 155236
rect 367094 155184 367100 155236
rect 367152 155224 367158 155236
rect 399018 155224 399024 155236
rect 367152 155196 399024 155224
rect 367152 155184 367158 155196
rect 399018 155184 399024 155196
rect 399076 155184 399082 155236
rect 401594 155184 401600 155236
rect 401652 155224 401658 155236
rect 425514 155224 425520 155236
rect 401652 155196 425520 155224
rect 401652 155184 401658 155196
rect 425514 155184 425520 155196
rect 425572 155184 425578 155236
rect 53374 155116 53380 155168
rect 53432 155156 53438 155168
rect 76926 155156 76932 155168
rect 53432 155128 76932 155156
rect 53432 155116 53438 155128
rect 76926 155116 76932 155128
rect 76984 155116 76990 155168
rect 86126 155116 86132 155168
rect 86184 155156 86190 155168
rect 183554 155156 183560 155168
rect 86184 155128 183560 155156
rect 86184 155116 86190 155128
rect 183554 155116 183560 155128
rect 183612 155116 183618 155168
rect 186682 155116 186688 155168
rect 186740 155156 186746 155168
rect 186740 155128 192892 155156
rect 186740 155116 186746 155128
rect 95418 155048 95424 155100
rect 95476 155088 95482 155100
rect 186314 155088 186320 155100
rect 95476 155060 186320 155088
rect 95476 155048 95482 155060
rect 186314 155048 186320 155060
rect 186372 155048 186378 155100
rect 186498 155048 186504 155100
rect 186556 155088 186562 155100
rect 191742 155088 191748 155100
rect 186556 155060 191748 155088
rect 186556 155048 186562 155060
rect 191742 155048 191748 155060
rect 191800 155048 191806 155100
rect 192864 155088 192892 155128
rect 192938 155116 192944 155168
rect 192996 155156 193002 155168
rect 266262 155156 266268 155168
rect 192996 155128 266268 155156
rect 192996 155116 193002 155128
rect 266262 155116 266268 155128
rect 266320 155116 266326 155168
rect 309962 155116 309968 155168
rect 310020 155156 310026 155168
rect 355502 155156 355508 155168
rect 310020 155128 355508 155156
rect 310020 155116 310026 155128
rect 355502 155116 355508 155128
rect 355560 155116 355566 155168
rect 194962 155088 194968 155100
rect 192864 155060 194968 155088
rect 194962 155048 194968 155060
rect 195020 155048 195026 155100
rect 196342 155048 196348 155100
rect 196400 155088 196406 155100
rect 268838 155088 268844 155100
rect 196400 155060 268844 155088
rect 196400 155048 196406 155060
rect 268838 155048 268844 155060
rect 268896 155048 268902 155100
rect 98730 154980 98736 155032
rect 98788 155020 98794 155032
rect 186222 155020 186228 155032
rect 98788 154992 186228 155020
rect 98788 154980 98794 154992
rect 186222 154980 186228 154992
rect 186280 154980 186286 155032
rect 186590 154980 186596 155032
rect 186648 155020 186654 155032
rect 194318 155020 194324 155032
rect 186648 154992 194324 155020
rect 186648 154980 186654 154992
rect 194318 154980 194324 154992
rect 194376 154980 194382 155032
rect 199654 154980 199660 155032
rect 199712 155020 199718 155032
rect 271414 155020 271420 155032
rect 199712 154992 271420 155020
rect 199712 154980 199718 154992
rect 271414 154980 271420 154992
rect 271472 154980 271478 155032
rect 99558 154912 99564 154964
rect 99616 154952 99622 154964
rect 186314 154952 186320 154964
rect 99616 154924 186320 154952
rect 99616 154912 99622 154924
rect 186314 154912 186320 154924
rect 186372 154912 186378 154964
rect 188246 154912 188252 154964
rect 188304 154952 188310 154964
rect 240686 154952 240692 154964
rect 188304 154924 240692 154952
rect 188304 154912 188310 154924
rect 240686 154912 240692 154924
rect 240744 154912 240750 154964
rect 80238 154844 80244 154896
rect 80296 154884 80302 154896
rect 86862 154884 86868 154896
rect 80296 154856 86868 154884
rect 80296 154844 80302 154856
rect 86862 154844 86868 154856
rect 86920 154844 86926 154896
rect 122282 154844 122288 154896
rect 122340 154884 122346 154896
rect 212258 154884 212264 154896
rect 122340 154856 212264 154884
rect 122340 154844 122346 154856
rect 212258 154844 212264 154856
rect 212316 154844 212322 154896
rect 231762 154844 231768 154896
rect 231820 154884 231826 154896
rect 277118 154884 277124 154896
rect 231820 154856 277124 154884
rect 231820 154844 231826 154856
rect 277118 154844 277124 154856
rect 277176 154844 277182 154896
rect 125778 154776 125784 154828
rect 125836 154816 125842 154828
rect 214834 154816 214840 154828
rect 125836 154788 214840 154816
rect 125836 154776 125842 154788
rect 214834 154776 214840 154788
rect 214892 154776 214898 154828
rect 216766 154776 216772 154828
rect 216824 154816 216830 154828
rect 261386 154816 261392 154828
rect 216824 154788 261392 154816
rect 216824 154776 216830 154788
rect 261386 154776 261392 154788
rect 261444 154776 261450 154828
rect 107286 154708 107292 154760
rect 107344 154748 107350 154760
rect 133322 154748 133328 154760
rect 107344 154720 133328 154748
rect 107344 154708 107350 154720
rect 133322 154708 133328 154720
rect 133380 154708 133386 154760
rect 155954 154708 155960 154760
rect 156012 154748 156018 154760
rect 238018 154748 238024 154760
rect 156012 154720 238024 154748
rect 156012 154708 156018 154720
rect 238018 154708 238024 154720
rect 238076 154708 238082 154760
rect 110506 154640 110512 154692
rect 110564 154680 110570 154692
rect 128354 154680 128360 154692
rect 110564 154652 128360 154680
rect 110564 154640 110570 154652
rect 128354 154640 128360 154652
rect 128412 154640 128418 154692
rect 162670 154640 162676 154692
rect 162728 154680 162734 154692
rect 243078 154680 243084 154692
rect 162728 154652 243084 154680
rect 162728 154640 162734 154652
rect 243078 154640 243084 154652
rect 243136 154640 243142 154692
rect 146202 154572 146208 154624
rect 146260 154612 146266 154624
rect 146260 154584 150756 154612
rect 146260 154572 146266 154584
rect 44174 154504 44180 154556
rect 44232 154544 44238 154556
rect 146478 154544 146484 154556
rect 44232 154516 146484 154544
rect 44232 154504 44238 154516
rect 146478 154504 146484 154516
rect 146536 154504 146542 154556
rect 150618 154544 150624 154556
rect 146680 154516 150624 154544
rect 41598 154436 41604 154488
rect 41656 154476 41662 154488
rect 146680 154476 146708 154516
rect 150618 154504 150624 154516
rect 150676 154504 150682 154556
rect 150728 154544 150756 154584
rect 151814 154572 151820 154624
rect 151872 154612 151878 154624
rect 151872 154584 156736 154612
rect 151872 154572 151878 154584
rect 156598 154544 156604 154556
rect 150728 154516 156604 154544
rect 156598 154504 156604 154516
rect 156656 154504 156662 154556
rect 156708 154544 156736 154584
rect 159358 154572 159364 154624
rect 159416 154612 159422 154624
rect 240134 154612 240140 154624
rect 159416 154584 240140 154612
rect 159416 154572 159422 154584
rect 240134 154572 240140 154584
rect 240192 154572 240198 154624
rect 156782 154544 156788 154556
rect 156708 154516 156788 154544
rect 156782 154504 156788 154516
rect 156840 154504 156846 154556
rect 157334 154504 157340 154556
rect 157392 154544 157398 154556
rect 225782 154544 225788 154556
rect 157392 154516 225788 154544
rect 157392 154504 157398 154516
rect 225782 154504 225788 154516
rect 225840 154504 225846 154556
rect 231854 154504 231860 154556
rect 231912 154544 231918 154556
rect 296438 154544 296444 154556
rect 231912 154516 296444 154544
rect 231912 154504 231918 154516
rect 296438 154504 296444 154516
rect 296496 154504 296502 154556
rect 353662 154504 353668 154556
rect 353720 154544 353726 154556
rect 388898 154544 388904 154556
rect 353720 154516 388904 154544
rect 353720 154504 353726 154516
rect 388898 154504 388904 154516
rect 388956 154504 388962 154556
rect 185118 154476 185124 154488
rect 41656 154448 146708 154476
rect 146772 154448 185124 154476
rect 41656 154436 41662 154448
rect 34514 154368 34520 154420
rect 34572 154408 34578 154420
rect 145374 154408 145380 154420
rect 34572 154380 145380 154408
rect 34572 154368 34578 154380
rect 145374 154368 145380 154380
rect 145432 154368 145438 154420
rect 37918 154300 37924 154352
rect 37976 154340 37982 154352
rect 145098 154340 145104 154352
rect 37976 154312 145104 154340
rect 37976 154300 37982 154312
rect 145098 154300 145104 154312
rect 145156 154300 145162 154352
rect 30374 154232 30380 154284
rect 30432 154272 30438 154284
rect 137094 154272 137100 154284
rect 30432 154244 137100 154272
rect 30432 154232 30438 154244
rect 137094 154232 137100 154244
rect 137152 154232 137158 154284
rect 146772 154272 146800 154448
rect 185118 154436 185124 154448
rect 185176 154436 185182 154488
rect 191282 154436 191288 154488
rect 191340 154476 191346 154488
rect 200114 154476 200120 154488
rect 191340 154448 200120 154476
rect 191340 154436 191346 154448
rect 200114 154436 200120 154448
rect 200172 154436 200178 154488
rect 218330 154436 218336 154488
rect 218388 154476 218394 154488
rect 285582 154476 285588 154488
rect 218388 154448 285588 154476
rect 218388 154436 218394 154448
rect 285582 154436 285588 154448
rect 285640 154436 285646 154488
rect 285674 154436 285680 154488
rect 285732 154476 285738 154488
rect 337470 154476 337476 154488
rect 285732 154448 337476 154476
rect 285732 154436 285738 154448
rect 337470 154436 337476 154448
rect 337528 154436 337534 154488
rect 356238 154436 356244 154488
rect 356296 154476 356302 154488
rect 391474 154476 391480 154488
rect 356296 154448 391480 154476
rect 356296 154436 356302 154448
rect 391474 154436 391480 154448
rect 391532 154436 391538 154488
rect 400306 154436 400312 154488
rect 400364 154476 400370 154488
rect 424870 154476 424876 154488
rect 400364 154448 424876 154476
rect 400364 154436 400370 154448
rect 424870 154436 424876 154448
rect 424928 154436 424934 154488
rect 188430 154408 188436 154420
rect 137204 154244 146800 154272
rect 146864 154380 188436 154408
rect 23474 154164 23480 154216
rect 23532 154204 23538 154216
rect 137002 154204 137008 154216
rect 23532 154176 137008 154204
rect 23532 154164 23538 154176
rect 137002 154164 137008 154176
rect 137060 154164 137066 154216
rect 13814 154096 13820 154148
rect 13872 154136 13878 154148
rect 126790 154136 126796 154148
rect 13872 154108 126796 154136
rect 13872 154096 13878 154108
rect 126790 154096 126796 154108
rect 126848 154096 126854 154148
rect 137204 154136 137232 154244
rect 146864 154204 146892 154380
rect 188430 154368 188436 154380
rect 188488 154368 188494 154420
rect 191466 154368 191472 154420
rect 191524 154408 191530 154420
rect 202690 154408 202696 154420
rect 191524 154380 202696 154408
rect 191524 154368 191530 154380
rect 202690 154368 202696 154380
rect 202748 154368 202754 154420
rect 208394 154368 208400 154420
rect 208452 154408 208458 154420
rect 278406 154408 278412 154420
rect 208452 154380 278412 154408
rect 208452 154368 208458 154380
rect 278406 154368 278412 154380
rect 278464 154368 278470 154420
rect 278866 154368 278872 154420
rect 278924 154408 278930 154420
rect 332410 154408 332416 154420
rect 278924 154380 332416 154408
rect 278924 154368 278930 154380
rect 332410 154368 332416 154380
rect 332468 154368 332474 154420
rect 349522 154368 349528 154420
rect 349580 154408 349586 154420
rect 386322 154408 386328 154420
rect 349580 154380 386328 154408
rect 349580 154368 349586 154380
rect 386322 154368 386328 154380
rect 386380 154368 386386 154420
rect 397454 154368 397460 154420
rect 397512 154408 397518 154420
rect 423030 154408 423036 154420
rect 397512 154380 423036 154408
rect 397512 154368 397518 154380
rect 423030 154368 423036 154380
rect 423088 154368 423094 154420
rect 146938 154300 146944 154352
rect 146996 154340 147002 154352
rect 191282 154340 191288 154352
rect 146996 154312 191288 154340
rect 146996 154300 147002 154312
rect 191282 154300 191288 154312
rect 191340 154300 191346 154352
rect 191374 154300 191380 154352
rect 191432 154340 191438 154352
rect 202046 154340 202052 154352
rect 191432 154312 202052 154340
rect 191432 154300 191438 154312
rect 202046 154300 202052 154312
rect 202104 154300 202110 154352
rect 204806 154300 204812 154352
rect 204864 154340 204870 154352
rect 275830 154340 275836 154352
rect 204864 154312 275836 154340
rect 204864 154300 204870 154312
rect 275830 154300 275836 154312
rect 275888 154300 275894 154352
rect 276198 154300 276204 154352
rect 276256 154340 276262 154352
rect 329926 154340 329932 154352
rect 276256 154312 329932 154340
rect 276256 154300 276262 154312
rect 329926 154300 329932 154312
rect 329984 154300 329990 154352
rect 346394 154300 346400 154352
rect 346452 154340 346458 154352
rect 383746 154340 383752 154352
rect 346452 154312 383752 154340
rect 346452 154300 346458 154312
rect 383746 154300 383752 154312
rect 383804 154300 383810 154352
rect 390646 154300 390652 154352
rect 390704 154340 390710 154352
rect 417142 154340 417148 154352
rect 390704 154312 417148 154340
rect 390704 154300 390710 154312
rect 417142 154300 417148 154312
rect 417200 154300 417206 154352
rect 185210 154272 185216 154284
rect 127084 154108 137232 154136
rect 137296 154176 146892 154204
rect 146956 154244 185216 154272
rect 9674 154028 9680 154080
rect 9732 154068 9738 154080
rect 126882 154068 126888 154080
rect 9732 154040 126888 154068
rect 9732 154028 9738 154040
rect 126882 154028 126888 154040
rect 126940 154028 126946 154080
rect 127084 154068 127112 154108
rect 137296 154068 137324 154176
rect 146846 154136 146852 154148
rect 126992 154040 127112 154068
rect 127728 154040 137324 154068
rect 137388 154108 146852 154136
rect 7098 153960 7104 154012
rect 7156 154000 7162 154012
rect 117958 154000 117964 154012
rect 7156 153972 117964 154000
rect 7156 153960 7162 153972
rect 117958 153960 117964 153972
rect 118016 153960 118022 154012
rect 121730 154000 121736 154012
rect 118068 153972 121736 154000
rect 2958 153892 2964 153944
rect 3016 153932 3022 153944
rect 118068 153932 118096 153972
rect 121730 153960 121736 153972
rect 121788 153960 121794 154012
rect 121822 153960 121828 154012
rect 121880 154000 121886 154012
rect 126992 154000 127020 154040
rect 127728 154000 127756 154040
rect 121880 153972 127020 154000
rect 127084 153972 127756 154000
rect 121880 153960 121886 153972
rect 3016 153904 118096 153932
rect 3016 153892 3022 153904
rect 118142 153892 118148 153944
rect 118200 153932 118206 153944
rect 124306 153932 124312 153944
rect 118200 153904 124312 153932
rect 118200 153892 118206 153904
rect 124306 153892 124312 153904
rect 124364 153892 124370 153944
rect 125502 153892 125508 153944
rect 125560 153932 125566 153944
rect 127084 153932 127112 153972
rect 127894 153960 127900 154012
rect 127952 154000 127958 154012
rect 137388 154000 137416 154108
rect 146846 154096 146852 154108
rect 146904 154096 146910 154148
rect 137462 154028 137468 154080
rect 137520 154068 137526 154080
rect 137520 154040 137600 154068
rect 137520 154028 137526 154040
rect 127952 153972 137416 154000
rect 137572 154000 137600 154040
rect 137646 154028 137652 154080
rect 137704 154068 137710 154080
rect 146956 154068 146984 154244
rect 185210 154232 185216 154244
rect 185268 154232 185274 154284
rect 185302 154232 185308 154284
rect 185360 154272 185366 154284
rect 258534 154272 258540 154284
rect 185360 154244 258540 154272
rect 185360 154232 185366 154244
rect 258534 154232 258540 154244
rect 258592 154232 258598 154284
rect 262214 154232 262220 154284
rect 262272 154272 262278 154284
rect 319530 154272 319536 154284
rect 262272 154244 319536 154272
rect 262272 154232 262278 154244
rect 319530 154232 319536 154244
rect 319588 154232 319594 154284
rect 336826 154232 336832 154284
rect 336884 154272 336890 154284
rect 376018 154272 376024 154284
rect 336884 154244 376024 154272
rect 336884 154232 336890 154244
rect 376018 154232 376024 154244
rect 376076 154232 376082 154284
rect 393314 154232 393320 154284
rect 393372 154272 393378 154284
rect 419718 154272 419724 154284
rect 393372 154244 419724 154272
rect 393372 154232 393378 154244
rect 419718 154232 419724 154244
rect 419776 154232 419782 154284
rect 147122 154164 147128 154216
rect 147180 154204 147186 154216
rect 152734 154204 152740 154216
rect 147180 154176 152740 154204
rect 147180 154164 147186 154176
rect 152734 154164 152740 154176
rect 152792 154164 152798 154216
rect 153286 154164 153292 154216
rect 153344 154204 153350 154216
rect 163498 154204 163504 154216
rect 153344 154176 163504 154204
rect 153344 154164 153350 154176
rect 163498 154164 163504 154176
rect 163556 154164 163562 154216
rect 165062 154164 165068 154216
rect 165120 154204 165126 154216
rect 168650 154204 168656 154216
rect 165120 154176 168656 154204
rect 165120 154164 165126 154176
rect 168650 154164 168656 154176
rect 168708 154164 168714 154216
rect 172514 154164 172520 154216
rect 172572 154204 172578 154216
rect 250806 154204 250812 154216
rect 172572 154176 250812 154204
rect 172572 154164 172578 154176
rect 250806 154164 250812 154176
rect 250864 154164 250870 154216
rect 255314 154164 255320 154216
rect 255372 154204 255378 154216
rect 314378 154204 314384 154216
rect 255372 154176 314384 154204
rect 255372 154164 255378 154176
rect 314378 154164 314384 154176
rect 314436 154164 314442 154216
rect 342806 154164 342812 154216
rect 342864 154204 342870 154216
rect 381170 154204 381176 154216
rect 342864 154176 381176 154204
rect 342864 154164 342870 154176
rect 381170 154164 381176 154176
rect 381228 154164 381234 154216
rect 386506 154164 386512 154216
rect 386564 154204 386570 154216
rect 414566 154204 414572 154216
rect 386564 154176 414572 154204
rect 386564 154164 386570 154176
rect 414566 154164 414572 154176
rect 414624 154164 414630 154216
rect 147030 154096 147036 154148
rect 147088 154136 147094 154148
rect 147088 154108 148272 154136
rect 147088 154096 147094 154108
rect 148134 154068 148140 154080
rect 137704 154040 146984 154068
rect 147048 154040 148140 154068
rect 137704 154028 137710 154040
rect 142338 154000 142344 154012
rect 137572 153972 142344 154000
rect 127952 153960 127958 153972
rect 142338 153960 142344 153972
rect 142396 153960 142402 154012
rect 145098 153960 145104 154012
rect 145156 154000 145162 154012
rect 147048 154000 147076 154040
rect 148134 154028 148140 154040
rect 148192 154028 148198 154080
rect 145156 153972 147076 154000
rect 148244 154000 148272 154108
rect 150066 154096 150072 154148
rect 150124 154136 150130 154148
rect 150124 154108 156736 154136
rect 150124 154096 150130 154108
rect 152642 154028 152648 154080
rect 152700 154068 152706 154080
rect 155770 154068 155776 154080
rect 152700 154040 155776 154068
rect 152700 154028 152706 154040
rect 155770 154028 155776 154040
rect 155828 154028 155834 154080
rect 153194 154000 153200 154012
rect 148244 153972 153200 154000
rect 145156 153960 145162 153972
rect 153194 153960 153200 153972
rect 153252 153960 153258 154012
rect 156708 154000 156736 154108
rect 156874 154096 156880 154148
rect 156932 154136 156938 154148
rect 166258 154136 166264 154148
rect 156932 154108 166264 154136
rect 156932 154096 156938 154108
rect 166258 154096 166264 154108
rect 166316 154096 166322 154148
rect 166350 154096 166356 154148
rect 166408 154136 166414 154148
rect 245654 154136 245660 154148
rect 166408 154108 245660 154136
rect 166408 154096 166414 154108
rect 245654 154096 245660 154108
rect 245712 154096 245718 154148
rect 248598 154096 248604 154148
rect 248656 154136 248662 154148
rect 309226 154136 309232 154148
rect 248656 154108 309232 154136
rect 248656 154096 248662 154108
rect 309226 154096 309232 154108
rect 309284 154096 309290 154148
rect 326706 154096 326712 154148
rect 326764 154136 326770 154148
rect 368290 154136 368296 154148
rect 326764 154108 368296 154136
rect 326764 154096 326770 154108
rect 368290 154096 368296 154108
rect 368348 154096 368354 154148
rect 383654 154096 383660 154148
rect 383712 154136 383718 154148
rect 411990 154136 411996 154148
rect 383712 154108 411996 154136
rect 383712 154096 383718 154108
rect 411990 154096 411996 154108
rect 412048 154096 412054 154148
rect 156782 154028 156788 154080
rect 156840 154068 156846 154080
rect 235442 154068 235448 154080
rect 156840 154040 235448 154068
rect 156840 154028 156846 154040
rect 235442 154028 235448 154040
rect 235500 154028 235506 154080
rect 241882 154028 241888 154080
rect 241940 154068 241946 154080
rect 304074 154068 304080 154080
rect 241940 154040 304080 154068
rect 241940 154028 241946 154040
rect 304074 154028 304080 154040
rect 304132 154028 304138 154080
rect 323302 154028 323308 154080
rect 323360 154068 323366 154080
rect 365806 154068 365812 154080
rect 323360 154040 365812 154068
rect 323360 154028 323366 154040
rect 365806 154028 365812 154040
rect 365864 154028 365870 154080
rect 376846 154028 376852 154080
rect 376904 154068 376910 154080
rect 406838 154068 406844 154080
rect 376904 154040 406844 154068
rect 376904 154028 376910 154040
rect 406838 154028 406844 154040
rect 406896 154028 406902 154080
rect 233510 154000 233516 154012
rect 156708 153972 233516 154000
rect 233510 153960 233516 153972
rect 233568 153960 233574 154012
rect 235074 153960 235080 154012
rect 235132 154000 235138 154012
rect 299014 154000 299020 154012
rect 235132 153972 299020 154000
rect 235132 153960 235138 153972
rect 299014 153960 299020 153972
rect 299072 153960 299078 154012
rect 319254 153960 319260 154012
rect 319312 154000 319318 154012
rect 363230 154000 363236 154012
rect 319312 153972 363236 154000
rect 319312 153960 319318 153972
rect 363230 153960 363236 153972
rect 363288 153960 363294 154012
rect 369946 153960 369952 154012
rect 370004 154000 370010 154012
rect 401594 154000 401600 154012
rect 370004 153972 401600 154000
rect 370004 153960 370010 153972
rect 401594 153960 401600 153972
rect 401652 153960 401658 154012
rect 125560 153904 127112 153932
rect 125560 153892 125566 153904
rect 127158 153892 127164 153944
rect 127216 153932 127222 153944
rect 129458 153932 129464 153944
rect 127216 153904 129464 153932
rect 127216 153892 127222 153904
rect 129458 153892 129464 153904
rect 129516 153892 129522 153944
rect 129918 153892 129924 153944
rect 129976 153932 129982 153944
rect 218054 153932 218060 153944
rect 129976 153904 218060 153932
rect 129976 153892 129982 153904
rect 218054 153892 218060 153904
rect 218112 153892 218118 153944
rect 225046 153892 225052 153944
rect 225104 153932 225110 153944
rect 291378 153932 291384 153944
rect 225104 153904 291384 153932
rect 225104 153892 225110 153904
rect 291378 153892 291384 153904
rect 291436 153892 291442 153944
rect 313274 153892 313280 153944
rect 313332 153932 313338 153944
rect 357802 153932 357808 153944
rect 313332 153904 357808 153932
rect 313332 153892 313338 153904
rect 357802 153892 357808 153904
rect 357860 153892 357866 153944
rect 360378 153892 360384 153944
rect 360436 153932 360442 153944
rect 394050 153932 394056 153944
rect 360436 153904 394056 153932
rect 360436 153892 360442 153904
rect 394050 153892 394056 153904
rect 394108 153892 394114 153944
rect 397362 153892 397368 153944
rect 397420 153932 397426 153944
rect 422478 153932 422484 153944
rect 397420 153904 422484 153932
rect 397420 153892 397426 153904
rect 422478 153892 422484 153904
rect 422536 153892 422542 153944
rect 474 153824 480 153876
rect 532 153864 538 153876
rect 119798 153864 119804 153876
rect 532 153836 119804 153864
rect 532 153824 538 153836
rect 119798 153824 119804 153836
rect 119856 153824 119862 153876
rect 119890 153824 119896 153876
rect 119948 153864 119954 153876
rect 209774 153864 209780 153876
rect 119948 153836 209780 153864
rect 119948 153824 119954 153836
rect 209774 153824 209780 153836
rect 209832 153824 209838 153876
rect 215294 153824 215300 153876
rect 215352 153864 215358 153876
rect 283650 153864 283656 153876
rect 215352 153836 283656 153864
rect 215352 153824 215358 153836
rect 283650 153824 283656 153836
rect 283708 153824 283714 153876
rect 285674 153824 285680 153876
rect 285732 153864 285738 153876
rect 286134 153864 286140 153876
rect 285732 153836 286140 153864
rect 285732 153824 285738 153836
rect 286134 153824 286140 153836
rect 286192 153824 286198 153876
rect 286226 153824 286232 153876
rect 286284 153864 286290 153876
rect 334894 153864 334900 153876
rect 286284 153836 334900 153864
rect 286284 153824 286290 153836
rect 334894 153824 334900 153836
rect 334952 153824 334958 153876
rect 339494 153824 339500 153876
rect 339552 153864 339558 153876
rect 378594 153864 378600 153876
rect 339552 153836 378600 153864
rect 339552 153824 339558 153836
rect 378594 153824 378600 153836
rect 378652 153824 378658 153876
rect 380158 153824 380164 153876
rect 380216 153864 380222 153876
rect 409414 153864 409420 153876
rect 380216 153836 409420 153864
rect 380216 153824 380222 153836
rect 409414 153824 409420 153836
rect 409472 153824 409478 153876
rect 48314 153756 48320 153808
rect 48372 153796 48378 153808
rect 152642 153796 152648 153808
rect 48372 153768 152648 153796
rect 48372 153756 48378 153768
rect 152642 153756 152648 153768
rect 152700 153756 152706 153808
rect 152734 153756 152740 153808
rect 152792 153796 152798 153808
rect 212902 153796 212908 153808
rect 152792 153768 212908 153796
rect 152792 153756 152798 153768
rect 212902 153756 212908 153768
rect 212960 153756 212966 153808
rect 222378 153756 222384 153808
rect 222436 153796 222442 153808
rect 288710 153796 288716 153808
rect 222436 153768 288716 153796
rect 222436 153756 222442 153768
rect 288710 153756 288716 153768
rect 288768 153756 288774 153808
rect 363046 153756 363052 153808
rect 363104 153796 363110 153808
rect 396534 153796 396540 153808
rect 363104 153768 396540 153796
rect 363104 153756 363110 153768
rect 396534 153756 396540 153768
rect 396592 153756 396598 153808
rect 426434 153756 426440 153808
rect 426492 153796 426498 153808
rect 432414 153796 432420 153808
rect 426492 153768 432420 153796
rect 426492 153756 426498 153768
rect 432414 153756 432420 153768
rect 432472 153756 432478 153808
rect 57974 153688 57980 153740
rect 58032 153728 58038 153740
rect 153286 153728 153292 153740
rect 58032 153700 153292 153728
rect 58032 153688 58038 153700
rect 153286 153688 153292 153700
rect 153344 153688 153350 153740
rect 154482 153688 154488 153740
rect 154540 153728 154546 153740
rect 156506 153728 156512 153740
rect 154540 153700 156512 153728
rect 154540 153688 154546 153700
rect 156506 153688 156512 153700
rect 156564 153688 156570 153740
rect 156598 153688 156604 153740
rect 156656 153728 156662 153740
rect 210418 153728 210424 153740
rect 156656 153700 210424 153728
rect 156656 153688 156662 153700
rect 210418 153688 210424 153700
rect 210476 153688 210482 153740
rect 229094 153688 229100 153740
rect 229152 153728 229158 153740
rect 293862 153728 293868 153740
rect 229152 153700 293868 153728
rect 229152 153688 229158 153700
rect 293862 153688 293868 153700
rect 293920 153688 293926 153740
rect 64874 153620 64880 153672
rect 64932 153660 64938 153672
rect 165062 153660 165068 153672
rect 64932 153632 165068 153660
rect 64932 153620 64938 153632
rect 165062 153620 165068 153632
rect 165120 153620 165126 153672
rect 166258 153620 166264 153672
rect 166316 153660 166322 153672
rect 215478 153660 215484 153672
rect 166316 153632 215484 153660
rect 166316 153620 166322 153632
rect 215478 153620 215484 153632
rect 215536 153620 215542 153672
rect 238846 153620 238852 153672
rect 238904 153660 238910 153672
rect 301590 153660 301596 153672
rect 238904 153632 301596 153660
rect 238904 153620 238910 153632
rect 301590 153620 301596 153632
rect 301648 153620 301654 153672
rect 82814 153552 82820 153604
rect 82872 153592 82878 153604
rect 182082 153592 182088 153604
rect 82872 153564 182088 153592
rect 82872 153552 82878 153564
rect 182082 153552 182088 153564
rect 182140 153552 182146 153604
rect 182174 153552 182180 153604
rect 182232 153592 182238 153604
rect 185026 153592 185032 153604
rect 182232 153564 185032 153592
rect 182232 153552 182238 153564
rect 185026 153552 185032 153564
rect 185084 153552 185090 153604
rect 185118 153552 185124 153604
rect 185176 153592 185182 153604
rect 188338 153592 188344 153604
rect 185176 153564 188344 153592
rect 185176 153552 185182 153564
rect 188338 153552 188344 153564
rect 188396 153552 188402 153604
rect 188430 153552 188436 153604
rect 188488 153592 188494 153604
rect 197538 153592 197544 153604
rect 188488 153564 197544 153592
rect 188488 153552 188494 153564
rect 197538 153552 197544 153564
rect 197596 153552 197602 153604
rect 243722 153592 243728 153604
rect 197648 153564 243728 153592
rect 102134 153484 102140 153536
rect 102192 153524 102198 153536
rect 196894 153524 196900 153536
rect 102192 153496 196900 153524
rect 102192 153484 102198 153496
rect 196894 153484 196900 153496
rect 196952 153484 196958 153536
rect 196986 153484 196992 153536
rect 197044 153524 197050 153536
rect 197648 153524 197676 153564
rect 243722 153552 243728 153564
rect 243780 153552 243786 153604
rect 245930 153552 245936 153604
rect 245988 153592 245994 153604
rect 306650 153592 306656 153604
rect 245988 153564 306656 153592
rect 245988 153552 245994 153564
rect 306650 153552 306656 153564
rect 306708 153552 306714 153604
rect 197044 153496 197676 153524
rect 197044 153484 197050 153496
rect 198918 153484 198924 153536
rect 198976 153524 198982 153536
rect 248874 153524 248880 153536
rect 198976 153496 248880 153524
rect 198976 153484 198982 153496
rect 248874 153484 248880 153496
rect 248932 153484 248938 153536
rect 252646 153484 252652 153536
rect 252704 153524 252710 153536
rect 311802 153524 311808 153536
rect 252704 153496 311808 153524
rect 252704 153484 252710 153496
rect 311802 153484 311808 153496
rect 311860 153484 311866 153536
rect 331214 153484 331220 153536
rect 331272 153524 331278 153536
rect 337010 153524 337016 153536
rect 331272 153496 337016 153524
rect 331272 153484 331278 153496
rect 337010 153484 337016 153496
rect 337068 153484 337074 153536
rect 104894 153416 104900 153468
rect 104952 153456 104958 153468
rect 199470 153456 199476 153468
rect 104952 153428 199476 153456
rect 104952 153416 104958 153428
rect 199470 153416 199476 153428
rect 199528 153416 199534 153468
rect 201402 153416 201408 153468
rect 201460 153456 201466 153468
rect 256602 153456 256608 153468
rect 201460 153428 256608 153456
rect 201460 153416 201466 153428
rect 256602 153416 256608 153428
rect 256660 153416 256666 153468
rect 265434 153416 265440 153468
rect 265492 153456 265498 153468
rect 322198 153456 322204 153468
rect 265492 153428 322204 153456
rect 265492 153416 265498 153428
rect 322198 153416 322204 153428
rect 322256 153416 322262 153468
rect 108298 153348 108304 153400
rect 108356 153388 108362 153400
rect 191374 153388 191380 153400
rect 108356 153360 191380 153388
rect 108356 153348 108362 153360
rect 191374 153348 191380 153360
rect 191432 153348 191438 153400
rect 194502 153348 194508 153400
rect 194560 153388 194566 153400
rect 238662 153388 238668 153400
rect 194560 153360 238668 153388
rect 194560 153348 194566 153360
rect 238662 153348 238668 153360
rect 238720 153348 238726 153400
rect 259454 153348 259460 153400
rect 259512 153388 259518 153400
rect 316954 153388 316960 153400
rect 259512 153360 316960 153388
rect 259512 153348 259518 153360
rect 316954 153348 316960 153360
rect 317012 153348 317018 153400
rect 437566 153348 437572 153400
rect 437624 153388 437630 153400
rect 437624 153360 438532 153388
rect 437624 153348 437630 153360
rect 114830 153280 114836 153332
rect 114888 153320 114894 153332
rect 118602 153320 118608 153332
rect 114888 153292 118608 153320
rect 114888 153280 114894 153292
rect 118602 153280 118608 153292
rect 118660 153280 118666 153332
rect 118786 153280 118792 153332
rect 118844 153320 118850 153332
rect 119890 153320 119896 153332
rect 118844 153292 119896 153320
rect 118844 153280 118850 153292
rect 119890 153280 119896 153292
rect 119948 153280 119954 153332
rect 119982 153280 119988 153332
rect 120040 153320 120046 153332
rect 207198 153320 207204 153332
rect 120040 153292 207204 153320
rect 120040 153280 120046 153292
rect 207198 153280 207204 153292
rect 207256 153280 207262 153332
rect 272886 153280 272892 153332
rect 272944 153320 272950 153332
rect 327258 153320 327264 153332
rect 272944 153292 327264 153320
rect 272944 153280 272950 153292
rect 327258 153280 327264 153292
rect 327316 153280 327322 153332
rect 425974 153280 425980 153332
rect 426032 153320 426038 153332
rect 431310 153320 431316 153332
rect 426032 153292 431316 153320
rect 426032 153280 426038 153292
rect 431310 153280 431316 153292
rect 431368 153280 431374 153332
rect 437446 153292 437796 153320
rect 115934 153212 115940 153264
rect 115992 153252 115998 153264
rect 207842 153252 207848 153264
rect 115992 153224 118556 153252
rect 115992 153212 115998 153224
rect 118528 153184 118556 153224
rect 118804 153224 207848 153252
rect 118804 153184 118832 153224
rect 207842 153212 207848 153224
rect 207900 153212 207906 153264
rect 269206 153212 269212 153264
rect 269264 153252 269270 153264
rect 324682 153252 324688 153264
rect 269264 153224 324688 153252
rect 269264 153212 269270 153224
rect 324682 153212 324688 153224
rect 324740 153212 324746 153264
rect 428090 153252 428096 153264
rect 427786 153224 428096 153252
rect 118528 153156 118832 153184
rect 120074 153144 120080 153196
rect 120132 153184 120138 153196
rect 205910 153184 205916 153196
rect 120132 153156 205916 153184
rect 120132 153144 120138 153156
rect 205910 153144 205916 153156
rect 205968 153144 205974 153196
rect 223850 153144 223856 153196
rect 223908 153184 223914 153196
rect 288066 153184 288072 153196
rect 223908 153156 288072 153184
rect 223908 153144 223914 153156
rect 288066 153144 288072 153156
rect 288124 153144 288130 153196
rect 288250 153144 288256 153196
rect 288308 153184 288314 153196
rect 289998 153184 290004 153196
rect 288308 153156 290004 153184
rect 288308 153144 288314 153156
rect 289998 153144 290004 153156
rect 290056 153144 290062 153196
rect 303706 153144 303712 153196
rect 303764 153184 303770 153196
rect 350994 153184 351000 153196
rect 303764 153156 351000 153184
rect 303764 153144 303770 153156
rect 350994 153144 351000 153156
rect 351052 153144 351058 153196
rect 352006 153144 352012 153196
rect 352064 153184 352070 153196
rect 388254 153184 388260 153196
rect 352064 153156 388260 153184
rect 352064 153144 352070 153156
rect 388254 153144 388260 153156
rect 388312 153144 388318 153196
rect 389174 153144 389180 153196
rect 389232 153184 389238 153196
rect 412634 153184 412640 153196
rect 389232 153156 412640 153184
rect 389232 153144 389238 153156
rect 412634 153144 412640 153156
rect 412692 153144 412698 153196
rect 413094 153144 413100 153196
rect 413152 153184 413158 153196
rect 427786 153184 427814 153224
rect 428090 153212 428096 153224
rect 428148 153212 428154 153264
rect 431862 153212 431868 153264
rect 431920 153252 431926 153264
rect 431920 153224 433012 153252
rect 431920 153212 431926 153224
rect 413152 153156 427814 153184
rect 413152 153144 413158 153156
rect 427906 153144 427912 153196
rect 427964 153184 427970 153196
rect 432690 153184 432696 153196
rect 427964 153156 432696 153184
rect 427964 153144 427970 153156
rect 432690 153144 432696 153156
rect 432748 153144 432754 153196
rect 432984 153184 433012 153224
rect 433794 153184 433800 153196
rect 432984 153156 433800 153184
rect 433794 153144 433800 153156
rect 433852 153144 433858 153196
rect 434346 153144 434352 153196
rect 434404 153184 434410 153196
rect 437446 153184 437474 153292
rect 434404 153156 437474 153184
rect 434404 153144 434410 153156
rect 86862 153076 86868 153128
rect 86920 153116 86926 153128
rect 180242 153116 180248 153128
rect 86920 153088 180248 153116
rect 86920 153076 86926 153088
rect 180242 153076 180248 153088
rect 180300 153076 180306 153128
rect 180794 153076 180800 153128
rect 180852 153116 180858 153128
rect 257246 153116 257252 153128
rect 180852 153088 257252 153116
rect 180852 153076 180858 153088
rect 257246 153076 257252 153088
rect 257304 153076 257310 153128
rect 264974 153076 264980 153128
rect 265032 153116 265038 153128
rect 321462 153116 321468 153128
rect 265032 153088 321468 153116
rect 265032 153076 265038 153088
rect 321462 153076 321468 153088
rect 321520 153076 321526 153128
rect 324222 153076 324228 153128
rect 324280 153116 324286 153128
rect 366358 153116 366364 153128
rect 324280 153088 366364 153116
rect 324280 153076 324286 153088
rect 366358 153076 366364 153088
rect 366416 153076 366422 153128
rect 368474 153076 368480 153128
rect 368532 153116 368538 153128
rect 400398 153116 400404 153128
rect 368532 153088 400404 153116
rect 368532 153076 368538 153088
rect 400398 153076 400404 153088
rect 400456 153076 400462 153128
rect 403250 153076 403256 153128
rect 403308 153116 403314 153128
rect 415854 153116 415860 153128
rect 403308 153088 415860 153116
rect 403308 153076 403314 153088
rect 415854 153076 415860 153088
rect 415912 153076 415918 153128
rect 419258 153076 419264 153128
rect 419316 153116 419322 153128
rect 432782 153116 432788 153128
rect 419316 153088 432788 153116
rect 419316 153076 419322 153088
rect 432782 153076 432788 153088
rect 432840 153076 432846 153128
rect 436094 153076 436100 153128
rect 436152 153116 436158 153128
rect 437566 153116 437572 153128
rect 436152 153088 437572 153116
rect 436152 153076 436158 153088
rect 437566 153076 437572 153088
rect 437624 153076 437630 153128
rect 437768 153116 437796 153292
rect 437842 153144 437848 153196
rect 437900 153184 437906 153196
rect 438394 153184 438400 153196
rect 437900 153156 438400 153184
rect 437900 153144 437906 153156
rect 438394 153144 438400 153156
rect 438452 153144 438458 153196
rect 438504 153184 438532 153360
rect 440160 153224 440648 153252
rect 440160 153184 440188 153224
rect 438504 153156 440188 153184
rect 440234 153144 440240 153196
rect 440292 153184 440298 153196
rect 440510 153184 440516 153196
rect 440292 153156 440516 153184
rect 440292 153144 440298 153156
rect 440510 153144 440516 153156
rect 440568 153144 440574 153196
rect 440620 153184 440648 153224
rect 441982 153212 441988 153264
rect 442040 153252 442046 153264
rect 442040 153224 442580 153252
rect 442040 153212 442046 153224
rect 442166 153184 442172 153196
rect 440620 153156 442172 153184
rect 442166 153144 442172 153156
rect 442224 153144 442230 153196
rect 442552 153184 442580 153224
rect 449250 153184 449256 153196
rect 442552 153156 449256 153184
rect 449250 153144 449256 153156
rect 449308 153144 449314 153196
rect 453850 153144 453856 153196
rect 453908 153184 453914 153196
rect 459462 153184 459468 153196
rect 453908 153156 459468 153184
rect 453908 153144 453914 153156
rect 459462 153144 459468 153156
rect 459520 153144 459526 153196
rect 461854 153144 461860 153196
rect 461912 153184 461918 153196
rect 465902 153184 465908 153196
rect 461912 153156 465908 153184
rect 461912 153144 461918 153156
rect 465902 153144 465908 153156
rect 465960 153144 465966 153196
rect 466454 153144 466460 153196
rect 466512 153184 466518 153196
rect 469766 153184 469772 153196
rect 466512 153156 469772 153184
rect 466512 153144 466518 153156
rect 469766 153144 469772 153156
rect 469824 153144 469830 153196
rect 471422 153144 471428 153196
rect 471480 153184 471486 153196
rect 472986 153184 472992 153196
rect 471480 153156 472992 153184
rect 471480 153144 471486 153156
rect 472986 153144 472992 153156
rect 473044 153144 473050 153196
rect 473354 153144 473360 153196
rect 473412 153184 473418 153196
rect 475562 153184 475568 153196
rect 473412 153156 475568 153184
rect 473412 153144 473418 153156
rect 475562 153144 475568 153156
rect 475620 153144 475626 153196
rect 476114 153144 476120 153196
rect 476172 153184 476178 153196
rect 478138 153184 478144 153196
rect 476172 153156 478144 153184
rect 476172 153144 476178 153156
rect 478138 153144 478144 153156
rect 478196 153144 478202 153196
rect 485682 153144 485688 153196
rect 485740 153184 485746 153196
rect 489638 153184 489644 153196
rect 485740 153156 489644 153184
rect 485740 153144 485746 153156
rect 489638 153144 489644 153156
rect 489696 153144 489702 153196
rect 490742 153144 490748 153196
rect 490800 153184 490806 153196
rect 493502 153184 493508 153196
rect 490800 153156 493508 153184
rect 490800 153144 490806 153156
rect 493502 153144 493508 153156
rect 493560 153144 493566 153196
rect 494054 153144 494060 153196
rect 494112 153184 494118 153196
rect 496078 153184 496084 153196
rect 494112 153156 496084 153184
rect 494112 153144 494118 153156
rect 496078 153144 496084 153156
rect 496136 153144 496142 153196
rect 496630 153144 496636 153196
rect 496688 153184 496694 153196
rect 498010 153184 498016 153196
rect 496688 153156 498016 153184
rect 496688 153144 496694 153156
rect 498010 153144 498016 153156
rect 498068 153144 498074 153196
rect 512914 153144 512920 153196
rect 512972 153184 512978 153196
rect 515214 153184 515220 153196
rect 512972 153156 515220 153184
rect 512972 153144 512978 153156
rect 515214 153144 515220 153156
rect 515272 153144 515278 153196
rect 437768 153088 442120 153116
rect 103514 153008 103520 153060
rect 103572 153048 103578 153060
rect 198182 153048 198188 153060
rect 103572 153020 198188 153048
rect 103572 153008 103578 153020
rect 198182 153008 198188 153020
rect 198240 153008 198246 153060
rect 215386 153008 215392 153060
rect 215444 153048 215450 153060
rect 279694 153048 279700 153060
rect 215444 153020 279700 153048
rect 215444 153008 215450 153020
rect 279694 153008 279700 153020
rect 279752 153008 279758 153060
rect 291470 153008 291476 153060
rect 291528 153048 291534 153060
rect 335722 153048 335728 153060
rect 291528 153020 335728 153048
rect 291528 153008 291534 153020
rect 335722 153008 335728 153020
rect 335780 153008 335786 153060
rect 335832 153020 336044 153048
rect 96614 152940 96620 152992
rect 96672 152980 96678 152992
rect 193030 152980 193036 152992
rect 96672 152952 193036 152980
rect 96672 152940 96678 152952
rect 193030 152940 193036 152952
rect 193088 152940 193094 152992
rect 203702 152940 203708 152992
rect 203760 152980 203766 152992
rect 267550 152980 267556 152992
rect 203760 152952 267556 152980
rect 203760 152940 203766 152952
rect 267550 152940 267556 152952
rect 267608 152940 267614 152992
rect 272150 152940 272156 152992
rect 272208 152980 272214 152992
rect 320726 152980 320732 152992
rect 272208 152952 320732 152980
rect 272208 152940 272214 152952
rect 320726 152940 320732 152952
rect 320784 152940 320790 152992
rect 330938 152940 330944 152992
rect 330996 152980 331002 152992
rect 335832 152980 335860 153020
rect 330996 152952 335860 152980
rect 336016 152980 336044 153020
rect 336090 153008 336096 153060
rect 336148 153048 336154 153060
rect 347130 153048 347136 153060
rect 336148 153020 347136 153048
rect 336148 153008 336154 153020
rect 347130 153008 347136 153020
rect 347188 153008 347194 153060
rect 349154 153008 349160 153060
rect 349212 153048 349218 153060
rect 385586 153048 385592 153060
rect 349212 153020 385592 153048
rect 349212 153008 349218 153020
rect 385586 153008 385592 153020
rect 385644 153008 385650 153060
rect 386230 153008 386236 153060
rect 386288 153048 386294 153060
rect 399754 153048 399760 153060
rect 386288 153020 399760 153048
rect 386288 153008 386294 153020
rect 399754 153008 399760 153020
rect 399812 153008 399818 153060
rect 406654 153008 406660 153060
rect 406712 153048 406718 153060
rect 429286 153048 429292 153060
rect 406712 153020 429292 153048
rect 406712 153008 406718 153020
rect 429286 153008 429292 153020
rect 429344 153008 429350 153060
rect 431862 153048 431868 153060
rect 430500 153020 431868 153048
rect 371510 152980 371516 152992
rect 336016 152952 371516 152980
rect 330996 152940 331002 152952
rect 371510 152940 371516 152952
rect 371568 152940 371574 152992
rect 372614 152940 372620 152992
rect 372672 152980 372678 152992
rect 403618 152980 403624 152992
rect 372672 152952 403624 152980
rect 372672 152940 372678 152952
rect 403618 152940 403624 152952
rect 403676 152940 403682 152992
rect 404354 152940 404360 152992
rect 404412 152980 404418 152992
rect 427630 152980 427636 152992
rect 404412 152952 427636 152980
rect 404412 152940 404418 152952
rect 427630 152940 427636 152952
rect 427688 152940 427694 152992
rect 428090 152940 428096 152992
rect 428148 152980 428154 152992
rect 430500 152980 430528 153020
rect 431862 153008 431868 153020
rect 431920 153008 431926 153060
rect 431954 153008 431960 153060
rect 432012 153048 432018 153060
rect 441982 153048 441988 153060
rect 432012 153020 441988 153048
rect 432012 153008 432018 153020
rect 441982 153008 441988 153020
rect 442040 153008 442046 153060
rect 442092 153048 442120 153088
rect 442534 153076 442540 153128
rect 442592 153116 442598 153128
rect 443546 153116 443552 153128
rect 442592 153088 443552 153116
rect 442592 153076 442598 153088
rect 443546 153076 443552 153088
rect 443604 153076 443610 153128
rect 444466 153076 444472 153128
rect 444524 153116 444530 153128
rect 458266 153116 458272 153128
rect 444524 153088 458272 153116
rect 444524 153076 444530 153088
rect 458266 153076 458272 153088
rect 458324 153076 458330 153128
rect 462958 153076 462964 153128
rect 463016 153116 463022 153128
rect 467282 153116 467288 153128
rect 463016 153088 467288 153116
rect 463016 153076 463022 153088
rect 467282 153076 467288 153088
rect 467340 153076 467346 153128
rect 471238 153076 471244 153128
rect 471296 153116 471302 153128
rect 473630 153116 473636 153128
rect 471296 153088 473636 153116
rect 471296 153076 471302 153088
rect 473630 153076 473636 153088
rect 473688 153076 473694 153128
rect 474826 153076 474832 153128
rect 474884 153116 474890 153128
rect 476942 153116 476948 153128
rect 474884 153088 476948 153116
rect 474884 153076 474890 153088
rect 476942 153076 476948 153088
rect 477000 153076 477006 153128
rect 484026 153076 484032 153128
rect 484084 153116 484090 153128
rect 488442 153116 488448 153128
rect 484084 153088 488448 153116
rect 484084 153076 484090 153088
rect 488442 153076 488448 153088
rect 488500 153076 488506 153128
rect 489914 153076 489920 153128
rect 489972 153116 489978 153128
rect 492858 153116 492864 153128
rect 489972 153088 492864 153116
rect 489972 153076 489978 153088
rect 492858 153076 492864 153088
rect 492916 153076 492922 153128
rect 494146 153076 494152 153128
rect 494204 153116 494210 153128
rect 496722 153116 496728 153128
rect 494204 153088 496728 153116
rect 494204 153076 494210 153088
rect 496722 153076 496728 153088
rect 496780 153076 496786 153128
rect 496814 153076 496820 153128
rect 496872 153116 496878 153128
rect 498654 153116 498660 153128
rect 496872 153088 498660 153116
rect 496872 153076 496878 153088
rect 498654 153076 498660 153088
rect 498712 153076 498718 153128
rect 510982 153076 510988 153128
rect 511040 153116 511046 153128
rect 513466 153116 513472 153128
rect 511040 153088 513472 153116
rect 511040 153076 511046 153088
rect 513466 153076 513472 153088
rect 513524 153076 513530 153128
rect 514202 153076 514208 153128
rect 514260 153116 514266 153128
rect 517422 153116 517428 153128
rect 514260 153088 517428 153116
rect 514260 153076 514266 153088
rect 517422 153076 517428 153088
rect 517480 153076 517486 153128
rect 442258 153048 442264 153060
rect 442092 153020 442264 153048
rect 442258 153008 442264 153020
rect 442316 153008 442322 153060
rect 449894 153048 449900 153060
rect 442460 153020 449900 153048
rect 428148 152952 430528 152980
rect 428148 152940 428154 152952
rect 430574 152940 430580 152992
rect 430632 152980 430638 152992
rect 442350 152980 442356 152992
rect 430632 152952 442356 152980
rect 430632 152940 430638 152952
rect 442350 152940 442356 152952
rect 442408 152940 442414 152992
rect 89806 152872 89812 152924
rect 89864 152912 89870 152924
rect 187878 152912 187884 152924
rect 89864 152884 187884 152912
rect 89864 152872 89870 152884
rect 187878 152872 187884 152884
rect 187936 152872 187942 152924
rect 191650 152872 191656 152924
rect 191708 152912 191714 152924
rect 208486 152912 208492 152924
rect 191708 152884 208492 152912
rect 191708 152872 191714 152884
rect 208486 152872 208492 152884
rect 208544 152872 208550 152924
rect 212442 152872 212448 152924
rect 212500 152912 212506 152924
rect 277762 152912 277768 152924
rect 212500 152884 277768 152912
rect 212500 152872 212506 152884
rect 277762 152872 277768 152884
rect 277820 152872 277826 152924
rect 285490 152872 285496 152924
rect 285548 152912 285554 152924
rect 335814 152912 335820 152924
rect 285548 152884 335820 152912
rect 285548 152872 285554 152884
rect 335814 152872 335820 152884
rect 335872 152872 335878 152924
rect 335906 152872 335912 152924
rect 335964 152912 335970 152924
rect 341334 152912 341340 152924
rect 335964 152884 341340 152912
rect 335964 152872 335970 152884
rect 341334 152872 341340 152884
rect 341392 152872 341398 152924
rect 341426 152872 341432 152924
rect 341484 152912 341490 152924
rect 377306 152912 377312 152924
rect 341484 152884 377312 152912
rect 341484 152872 341490 152884
rect 377306 152872 377312 152884
rect 377364 152872 377370 152924
rect 378226 152872 378232 152924
rect 378284 152912 378290 152924
rect 379882 152912 379888 152924
rect 378284 152884 379888 152912
rect 378284 152872 378290 152884
rect 379882 152872 379888 152884
rect 379940 152872 379946 152924
rect 380894 152872 380900 152924
rect 380952 152912 380958 152924
rect 410058 152912 410064 152924
rect 380952 152884 410064 152912
rect 380952 152872 380958 152884
rect 410058 152872 410064 152884
rect 410116 152872 410122 152924
rect 411254 152872 411260 152924
rect 411312 152912 411318 152924
rect 433150 152912 433156 152924
rect 411312 152884 433156 152912
rect 411312 152872 411318 152884
rect 433150 152872 433156 152884
rect 433208 152872 433214 152924
rect 433518 152872 433524 152924
rect 433576 152912 433582 152924
rect 442460 152912 442488 153020
rect 449894 153008 449900 153020
rect 449952 153008 449958 153060
rect 456886 153008 456892 153060
rect 456944 153048 456950 153060
rect 460750 153048 460756 153060
rect 456944 153020 460756 153048
rect 456944 153008 456950 153020
rect 460750 153008 460756 153020
rect 460808 153008 460814 153060
rect 463510 153008 463516 153060
rect 463568 153048 463574 153060
rect 466546 153048 466552 153060
rect 463568 153020 466552 153048
rect 463568 153008 463574 153020
rect 466546 153008 466552 153020
rect 466604 153008 466610 153060
rect 466638 153008 466644 153060
rect 466696 153048 466702 153060
rect 470410 153048 470416 153060
rect 466696 153020 470416 153048
rect 466696 153008 466702 153020
rect 470410 153008 470416 153020
rect 470468 153008 470474 153060
rect 472342 153008 472348 153060
rect 472400 153048 472406 153060
rect 474918 153048 474924 153060
rect 472400 153020 474924 153048
rect 472400 153008 472406 153020
rect 474918 153008 474924 153020
rect 474976 153008 474982 153060
rect 484486 153008 484492 153060
rect 484544 153048 484550 153060
rect 488994 153048 489000 153060
rect 484544 153020 489000 153048
rect 484544 153008 484550 153020
rect 488994 153008 489000 153020
rect 489052 153008 489058 153060
rect 492674 153008 492680 153060
rect 492732 153048 492738 153060
rect 495434 153048 495440 153060
rect 492732 153020 495440 153048
rect 492732 153008 492738 153020
rect 495434 153008 495440 153020
rect 495492 153008 495498 153060
rect 495526 153008 495532 153060
rect 495584 153048 495590 153060
rect 497366 153048 497372 153060
rect 495584 153020 497372 153048
rect 495584 153008 495590 153020
rect 497366 153008 497372 153020
rect 497424 153008 497430 153060
rect 442534 152940 442540 152992
rect 442592 152980 442598 152992
rect 447962 152980 447968 152992
rect 442592 152952 447968 152980
rect 442592 152940 442598 152952
rect 447962 152940 447968 152952
rect 448020 152940 448026 152992
rect 463878 152940 463884 152992
rect 463936 152980 463942 152992
rect 468386 152980 468392 152992
rect 463936 152952 468392 152980
rect 463936 152940 463942 152952
rect 468386 152940 468392 152952
rect 468444 152940 468450 152992
rect 472434 152940 472440 152992
rect 472492 152980 472498 152992
rect 474274 152980 474280 152992
rect 472492 152952 474280 152980
rect 472492 152940 472498 152952
rect 474274 152940 474280 152952
rect 474332 152940 474338 152992
rect 483106 152940 483112 152992
rect 483164 152980 483170 152992
rect 487798 152980 487804 152992
rect 483164 152952 487804 152980
rect 483164 152940 483170 152952
rect 487798 152940 487804 152952
rect 487856 152940 487862 152992
rect 491662 152940 491668 152992
rect 491720 152980 491726 152992
rect 494790 152980 494796 152992
rect 491720 152952 494796 152980
rect 491720 152940 491726 152952
rect 494790 152940 494796 152952
rect 494848 152940 494854 152992
rect 512270 152940 512276 152992
rect 512328 152980 512334 152992
rect 514754 152980 514760 152992
rect 512328 152952 514760 152980
rect 512328 152940 512334 152952
rect 514754 152940 514760 152952
rect 514812 152940 514818 152992
rect 433576 152884 442488 152912
rect 433576 152872 433582 152884
rect 443178 152872 443184 152924
rect 443236 152912 443242 152924
rect 451182 152912 451188 152924
rect 443236 152884 451188 152912
rect 443236 152872 443242 152884
rect 451182 152872 451188 152884
rect 451240 152872 451246 152924
rect 459646 152872 459652 152924
rect 459704 152912 459710 152924
rect 464614 152912 464620 152924
rect 459704 152884 464620 152912
rect 459704 152872 459710 152884
rect 464614 152872 464620 152884
rect 464672 152872 464678 152924
rect 465074 152872 465080 152924
rect 465132 152912 465138 152924
rect 469122 152912 469128 152924
rect 465132 152884 469128 152912
rect 465132 152872 465138 152884
rect 469122 152872 469128 152884
rect 469180 152872 469186 152924
rect 491294 152872 491300 152924
rect 491352 152912 491358 152924
rect 494146 152912 494152 152924
rect 491352 152884 494152 152912
rect 491352 152872 491358 152884
rect 494146 152872 494152 152884
rect 494204 152872 494210 152924
rect 513558 152872 513564 152924
rect 513616 152912 513622 152924
rect 516134 152912 516140 152924
rect 513616 152884 516140 152912
rect 513616 152872 513622 152884
rect 516134 152872 516140 152884
rect 516192 152872 516198 152924
rect 66254 152804 66260 152856
rect 66312 152844 66318 152856
rect 169938 152844 169944 152856
rect 66312 152816 169944 152844
rect 66312 152804 66318 152816
rect 169938 152804 169944 152816
rect 169996 152804 170002 152856
rect 173894 152804 173900 152856
rect 173952 152844 173958 152856
rect 252094 152844 252100 152856
rect 173952 152816 252100 152844
rect 173952 152804 173958 152816
rect 252094 152804 252100 152816
rect 252152 152804 252158 152856
rect 257706 152804 257712 152856
rect 257764 152844 257770 152856
rect 315666 152844 315672 152856
rect 257764 152816 315672 152844
rect 257764 152804 257770 152816
rect 315666 152804 315672 152816
rect 315724 152804 315730 152856
rect 317046 152804 317052 152856
rect 317104 152844 317110 152856
rect 318242 152844 318248 152856
rect 317104 152816 318248 152844
rect 317104 152804 317110 152816
rect 318242 152804 318248 152816
rect 318300 152804 318306 152856
rect 318334 152804 318340 152856
rect 318392 152844 318398 152856
rect 361942 152844 361948 152856
rect 318392 152816 361948 152844
rect 318392 152804 318398 152816
rect 361942 152804 361948 152816
rect 362000 152804 362006 152856
rect 365714 152804 365720 152856
rect 365772 152844 365778 152856
rect 367002 152844 367008 152856
rect 365772 152816 367008 152844
rect 365772 152804 365778 152816
rect 367002 152804 367008 152816
rect 367060 152804 367066 152856
rect 367186 152804 367192 152856
rect 367244 152844 367250 152856
rect 368934 152844 368940 152856
rect 367244 152816 368940 152844
rect 367244 152804 367250 152816
rect 368934 152804 368940 152816
rect 368992 152804 368998 152856
rect 369026 152804 369032 152856
rect 369084 152844 369090 152856
rect 397178 152844 397184 152856
rect 369084 152816 397184 152844
rect 369084 152804 369090 152816
rect 397178 152804 397184 152816
rect 397236 152804 397242 152856
rect 401686 152804 401692 152856
rect 401744 152844 401750 152856
rect 426158 152844 426164 152856
rect 401744 152816 426164 152844
rect 401744 152804 401750 152816
rect 426158 152804 426164 152816
rect 426216 152804 426222 152856
rect 426342 152804 426348 152856
rect 426400 152844 426406 152856
rect 426400 152816 430160 152844
rect 426400 152804 426406 152816
rect 26418 152736 26424 152788
rect 26476 152776 26482 152788
rect 139118 152776 139124 152788
rect 26476 152748 139124 152776
rect 26476 152736 26482 152748
rect 139118 152736 139124 152748
rect 139176 152736 139182 152788
rect 139394 152736 139400 152788
rect 139452 152776 139458 152788
rect 141694 152776 141700 152788
rect 139452 152748 141700 152776
rect 139452 152736 139458 152748
rect 141694 152736 141700 152748
rect 141752 152736 141758 152788
rect 146846 152776 146852 152788
rect 141804 152748 146852 152776
rect 22186 152668 22192 152720
rect 22244 152708 22250 152720
rect 135898 152708 135904 152720
rect 22244 152680 135904 152708
rect 22244 152668 22250 152680
rect 135898 152668 135904 152680
rect 135956 152668 135962 152720
rect 141804 152708 141832 152748
rect 146846 152736 146852 152748
rect 146904 152736 146910 152788
rect 149054 152736 149060 152788
rect 149112 152776 149118 152788
rect 231578 152776 231584 152788
rect 149112 152748 231584 152776
rect 149112 152736 149118 152748
rect 231578 152736 231584 152748
rect 231636 152736 231642 152788
rect 240318 152736 240324 152788
rect 240376 152776 240382 152788
rect 241882 152776 241888 152788
rect 240376 152748 241888 152776
rect 240376 152736 240382 152748
rect 241882 152736 241888 152748
rect 241940 152736 241946 152788
rect 244366 152736 244372 152788
rect 244424 152776 244430 152788
rect 306006 152776 306012 152788
rect 244424 152748 306012 152776
rect 244424 152736 244430 152748
rect 306006 152736 306012 152748
rect 306064 152736 306070 152788
rect 307662 152736 307668 152788
rect 307720 152776 307726 152788
rect 352282 152776 352288 152788
rect 307720 152748 352288 152776
rect 307720 152736 307726 152748
rect 352282 152736 352288 152748
rect 352340 152736 352346 152788
rect 357434 152736 357440 152788
rect 357492 152776 357498 152788
rect 359366 152776 359372 152788
rect 357492 152748 359372 152776
rect 357492 152736 357498 152748
rect 359366 152736 359372 152748
rect 359424 152736 359430 152788
rect 359458 152736 359464 152788
rect 359516 152776 359522 152788
rect 390186 152776 390192 152788
rect 359516 152748 390192 152776
rect 359516 152736 359522 152748
rect 390186 152736 390192 152748
rect 390244 152736 390250 152788
rect 415210 152776 415216 152788
rect 394160 152748 415216 152776
rect 136008 152680 141832 152708
rect 15194 152600 15200 152652
rect 15252 152640 15258 152652
rect 130746 152640 130752 152652
rect 15252 152612 130752 152640
rect 15252 152600 15258 152612
rect 130746 152600 130752 152612
rect 130804 152600 130810 152652
rect 135162 152600 135168 152652
rect 135220 152640 135226 152652
rect 136008 152640 136036 152680
rect 141878 152668 141884 152720
rect 141936 152708 141942 152720
rect 151906 152708 151912 152720
rect 141936 152680 151912 152708
rect 141936 152668 141942 152680
rect 151906 152668 151912 152680
rect 151964 152668 151970 152720
rect 153562 152668 153568 152720
rect 153620 152708 153626 152720
rect 236730 152708 236736 152720
rect 153620 152680 236736 152708
rect 153620 152668 153626 152680
rect 236730 152668 236736 152680
rect 236788 152668 236794 152720
rect 247034 152668 247040 152720
rect 247092 152708 247098 152720
rect 307938 152708 307944 152720
rect 247092 152680 307944 152708
rect 247092 152668 247098 152680
rect 307938 152668 307944 152680
rect 307996 152668 308002 152720
rect 311526 152668 311532 152720
rect 311584 152708 311590 152720
rect 356790 152708 356796 152720
rect 311584 152680 356796 152708
rect 311584 152668 311590 152680
rect 356790 152668 356796 152680
rect 356848 152668 356854 152720
rect 358814 152668 358820 152720
rect 358872 152708 358878 152720
rect 393406 152708 393412 152720
rect 358872 152680 393412 152708
rect 358872 152668 358878 152680
rect 393406 152668 393412 152680
rect 393464 152668 393470 152720
rect 135220 152612 136036 152640
rect 135220 152600 135226 152612
rect 136910 152600 136916 152652
rect 136968 152640 136974 152652
rect 137186 152640 137192 152652
rect 136968 152612 137192 152640
rect 136968 152600 136974 152612
rect 137186 152600 137192 152612
rect 137244 152600 137250 152652
rect 216122 152640 216128 152652
rect 137296 152612 216128 152640
rect 19334 152532 19340 152584
rect 19392 152572 19398 152584
rect 133966 152572 133972 152584
rect 19392 152544 133972 152572
rect 19392 152532 19398 152544
rect 133966 152532 133972 152544
rect 134024 152532 134030 152584
rect 2866 152464 2872 152516
rect 2924 152504 2930 152516
rect 121086 152504 121092 152516
rect 2924 152476 121092 152504
rect 2924 152464 2930 152476
rect 121086 152464 121092 152476
rect 121144 152464 121150 152516
rect 129734 152464 129740 152516
rect 129792 152504 129798 152516
rect 137296 152504 137324 152612
rect 216122 152600 216128 152612
rect 216180 152600 216186 152652
rect 220446 152600 220452 152652
rect 220504 152640 220510 152652
rect 284846 152640 284852 152652
rect 220504 152612 284852 152640
rect 220504 152600 220510 152612
rect 284846 152600 284852 152612
rect 284904 152600 284910 152652
rect 285766 152600 285772 152652
rect 285824 152640 285830 152652
rect 291838 152640 291844 152652
rect 285824 152612 291844 152640
rect 285824 152600 285830 152612
rect 291838 152600 291844 152612
rect 291896 152600 291902 152652
rect 292206 152600 292212 152652
rect 292264 152640 292270 152652
rect 341978 152640 341984 152652
rect 292264 152612 341984 152640
rect 292264 152600 292270 152612
rect 341978 152600 341984 152612
rect 342036 152600 342042 152652
rect 342254 152600 342260 152652
rect 342312 152640 342318 152652
rect 343910 152640 343916 152652
rect 342312 152612 343916 152640
rect 342312 152600 342318 152612
rect 343910 152600 343916 152612
rect 343968 152600 343974 152652
rect 345290 152600 345296 152652
rect 345348 152640 345354 152652
rect 382458 152640 382464 152652
rect 345348 152612 382464 152640
rect 345348 152600 345354 152612
rect 382458 152600 382464 152612
rect 382516 152600 382522 152652
rect 386414 152600 386420 152652
rect 386472 152640 386478 152652
rect 386472 152612 389864 152640
rect 386472 152600 386478 152612
rect 140774 152532 140780 152584
rect 140832 152572 140838 152584
rect 140832 152544 142154 152572
rect 140832 152532 140838 152544
rect 129792 152476 137324 152504
rect 129792 152464 129798 152476
rect 137554 152464 137560 152516
rect 137612 152504 137618 152516
rect 141142 152504 141148 152516
rect 137612 152476 141148 152504
rect 137612 152464 137618 152476
rect 141142 152464 141148 152476
rect 141200 152464 141206 152516
rect 142126 152504 142154 152544
rect 146938 152532 146944 152584
rect 146996 152572 147002 152584
rect 221274 152572 221280 152584
rect 146996 152544 221280 152572
rect 146996 152532 147002 152544
rect 221274 152532 221280 152544
rect 221332 152532 221338 152584
rect 225230 152532 225236 152584
rect 225288 152572 225294 152584
rect 229002 152572 229008 152584
rect 225288 152544 229008 152572
rect 225288 152532 225294 152544
rect 229002 152532 229008 152544
rect 229060 152532 229066 152584
rect 234154 152532 234160 152584
rect 234212 152572 234218 152584
rect 297726 152572 297732 152584
rect 234212 152544 297732 152572
rect 234212 152532 234218 152544
rect 297726 152532 297732 152544
rect 297784 152532 297790 152584
rect 304810 152532 304816 152584
rect 304868 152572 304874 152584
rect 351638 152572 351644 152584
rect 304868 152544 351644 152572
rect 304868 152532 304874 152544
rect 351638 152532 351644 152544
rect 351696 152532 351702 152584
rect 354490 152532 354496 152584
rect 354548 152572 354554 152584
rect 389542 152572 389548 152584
rect 354548 152544 389548 152572
rect 354548 152532 354554 152544
rect 389542 152532 389548 152544
rect 389600 152532 389606 152584
rect 389836 152572 389864 152612
rect 390370 152600 390376 152652
rect 390428 152640 390434 152652
rect 394160 152640 394188 152748
rect 415210 152736 415216 152748
rect 415268 152736 415274 152788
rect 415394 152736 415400 152788
rect 415452 152776 415458 152788
rect 427814 152776 427820 152788
rect 415452 152748 427820 152776
rect 415452 152736 415458 152748
rect 427814 152736 427820 152748
rect 427872 152736 427878 152788
rect 430022 152776 430028 152788
rect 427924 152748 430028 152776
rect 395522 152668 395528 152720
rect 395580 152708 395586 152720
rect 397822 152708 397828 152720
rect 395580 152680 397828 152708
rect 395580 152668 395586 152680
rect 397822 152668 397828 152680
rect 397880 152668 397886 152720
rect 399110 152668 399116 152720
rect 399168 152708 399174 152720
rect 424226 152708 424232 152720
rect 399168 152680 424232 152708
rect 399168 152668 399174 152680
rect 424226 152668 424232 152680
rect 424284 152668 424290 152720
rect 413922 152640 413928 152652
rect 390428 152612 394188 152640
rect 394712 152612 413928 152640
rect 390428 152600 390434 152612
rect 394712 152572 394740 152612
rect 413922 152600 413928 152612
rect 413980 152600 413986 152652
rect 414382 152600 414388 152652
rect 414440 152640 414446 152652
rect 427924 152640 427952 152748
rect 430022 152736 430028 152748
rect 430080 152736 430086 152788
rect 430132 152776 430160 152816
rect 430206 152804 430212 152856
rect 430264 152844 430270 152856
rect 447318 152844 447324 152856
rect 430264 152816 447324 152844
rect 430264 152804 430270 152816
rect 447318 152804 447324 152816
rect 447376 152804 447382 152856
rect 510338 152804 510344 152856
rect 510396 152844 510402 152856
rect 511994 152844 512000 152856
rect 510396 152816 512000 152844
rect 510396 152804 510402 152816
rect 511994 152804 512000 152816
rect 512052 152804 512058 152856
rect 434530 152776 434536 152788
rect 430132 152748 434536 152776
rect 434530 152736 434536 152748
rect 434588 152736 434594 152788
rect 434714 152736 434720 152788
rect 434772 152776 434778 152788
rect 434772 152748 438808 152776
rect 434772 152736 434778 152748
rect 428182 152668 428188 152720
rect 428240 152708 428246 152720
rect 438780 152708 438808 152748
rect 438854 152736 438860 152788
rect 438912 152776 438918 152788
rect 454402 152776 454408 152788
rect 438912 152748 454408 152776
rect 438912 152736 438918 152748
rect 454402 152736 454408 152748
rect 454460 152736 454466 152788
rect 511626 152736 511632 152788
rect 511684 152776 511690 152788
rect 513742 152776 513748 152788
rect 511684 152748 513748 152776
rect 511684 152736 511690 152748
rect 513742 152736 513748 152748
rect 513800 152736 513806 152788
rect 440234 152708 440240 152720
rect 428240 152680 437474 152708
rect 438780 152680 440240 152708
rect 428240 152668 428246 152680
rect 437106 152640 437112 152652
rect 414440 152612 427952 152640
rect 428016 152612 437112 152640
rect 414440 152600 414446 152612
rect 389836 152544 394740 152572
rect 394878 152532 394884 152584
rect 394936 152572 394942 152584
rect 420362 152572 420368 152584
rect 394936 152544 420368 152572
rect 394936 152532 394942 152544
rect 420362 152532 420368 152544
rect 420420 152532 420426 152584
rect 423398 152532 423404 152584
rect 423456 152572 423462 152584
rect 428016 152572 428044 152612
rect 437106 152600 437112 152612
rect 437164 152600 437170 152652
rect 437446 152640 437474 152680
rect 440234 152668 440240 152680
rect 440292 152668 440298 152720
rect 440326 152668 440332 152720
rect 440384 152708 440390 152720
rect 445478 152708 445484 152720
rect 440384 152680 445484 152708
rect 440384 152668 440390 152680
rect 445478 152668 445484 152680
rect 445536 152668 445542 152720
rect 441430 152640 441436 152652
rect 437446 152612 441436 152640
rect 441430 152600 441436 152612
rect 441488 152600 441494 152652
rect 441614 152600 441620 152652
rect 441672 152640 441678 152652
rect 444742 152640 444748 152652
rect 441672 152612 444748 152640
rect 441672 152600 441678 152612
rect 444742 152600 444748 152612
rect 444800 152600 444806 152652
rect 459554 152600 459560 152652
rect 459612 152640 459618 152652
rect 465258 152640 465264 152652
rect 459612 152612 465264 152640
rect 459612 152600 459618 152612
rect 465258 152600 465264 152612
rect 465316 152600 465322 152652
rect 423456 152544 428044 152572
rect 423456 152532 423462 152544
rect 429838 152532 429844 152584
rect 429896 152572 429902 152584
rect 441522 152572 441528 152584
rect 429896 152544 441528 152572
rect 429896 152532 429902 152544
rect 441522 152532 441528 152544
rect 441580 152532 441586 152584
rect 442074 152532 442080 152584
rect 442132 152572 442138 152584
rect 444650 152572 444656 152584
rect 442132 152544 444656 152572
rect 442132 152532 442138 152544
rect 444650 152532 444656 152544
rect 444708 152532 444714 152584
rect 445570 152532 445576 152584
rect 445628 152572 445634 152584
rect 456978 152572 456984 152584
rect 445628 152544 456984 152572
rect 445628 152532 445634 152544
rect 456978 152532 456984 152544
rect 457036 152532 457042 152584
rect 458174 152532 458180 152584
rect 458232 152572 458238 152584
rect 463970 152572 463976 152584
rect 458232 152544 463976 152572
rect 458232 152532 458238 152544
rect 463970 152532 463976 152544
rect 464028 152532 464034 152584
rect 226426 152504 226432 152516
rect 142126 152476 226432 152504
rect 226426 152464 226432 152476
rect 226484 152464 226490 152516
rect 227898 152464 227904 152516
rect 227956 152504 227962 152516
rect 293218 152504 293224 152516
rect 227956 152476 293224 152504
rect 227956 152464 227962 152476
rect 293218 152464 293224 152476
rect 293276 152464 293282 152516
rect 298646 152464 298652 152516
rect 298704 152504 298710 152516
rect 335906 152504 335912 152516
rect 298704 152476 335912 152504
rect 298704 152464 298710 152476
rect 335906 152464 335912 152476
rect 335964 152464 335970 152516
rect 335998 152464 336004 152516
rect 336056 152504 336062 152516
rect 346486 152504 346492 152516
rect 336056 152476 346492 152504
rect 336056 152464 336062 152476
rect 346486 152464 346492 152476
rect 346544 152464 346550 152516
rect 347958 152464 347964 152516
rect 348016 152504 348022 152516
rect 385034 152504 385040 152516
rect 348016 152476 385040 152504
rect 348016 152464 348022 152476
rect 385034 152464 385040 152476
rect 385092 152464 385098 152516
rect 385310 152464 385316 152516
rect 385368 152504 385374 152516
rect 387610 152504 387616 152516
rect 385368 152476 387616 152504
rect 385368 152464 385374 152476
rect 387610 152464 387616 152476
rect 387668 152464 387674 152516
rect 393130 152464 393136 152516
rect 393188 152504 393194 152516
rect 419074 152504 419080 152516
rect 393188 152476 419080 152504
rect 393188 152464 393194 152476
rect 419074 152464 419080 152476
rect 419132 152464 419138 152516
rect 421190 152464 421196 152516
rect 421248 152504 421254 152516
rect 432598 152504 432604 152516
rect 421248 152476 432604 152504
rect 421248 152464 421254 152476
rect 432598 152464 432604 152476
rect 432656 152464 432662 152516
rect 432690 152464 432696 152516
rect 432748 152504 432754 152516
rect 432748 152476 436140 152504
rect 432748 152464 432754 152476
rect 59998 152396 60004 152448
rect 60056 152436 60062 152448
rect 144270 152436 144276 152448
rect 60056 152408 144276 152436
rect 60056 152396 60062 152408
rect 144270 152396 144276 152408
rect 144328 152396 144334 152448
rect 144822 152396 144828 152448
rect 144880 152436 144886 152448
rect 162210 152436 162216 152448
rect 144880 152408 162216 152436
rect 144880 152396 144886 152408
rect 162210 152396 162216 152408
rect 162268 152396 162274 152448
rect 164326 152396 164332 152448
rect 164384 152436 164390 152448
rect 244366 152436 244372 152448
rect 164384 152408 244372 152436
rect 164384 152396 164390 152408
rect 244366 152396 244372 152408
rect 244424 152396 244430 152448
rect 251174 152396 251180 152448
rect 251232 152436 251238 152448
rect 311158 152436 311164 152448
rect 251232 152408 311164 152436
rect 251232 152396 251238 152408
rect 311158 152396 311164 152408
rect 311216 152396 311222 152448
rect 311986 152396 311992 152448
rect 312044 152436 312050 152448
rect 356146 152436 356152 152448
rect 312044 152408 356152 152436
rect 312044 152396 312050 152408
rect 356146 152396 356152 152408
rect 356204 152396 356210 152448
rect 361574 152396 361580 152448
rect 361632 152436 361638 152448
rect 395338 152436 395344 152448
rect 361632 152408 395344 152436
rect 361632 152396 361638 152408
rect 395338 152396 395344 152408
rect 395396 152396 395402 152448
rect 398834 152396 398840 152448
rect 398892 152436 398898 152448
rect 413278 152436 413284 152448
rect 398892 152408 413284 152436
rect 398892 152396 398898 152408
rect 413278 152396 413284 152408
rect 413336 152396 413342 152448
rect 413830 152396 413836 152448
rect 413888 152436 413894 152448
rect 416498 152436 416504 152448
rect 413888 152408 416504 152436
rect 413888 152396 413894 152408
rect 416498 152396 416504 152408
rect 416556 152396 416562 152448
rect 418430 152396 418436 152448
rect 418488 152436 418494 152448
rect 418488 152408 429976 152436
rect 418488 152396 418494 152408
rect 113174 152328 113180 152380
rect 113232 152368 113238 152380
rect 120074 152368 120080 152380
rect 113232 152340 120080 152368
rect 113232 152328 113238 152340
rect 120074 152328 120080 152340
rect 120132 152328 120138 152380
rect 120166 152328 120172 152380
rect 120224 152368 120230 152380
rect 211062 152368 211068 152380
rect 120224 152340 211068 152368
rect 120224 152328 120230 152340
rect 211062 152328 211068 152340
rect 211120 152328 211126 152380
rect 221734 152328 221740 152380
rect 221792 152368 221798 152380
rect 282914 152368 282920 152380
rect 221792 152340 282920 152368
rect 221792 152328 221798 152340
rect 282914 152328 282920 152340
rect 282972 152328 282978 152380
rect 283190 152328 283196 152380
rect 283248 152368 283254 152380
rect 287422 152368 287428 152380
rect 283248 152340 287428 152368
rect 283248 152328 283254 152340
rect 287422 152328 287428 152340
rect 287480 152328 287486 152380
rect 291838 152328 291844 152380
rect 291896 152368 291902 152380
rect 336182 152368 336188 152380
rect 291896 152340 336188 152368
rect 291896 152328 291902 152340
rect 336182 152328 336188 152340
rect 336240 152328 336246 152380
rect 343634 152328 343640 152380
rect 343692 152368 343698 152380
rect 380526 152368 380532 152380
rect 343692 152340 380532 152368
rect 343692 152328 343698 152340
rect 380526 152328 380532 152340
rect 380584 152328 380590 152380
rect 381446 152328 381452 152380
rect 381504 152368 381510 152380
rect 410702 152368 410708 152380
rect 381504 152340 410708 152368
rect 381504 152328 381510 152340
rect 410702 152328 410708 152340
rect 410760 152328 410766 152380
rect 413186 152328 413192 152380
rect 413244 152368 413250 152380
rect 421650 152368 421656 152380
rect 413244 152340 421656 152368
rect 413244 152328 413250 152340
rect 421650 152328 421656 152340
rect 421708 152328 421714 152380
rect 425146 152328 425152 152380
rect 425204 152368 425210 152380
rect 429948 152368 429976 152408
rect 430022 152396 430028 152448
rect 430080 152436 430086 152448
rect 435726 152436 435732 152448
rect 430080 152408 435732 152436
rect 430080 152396 430086 152408
rect 435726 152396 435732 152408
rect 435784 152396 435790 152448
rect 436112 152436 436140 152476
rect 436186 152464 436192 152516
rect 436244 152504 436250 152516
rect 444558 152504 444564 152516
rect 436244 152476 444564 152504
rect 436244 152464 436250 152476
rect 444558 152464 444564 152476
rect 444616 152464 444622 152516
rect 445478 152464 445484 152516
rect 445536 152504 445542 152516
rect 455690 152504 455696 152516
rect 445536 152476 455696 152504
rect 445536 152464 445542 152476
rect 455690 152464 455696 152476
rect 455748 152464 455754 152516
rect 436370 152436 436376 152448
rect 436112 152408 436376 152436
rect 436370 152396 436376 152408
rect 436428 152396 436434 152448
rect 437474 152396 437480 152448
rect 437532 152436 437538 152448
rect 444466 152436 444472 152448
rect 437532 152408 444472 152436
rect 437532 152396 437538 152408
rect 444466 152396 444472 152408
rect 444524 152396 444530 152448
rect 453758 152436 453764 152448
rect 444944 152408 453764 152436
rect 438302 152368 438308 152380
rect 425204 152340 428228 152368
rect 429948 152340 438308 152368
rect 425204 152328 425210 152340
rect 56502 152260 56508 152312
rect 56560 152300 56566 152312
rect 141050 152300 141056 152312
rect 56560 152272 141056 152300
rect 56560 152260 56566 152272
rect 141050 152260 141056 152272
rect 141108 152260 141114 152312
rect 141142 152260 141148 152312
rect 141200 152300 141206 152312
rect 146938 152300 146944 152312
rect 141200 152272 146944 152300
rect 141200 152260 141206 152272
rect 146938 152260 146944 152272
rect 146996 152260 147002 152312
rect 150434 152260 150440 152312
rect 150492 152300 150498 152312
rect 167362 152300 167368 152312
rect 150492 152272 167368 152300
rect 150492 152260 150498 152272
rect 167362 152260 167368 152272
rect 167420 152260 167426 152312
rect 172606 152260 172612 152312
rect 172664 152300 172670 152312
rect 249518 152300 249524 152312
rect 172664 152272 249524 152300
rect 172664 152260 172670 152272
rect 249518 152260 249524 152272
rect 249576 152260 249582 152312
rect 255498 152260 255504 152312
rect 255556 152300 255562 152312
rect 313090 152300 313096 152312
rect 255556 152272 313096 152300
rect 255556 152260 255562 152272
rect 313090 152260 313096 152272
rect 313148 152260 313154 152312
rect 320266 152260 320272 152312
rect 320324 152300 320330 152312
rect 323118 152300 323124 152312
rect 320324 152272 323124 152300
rect 320324 152260 320330 152272
rect 323118 152260 323124 152272
rect 323176 152260 323182 152312
rect 361298 152300 361304 152312
rect 323228 152272 361304 152300
rect 76926 152192 76932 152244
rect 76984 152232 76990 152244
rect 159634 152232 159640 152244
rect 76984 152204 159640 152232
rect 76984 152192 76990 152204
rect 159634 152192 159640 152204
rect 159692 152192 159698 152244
rect 160186 152192 160192 152244
rect 160244 152232 160250 152244
rect 177666 152232 177672 152244
rect 160244 152204 177672 152232
rect 160244 152192 160250 152204
rect 177666 152192 177672 152204
rect 177724 152192 177730 152244
rect 187970 152192 187976 152244
rect 188028 152232 188034 152244
rect 262398 152232 262404 152244
rect 188028 152204 262404 152232
rect 188028 152192 188034 152204
rect 262398 152192 262404 152204
rect 262456 152192 262462 152244
rect 266354 152192 266360 152244
rect 266412 152232 266418 152244
rect 320818 152232 320824 152244
rect 266412 152204 320824 152232
rect 266412 152192 266418 152204
rect 320818 152192 320824 152204
rect 320876 152192 320882 152244
rect 320910 152192 320916 152244
rect 320968 152232 320974 152244
rect 323228 152232 323256 152272
rect 361298 152260 361304 152272
rect 361356 152260 361362 152312
rect 364518 152260 364524 152312
rect 364576 152300 364582 152312
rect 369026 152300 369032 152312
rect 364576 152272 369032 152300
rect 364576 152260 364582 152272
rect 369026 152260 369032 152272
rect 369084 152260 369090 152312
rect 398466 152300 398472 152312
rect 369136 152272 398472 152300
rect 320968 152204 323256 152232
rect 320968 152192 320974 152204
rect 324314 152192 324320 152244
rect 324372 152232 324378 152244
rect 367002 152232 367008 152244
rect 324372 152204 367008 152232
rect 324372 152192 324378 152204
rect 367002 152192 367008 152204
rect 367060 152192 367066 152244
rect 367094 152192 367100 152244
rect 367152 152232 367158 152244
rect 369136 152232 369164 152272
rect 398466 152260 398472 152272
rect 398524 152260 398530 152312
rect 398558 152260 398564 152312
rect 398616 152300 398622 152312
rect 408126 152300 408132 152312
rect 398616 152272 408132 152300
rect 398616 152260 398622 152272
rect 408126 152260 408132 152272
rect 408184 152260 408190 152312
rect 410886 152260 410892 152312
rect 410944 152300 410950 152312
rect 428200 152300 428228 152340
rect 438302 152328 438308 152340
rect 438360 152328 438366 152380
rect 438394 152328 438400 152380
rect 438452 152368 438458 152380
rect 444944 152368 444972 152408
rect 453758 152396 453764 152408
rect 453816 152396 453822 152448
rect 438452 152340 444972 152368
rect 438452 152328 438458 152340
rect 445110 152328 445116 152380
rect 445168 152368 445174 152380
rect 456334 152368 456340 152380
rect 445168 152340 456340 152368
rect 445168 152328 445174 152340
rect 456334 152328 456340 152340
rect 456392 152328 456398 152380
rect 432690 152300 432696 152312
rect 410944 152272 428044 152300
rect 428200 152272 432696 152300
rect 410944 152260 410950 152272
rect 367152 152204 369164 152232
rect 367152 152192 367158 152204
rect 371326 152192 371332 152244
rect 371384 152232 371390 152244
rect 402330 152232 402336 152244
rect 371384 152204 402336 152232
rect 371384 152192 371390 152204
rect 402330 152192 402336 152204
rect 402388 152192 402394 152244
rect 405826 152192 405832 152244
rect 405884 152232 405890 152244
rect 408770 152232 408776 152244
rect 405884 152204 408776 152232
rect 405884 152192 405890 152204
rect 408770 152192 408776 152204
rect 408828 152192 408834 152244
rect 409230 152192 409236 152244
rect 409288 152232 409294 152244
rect 426710 152232 426716 152244
rect 409288 152204 426716 152232
rect 409288 152192 409294 152204
rect 426710 152192 426716 152204
rect 426768 152192 426774 152244
rect 84746 152124 84752 152176
rect 84804 152164 84810 152176
rect 164786 152164 164792 152176
rect 84804 152136 164792 152164
rect 84804 152124 84810 152136
rect 164786 152124 164792 152136
rect 164844 152124 164850 152176
rect 166994 152124 167000 152176
rect 167052 152164 167058 152176
rect 182726 152164 182732 152176
rect 167052 152136 182732 152164
rect 167052 152124 167058 152136
rect 182726 152124 182732 152136
rect 182784 152124 182790 152176
rect 192662 152124 192668 152176
rect 192720 152164 192726 152176
rect 213546 152164 213552 152176
rect 192720 152136 213552 152164
rect 192720 152124 192726 152136
rect 213546 152124 213552 152136
rect 213604 152124 213610 152176
rect 213822 152124 213828 152176
rect 213880 152164 213886 152176
rect 274542 152164 274548 152176
rect 213880 152136 274548 152164
rect 213880 152124 213886 152136
rect 274542 152124 274548 152136
rect 274600 152124 274606 152176
rect 278774 152124 278780 152176
rect 278832 152164 278838 152176
rect 331766 152164 331772 152176
rect 278832 152136 331772 152164
rect 278832 152124 278838 152136
rect 331766 152124 331772 152136
rect 331824 152124 331830 152176
rect 335814 152124 335820 152176
rect 335872 152164 335878 152176
rect 336826 152164 336832 152176
rect 335872 152136 336832 152164
rect 335872 152124 335878 152136
rect 336826 152124 336832 152136
rect 336884 152124 336890 152176
rect 336918 152124 336924 152176
rect 336976 152164 336982 152176
rect 372798 152164 372804 152176
rect 336976 152136 372804 152164
rect 336976 152124 336982 152136
rect 372798 152124 372804 152136
rect 372856 152124 372862 152176
rect 384942 152124 384948 152176
rect 385000 152164 385006 152176
rect 392118 152164 392124 152176
rect 385000 152136 392124 152164
rect 385000 152124 385006 152136
rect 392118 152124 392124 152136
rect 392176 152124 392182 152176
rect 394326 152124 394332 152176
rect 394384 152164 394390 152176
rect 417786 152164 417792 152176
rect 394384 152136 417792 152164
rect 394384 152124 394390 152136
rect 417786 152124 417792 152136
rect 417844 152124 417850 152176
rect 419626 152124 419632 152176
rect 419684 152164 419690 152176
rect 427722 152164 427728 152176
rect 419684 152136 427728 152164
rect 419684 152124 419690 152136
rect 427722 152124 427728 152136
rect 427780 152124 427786 152176
rect 428016 152164 428044 152272
rect 432690 152260 432696 152272
rect 432748 152260 432754 152312
rect 432782 152260 432788 152312
rect 432840 152300 432846 152312
rect 438946 152300 438952 152312
rect 432840 152272 438952 152300
rect 432840 152260 432846 152272
rect 438946 152260 438952 152272
rect 439004 152260 439010 152312
rect 440510 152260 440516 152312
rect 440568 152300 440574 152312
rect 455046 152300 455052 152312
rect 440568 152272 455052 152300
rect 440568 152260 440574 152272
rect 455046 152260 455052 152272
rect 455104 152260 455110 152312
rect 455506 152260 455512 152312
rect 455564 152300 455570 152312
rect 462038 152300 462044 152312
rect 455564 152272 462044 152300
rect 455564 152260 455570 152272
rect 462038 152260 462044 152272
rect 462096 152260 462102 152312
rect 429378 152192 429384 152244
rect 429436 152232 429442 152244
rect 446674 152232 446680 152244
rect 429436 152204 446680 152232
rect 429436 152192 429442 152204
rect 446674 152192 446680 152204
rect 446732 152192 446738 152244
rect 456794 152192 456800 152244
rect 456852 152232 456858 152244
rect 463326 152232 463332 152244
rect 456852 152204 463332 152232
rect 456852 152192 456858 152204
rect 463326 152192 463332 152204
rect 463384 152192 463390 152244
rect 431218 152164 431224 152176
rect 428016 152136 431224 152164
rect 431218 152124 431224 152136
rect 431276 152124 431282 152176
rect 431310 152124 431316 152176
rect 431368 152164 431374 152176
rect 444098 152164 444104 152176
rect 431368 152136 444104 152164
rect 431368 152124 431374 152136
rect 444098 152124 444104 152136
rect 444156 152124 444162 152176
rect 450538 152164 450544 152176
rect 444944 152136 450544 152164
rect 75822 152056 75828 152108
rect 75880 152096 75886 152108
rect 154482 152096 154488 152108
rect 75880 152068 154488 152096
rect 75880 152056 75886 152068
rect 154482 152056 154488 152068
rect 154540 152056 154546 152108
rect 156046 152056 156052 152108
rect 156104 152096 156110 152108
rect 172514 152096 172520 152108
rect 156104 152068 172520 152096
rect 156104 152056 156110 152068
rect 172514 152056 172520 152068
rect 172572 152056 172578 152108
rect 185578 152056 185584 152108
rect 185636 152096 185642 152108
rect 200758 152096 200764 152108
rect 185636 152068 200764 152096
rect 185636 152056 185642 152068
rect 200758 152056 200764 152068
rect 200816 152056 200822 152108
rect 272702 152096 272708 152108
rect 219406 152068 272708 152096
rect 71774 151988 71780 152040
rect 71832 152028 71838 152040
rect 149422 152028 149428 152040
rect 71832 152000 149428 152028
rect 71832 151988 71838 152000
rect 149422 151988 149428 152000
rect 149480 151988 149486 152040
rect 169754 151988 169760 152040
rect 169812 152028 169818 152040
rect 185302 152028 185308 152040
rect 169812 152000 185308 152028
rect 169812 151988 169818 152000
rect 185302 151988 185308 152000
rect 185360 151988 185366 152040
rect 195146 151988 195152 152040
rect 195204 152028 195210 152040
rect 218698 152028 218704 152040
rect 195204 152000 218704 152028
rect 195204 151988 195210 152000
rect 218698 151988 218704 152000
rect 218756 151988 218762 152040
rect 109034 151920 109040 151972
rect 109092 151960 109098 151972
rect 128170 151960 128176 151972
rect 109092 151932 128176 151960
rect 109092 151920 109098 151932
rect 128170 151920 128176 151932
rect 128228 151920 128234 151972
rect 128354 151920 128360 151972
rect 128412 151960 128418 151972
rect 203334 151960 203340 151972
rect 128412 151932 203340 151960
rect 128412 151920 128418 151932
rect 203334 151920 203340 151932
rect 203392 151920 203398 151972
rect 212718 151920 212724 151972
rect 212776 151960 212782 151972
rect 219406 151960 219434 152068
rect 272702 152056 272708 152068
rect 272760 152056 272766 152108
rect 272794 152056 272800 152108
rect 272852 152096 272858 152108
rect 325970 152096 325976 152108
rect 272852 152068 325976 152096
rect 272852 152056 272858 152068
rect 325970 152056 325976 152068
rect 326028 152056 326034 152108
rect 335354 152056 335360 152108
rect 335412 152096 335418 152108
rect 375374 152096 375380 152108
rect 335412 152068 375380 152096
rect 335412 152056 335418 152068
rect 375374 152056 375380 152068
rect 375432 152056 375438 152108
rect 382274 152056 382280 152108
rect 382332 152096 382338 152108
rect 386966 152096 386972 152108
rect 382332 152068 386972 152096
rect 382332 152056 382338 152068
rect 386966 152056 386972 152068
rect 387024 152056 387030 152108
rect 388346 152056 388352 152108
rect 388404 152096 388410 152108
rect 407482 152096 407488 152108
rect 388404 152068 407488 152096
rect 388404 152056 388410 152068
rect 407482 152056 407488 152068
rect 407540 152056 407546 152108
rect 408494 152056 408500 152108
rect 408552 152096 408558 152108
rect 423582 152096 423588 152108
rect 408552 152068 423588 152096
rect 408552 152056 408558 152068
rect 423582 152056 423588 152068
rect 423640 152056 423646 152108
rect 423674 152056 423680 152108
rect 423732 152096 423738 152108
rect 426342 152096 426348 152108
rect 423732 152068 426348 152096
rect 423732 152056 423738 152068
rect 426342 152056 426348 152068
rect 426400 152056 426406 152108
rect 432414 152056 432420 152108
rect 432472 152096 432478 152108
rect 444742 152096 444748 152108
rect 432472 152068 444748 152096
rect 432472 152056 432478 152068
rect 444742 152056 444748 152068
rect 444800 152056 444806 152108
rect 242802 151988 242808 152040
rect 242860 152028 242866 152040
rect 300946 152028 300952 152040
rect 242860 152000 300952 152028
rect 242860 151988 242866 152000
rect 300946 151988 300952 152000
rect 301004 151988 301010 152040
rect 301038 151988 301044 152040
rect 301096 152028 301102 152040
rect 335998 152028 336004 152040
rect 301096 152000 336004 152028
rect 301096 151988 301102 152000
rect 335998 151988 336004 152000
rect 336056 151988 336062 152040
rect 338086 152000 340874 152028
rect 212776 151932 219434 151960
rect 212776 151920 212782 151932
rect 243354 151920 243360 151972
rect 243412 151960 243418 151972
rect 302878 151960 302884 151972
rect 243412 151932 302884 151960
rect 243412 151920 243418 151932
rect 302878 151920 302884 151932
rect 302936 151920 302942 151972
rect 317414 151920 317420 151972
rect 317472 151960 317478 151972
rect 320910 151960 320916 151972
rect 317472 151932 320916 151960
rect 317472 151920 317478 151932
rect 320910 151920 320916 151932
rect 320968 151920 320974 151972
rect 321554 151920 321560 151972
rect 321612 151960 321618 151972
rect 325602 151960 325608 151972
rect 321612 151932 325608 151960
rect 321612 151920 321618 151932
rect 325602 151920 325608 151932
rect 325660 151920 325666 151972
rect 325878 151920 325884 151972
rect 325936 151960 325942 151972
rect 338086 151960 338114 152000
rect 325936 151932 338114 151960
rect 340846 151960 340874 152000
rect 342438 151988 342444 152040
rect 342496 152028 342502 152040
rect 344554 152028 344560 152040
rect 342496 152000 344560 152028
rect 342496 151988 342502 152000
rect 344554 151988 344560 152000
rect 344612 151988 344618 152040
rect 354674 151988 354680 152040
rect 354732 152028 354738 152040
rect 359458 152028 359464 152040
rect 354732 152000 359464 152028
rect 354732 151988 354738 152000
rect 359458 151988 359464 152000
rect 359516 151988 359522 152040
rect 378778 151988 378784 152040
rect 378836 152028 378842 152040
rect 384390 152028 384396 152040
rect 378836 152000 384396 152028
rect 378836 151988 378842 152000
rect 384390 151988 384396 152000
rect 384448 151988 384454 152040
rect 385770 151988 385776 152040
rect 385828 152028 385834 152040
rect 394694 152028 394700 152040
rect 385828 152000 394700 152028
rect 385828 151988 385834 152000
rect 394694 151988 394700 152000
rect 394752 151988 394758 152040
rect 404722 151988 404728 152040
rect 404780 152028 404786 152040
rect 421006 152028 421012 152040
rect 404780 152000 421012 152028
rect 404780 151988 404786 152000
rect 421006 151988 421012 152000
rect 421064 151988 421070 152040
rect 426802 152028 426808 152040
rect 422266 152000 426808 152028
rect 367646 151960 367652 151972
rect 340846 151932 367652 151960
rect 325936 151920 325942 151932
rect 367646 151920 367652 151932
rect 367704 151920 367710 151972
rect 375466 151920 375472 151972
rect 375524 151960 375530 151972
rect 405550 151960 405556 151972
rect 375524 151932 405556 151960
rect 375524 151920 375530 151932
rect 405550 151920 405556 151932
rect 405608 151920 405614 151972
rect 416590 151920 416596 151972
rect 416648 151960 416654 151972
rect 422266 151960 422294 152000
rect 426802 151988 426808 152000
rect 426860 151988 426866 152040
rect 432690 151988 432696 152040
rect 432748 152028 432754 152040
rect 443454 152028 443460 152040
rect 432748 152000 443460 152028
rect 432748 151988 432754 152000
rect 443454 151988 443460 152000
rect 443512 151988 443518 152040
rect 443546 151988 443552 152040
rect 443604 152028 443610 152040
rect 444944 152028 444972 152136
rect 450538 152124 450544 152136
rect 450596 152124 450602 152176
rect 455874 152124 455880 152176
rect 455932 152164 455938 152176
rect 461394 152164 461400 152176
rect 455932 152136 461400 152164
rect 455932 152124 455938 152136
rect 461394 152124 461400 152136
rect 461452 152124 461458 152176
rect 446306 152056 446312 152108
rect 446364 152096 446370 152108
rect 460106 152096 460112 152108
rect 446364 152068 460112 152096
rect 446364 152056 446370 152068
rect 460106 152056 460112 152068
rect 460164 152056 460170 152108
rect 443604 152000 444972 152028
rect 443604 151988 443610 152000
rect 445294 151988 445300 152040
rect 445352 152028 445358 152040
rect 458818 152028 458824 152040
rect 445352 152000 458824 152028
rect 445352 151988 445358 152000
rect 458818 151988 458824 152000
rect 458876 151988 458882 152040
rect 485774 151988 485780 152040
rect 485832 152028 485838 152040
rect 490282 152028 490288 152040
rect 485832 152000 490288 152028
rect 485832 151988 485838 152000
rect 490282 151988 490288 152000
rect 490340 151988 490346 152040
rect 516686 151988 516692 152040
rect 516744 152028 516750 152040
rect 520274 152028 520280 152040
rect 516744 152000 520280 152028
rect 516744 151988 516750 152000
rect 520274 151988 520280 152000
rect 520332 151988 520338 152040
rect 416648 151932 422294 151960
rect 416648 151920 416654 151932
rect 422570 151920 422576 151972
rect 422628 151960 422634 151972
rect 429838 151960 429844 151972
rect 422628 151932 429844 151960
rect 422628 151920 422634 151932
rect 429838 151920 429844 151932
rect 429896 151920 429902 151972
rect 434530 151920 434536 151972
rect 434588 151960 434594 151972
rect 439590 151960 439596 151972
rect 434588 151932 439596 151960
rect 434588 151920 434594 151932
rect 439590 151920 439596 151932
rect 439648 151920 439654 151972
rect 440234 151920 440240 151972
rect 440292 151960 440298 151972
rect 451090 151960 451096 151972
rect 440292 151932 451096 151960
rect 440292 151920 440298 151932
rect 451090 151920 451096 151932
rect 451148 151920 451154 151972
rect 451182 151920 451188 151972
rect 451240 151960 451246 151972
rect 457622 151960 457628 151972
rect 451240 151932 457628 151960
rect 451240 151920 451246 151932
rect 457622 151920 457628 151932
rect 457680 151920 457686 151972
rect 469214 151920 469220 151972
rect 469272 151960 469278 151972
rect 472342 151960 472348 151972
rect 469272 151932 472348 151960
rect 469272 151920 469278 151932
rect 472342 151920 472348 151932
rect 472400 151920 472406 151972
rect 487338 151920 487344 151972
rect 487396 151960 487402 151972
rect 490926 151960 490932 151972
rect 487396 151932 490932 151960
rect 487396 151920 487402 151932
rect 490926 151920 490932 151932
rect 490984 151920 490990 151972
rect 509050 151920 509056 151972
rect 509108 151960 509114 151972
rect 510890 151960 510896 151972
rect 509108 151932 510896 151960
rect 509108 151920 509114 151932
rect 510890 151920 510896 151932
rect 510948 151920 510954 151972
rect 515490 151920 515496 151972
rect 515548 151960 515554 151972
rect 518986 151960 518992 151972
rect 515548 151932 518992 151960
rect 515548 151920 515554 151932
rect 518986 151920 518992 151932
rect 519044 151920 519050 151972
rect 30190 151852 30196 151904
rect 30248 151892 30254 151904
rect 74534 151892 74540 151904
rect 30248 151864 74540 151892
rect 30248 151852 30254 151864
rect 74534 151852 74540 151864
rect 74592 151852 74598 151904
rect 107562 151852 107568 151904
rect 107620 151892 107626 151904
rect 175090 151892 175096 151904
rect 107620 151864 175096 151892
rect 107620 151852 107626 151864
rect 175090 151852 175096 151864
rect 175148 151852 175154 151904
rect 176654 151852 176660 151904
rect 176712 151892 176718 151904
rect 190454 151892 190460 151904
rect 176712 151864 190460 151892
rect 176712 151852 176718 151864
rect 190454 151852 190460 151864
rect 190512 151852 190518 151904
rect 261018 151852 261024 151904
rect 261076 151892 261082 151904
rect 316310 151892 316316 151904
rect 261076 151864 316316 151892
rect 261076 151852 261082 151864
rect 316310 151852 316316 151864
rect 316368 151852 316374 151904
rect 320726 151852 320732 151904
rect 320784 151892 320790 151904
rect 326614 151892 326620 151904
rect 320784 151864 326620 151892
rect 320784 151852 320790 151864
rect 326614 151852 326620 151864
rect 326672 151852 326678 151904
rect 331122 151892 331128 151904
rect 328288 151864 331128 151892
rect 33594 151784 33600 151836
rect 33652 151824 33658 151836
rect 84194 151824 84200 151836
rect 33652 151796 84200 151824
rect 33652 151784 33658 151796
rect 84194 151784 84200 151796
rect 84252 151784 84258 151836
rect 105814 151784 105820 151836
rect 105872 151824 105878 151836
rect 109770 151824 109776 151836
rect 105872 151796 109776 151824
rect 105872 151784 105878 151796
rect 109770 151784 109776 151796
rect 109828 151784 109834 151836
rect 109862 151784 109868 151836
rect 109920 151824 109926 151836
rect 138474 151824 138480 151836
rect 109920 151796 138480 151824
rect 109920 151784 109926 151796
rect 138474 151784 138480 151796
rect 138532 151784 138538 151836
rect 138566 151784 138572 151836
rect 138624 151824 138630 151836
rect 141878 151824 141884 151836
rect 138624 151796 141884 151824
rect 138624 151784 138630 151796
rect 141878 151784 141884 151796
rect 141936 151784 141942 151836
rect 142246 151784 142252 151836
rect 142304 151824 142310 151836
rect 157058 151824 157064 151836
rect 142304 151796 157064 151824
rect 142304 151784 142310 151796
rect 157058 151784 157064 151796
rect 157116 151784 157122 151836
rect 183094 151784 183100 151836
rect 183152 151824 183158 151836
rect 195606 151824 195612 151836
rect 183152 151796 195612 151824
rect 183152 151784 183158 151796
rect 195606 151784 195612 151796
rect 195664 151784 195670 151836
rect 277394 151784 277400 151836
rect 277452 151824 277458 151836
rect 328288 151824 328316 151864
rect 331122 151852 331128 151864
rect 331180 151852 331186 151904
rect 332594 151852 332600 151904
rect 332652 151892 332658 151904
rect 336918 151892 336924 151904
rect 332652 151864 336924 151892
rect 332652 151852 332658 151864
rect 336918 151852 336924 151864
rect 336976 151852 336982 151904
rect 337010 151852 337016 151904
rect 337068 151892 337074 151904
rect 372154 151892 372160 151904
rect 337068 151864 372160 151892
rect 337068 151852 337074 151864
rect 372154 151852 372160 151864
rect 372212 151852 372218 151904
rect 396166 151852 396172 151904
rect 396224 151892 396230 151904
rect 402974 151892 402980 151904
rect 396224 151864 402980 151892
rect 396224 151852 396230 151864
rect 402974 151852 402980 151864
rect 403032 151852 403038 151904
rect 404262 151852 404268 151904
rect 404320 151892 404326 151904
rect 418430 151892 418436 151904
rect 404320 151864 418436 151892
rect 404320 151852 404326 151864
rect 418430 151852 418436 151864
rect 418488 151852 418494 151904
rect 419534 151852 419540 151904
rect 419592 151892 419598 151904
rect 437014 151892 437020 151904
rect 419592 151864 437020 151892
rect 419592 151852 419598 151864
rect 437014 151852 437020 151864
rect 437072 151852 437078 151904
rect 437106 151852 437112 151904
rect 437164 151892 437170 151904
rect 442166 151892 442172 151904
rect 437164 151864 442172 151892
rect 437164 151852 437170 151864
rect 442166 151852 442172 151864
rect 442224 151852 442230 151904
rect 442258 151852 442264 151904
rect 442316 151892 442322 151904
rect 442316 151864 444788 151892
rect 442316 151852 442322 151864
rect 362586 151824 362592 151836
rect 277452 151796 328316 151824
rect 328426 151796 362592 151824
rect 277452 151784 277458 151796
rect 325602 151716 325608 151768
rect 325660 151756 325666 151768
rect 328426 151756 328454 151796
rect 362586 151784 362592 151796
rect 362644 151784 362650 151836
rect 363138 151784 363144 151836
rect 363196 151824 363202 151836
rect 364518 151824 364524 151836
rect 363196 151796 364524 151824
rect 363196 151784 363202 151796
rect 364518 151784 364524 151796
rect 364576 151784 364582 151836
rect 388438 151784 388444 151836
rect 388496 151824 388502 151836
rect 404906 151824 404912 151836
rect 388496 151796 404912 151824
rect 388496 151784 388502 151796
rect 404906 151784 404912 151796
rect 404964 151784 404970 151836
rect 417418 151784 417424 151836
rect 417476 151824 417482 151836
rect 431862 151824 431868 151836
rect 417476 151796 427814 151824
rect 417476 151784 417482 151796
rect 325660 151728 328454 151756
rect 325660 151716 325666 151728
rect 427786 151688 427814 151796
rect 428200 151796 431868 151824
rect 428200 151688 428228 151796
rect 431862 151784 431868 151796
rect 431920 151784 431926 151836
rect 432598 151784 432604 151836
rect 432656 151824 432662 151836
rect 440878 151824 440884 151836
rect 432656 151796 440884 151824
rect 432656 151784 432662 151796
rect 440878 151784 440884 151796
rect 440936 151784 440942 151836
rect 441430 151784 441436 151836
rect 441488 151824 441494 151836
rect 444760 151824 444788 151864
rect 444834 151852 444840 151904
rect 444892 151892 444898 151904
rect 452470 151892 452476 151904
rect 444892 151864 452476 151892
rect 444892 151852 444898 151864
rect 452470 151852 452476 151864
rect 452528 151852 452534 151904
rect 467834 151852 467840 151904
rect 467892 151892 467898 151904
rect 471054 151892 471060 151904
rect 467892 151864 471060 151892
rect 467892 151852 467898 151864
rect 471054 151852 471060 151864
rect 471112 151852 471118 151904
rect 488534 151852 488540 151904
rect 488592 151892 488598 151904
rect 492214 151892 492220 151904
rect 488592 151864 492220 151892
rect 488592 151852 488598 151864
rect 492214 151852 492220 151864
rect 492272 151852 492278 151904
rect 507762 151852 507768 151904
rect 507820 151892 507826 151904
rect 509510 151892 509516 151904
rect 507820 151864 509516 151892
rect 507820 151852 507826 151864
rect 509510 151852 509516 151864
rect 509568 151852 509574 151904
rect 516042 151852 516048 151904
rect 516100 151892 516106 151904
rect 519906 151892 519912 151904
rect 516100 151864 519912 151892
rect 516100 151852 516106 151864
rect 519906 151852 519912 151864
rect 519964 151852 519970 151904
rect 451826 151824 451832 151836
rect 441488 151796 444696 151824
rect 444760 151796 451832 151824
rect 441488 151784 441494 151796
rect 427786 151660 428228 151688
rect 444668 151688 444696 151796
rect 451826 151784 451832 151796
rect 451884 151784 451890 151836
rect 457162 151784 457168 151836
rect 457220 151824 457226 151836
rect 462682 151824 462688 151836
rect 457220 151796 462688 151824
rect 457220 151784 457226 151796
rect 462682 151784 462688 151796
rect 462740 151784 462746 151836
rect 464338 151784 464344 151836
rect 464396 151824 464402 151836
rect 467742 151824 467748 151836
rect 464396 151796 467748 151824
rect 464396 151784 464402 151796
rect 467742 151784 467748 151796
rect 467800 151784 467806 151836
rect 467926 151784 467932 151836
rect 467984 151824 467990 151836
rect 471698 151824 471704 151836
rect 467984 151796 471704 151824
rect 467984 151784 467990 151796
rect 471698 151784 471704 151796
rect 471756 151784 471762 151836
rect 488166 151784 488172 151836
rect 488224 151824 488230 151836
rect 491570 151824 491576 151836
rect 488224 151796 491576 151824
rect 488224 151784 488230 151796
rect 491570 151784 491576 151796
rect 491628 151784 491634 151836
rect 499114 151784 499120 151836
rect 499172 151824 499178 151836
rect 499942 151824 499948 151836
rect 499172 151796 499948 151824
rect 499172 151784 499178 151796
rect 499942 151784 499948 151796
rect 500000 151784 500006 151836
rect 517422 151784 517428 151836
rect 517480 151824 517486 151836
rect 521562 151824 521568 151836
rect 517480 151796 521568 151824
rect 517480 151784 517486 151796
rect 521562 151784 521568 151796
rect 521620 151784 521626 151836
rect 446030 151688 446036 151700
rect 444668 151660 446036 151688
rect 446030 151648 446036 151660
rect 446088 151648 446094 151700
rect 84194 151376 84200 151428
rect 84252 151416 84258 151428
rect 117222 151416 117228 151428
rect 84252 151388 117228 151416
rect 84252 151376 84258 151388
rect 117222 151376 117228 151388
rect 117280 151376 117286 151428
rect 74534 151308 74540 151360
rect 74592 151348 74598 151360
rect 117130 151348 117136 151360
rect 74592 151320 117136 151348
rect 74592 151308 74598 151320
rect 117130 151308 117136 151320
rect 117188 151308 117194 151360
rect 68002 151240 68008 151292
rect 68060 151280 68066 151292
rect 112806 151280 112812 151292
rect 68060 151252 112812 151280
rect 68060 151240 68066 151252
rect 112806 151240 112812 151252
rect 112864 151240 112870 151292
rect 64506 151172 64512 151224
rect 64564 151212 64570 151224
rect 112714 151212 112720 151224
rect 64564 151184 112720 151212
rect 64564 151172 64570 151184
rect 112714 151172 112720 151184
rect 112772 151172 112778 151224
rect 61102 151104 61108 151156
rect 61160 151144 61166 151156
rect 112622 151144 112628 151156
rect 61160 151116 112628 151144
rect 61160 151104 61166 151116
rect 112622 151104 112628 151116
rect 112680 151104 112686 151156
rect 57698 151036 57704 151088
rect 57756 151076 57762 151088
rect 112530 151076 112536 151088
rect 57756 151048 112536 151076
rect 57756 151036 57762 151048
rect 112530 151036 112536 151048
rect 112588 151036 112594 151088
rect 54202 150968 54208 151020
rect 54260 151008 54266 151020
rect 111610 151008 111616 151020
rect 54260 150980 111616 151008
rect 54260 150968 54266 150980
rect 111610 150968 111616 150980
rect 111668 150968 111674 151020
rect 50798 150900 50804 150952
rect 50856 150940 50862 150952
rect 112438 150940 112444 150952
rect 50856 150912 112444 150940
rect 50856 150900 50862 150912
rect 112438 150900 112444 150912
rect 112496 150900 112502 150952
rect 47302 150832 47308 150884
rect 47360 150872 47366 150884
rect 111518 150872 111524 150884
rect 47360 150844 111524 150872
rect 47360 150832 47366 150844
rect 111518 150832 111524 150844
rect 111576 150832 111582 150884
rect 43898 150764 43904 150816
rect 43956 150804 43962 150816
rect 111426 150804 111432 150816
rect 43956 150776 111432 150804
rect 43956 150764 43962 150776
rect 111426 150764 111432 150776
rect 111484 150764 111490 150816
rect 40494 150696 40500 150748
rect 40552 150736 40558 150748
rect 111334 150736 111340 150748
rect 40552 150708 111340 150736
rect 40552 150696 40558 150708
rect 111334 150696 111340 150708
rect 111392 150696 111398 150748
rect 36998 150628 37004 150680
rect 37056 150668 37062 150680
rect 111242 150668 111248 150680
rect 37056 150640 111248 150668
rect 37056 150628 37062 150640
rect 111242 150628 111248 150640
rect 111300 150628 111306 150680
rect 19794 150560 19800 150612
rect 19852 150600 19858 150612
rect 116854 150600 116860 150612
rect 19852 150572 116860 150600
rect 19852 150560 19858 150572
rect 116854 150560 116860 150572
rect 116912 150560 116918 150612
rect 16390 150492 16396 150544
rect 16448 150532 16454 150544
rect 116762 150532 116768 150544
rect 16448 150504 116768 150532
rect 16448 150492 16454 150504
rect 116762 150492 116768 150504
rect 116820 150492 116826 150544
rect 2682 150424 2688 150476
rect 2740 150464 2746 150476
rect 111058 150464 111064 150476
rect 2740 150436 111064 150464
rect 2740 150424 2746 150436
rect 111058 150424 111064 150436
rect 111116 150424 111122 150476
rect 263686 150288 263692 150340
rect 263744 150328 263750 150340
rect 263744 150300 264422 150328
rect 263744 150288 263750 150300
rect 264394 150204 264422 150300
rect 122834 150152 122840 150204
rect 122892 150192 122898 150204
rect 123708 150192 123714 150204
rect 122892 150164 123714 150192
rect 122892 150152 122898 150164
rect 123708 150152 123714 150164
rect 123766 150152 123772 150204
rect 146386 150152 146392 150204
rect 146444 150192 146450 150204
rect 147536 150192 147542 150204
rect 146444 150164 147542 150192
rect 146444 150152 146450 150164
rect 147536 150152 147542 150164
rect 147594 150152 147600 150204
rect 147674 150152 147680 150204
rect 147732 150192 147738 150204
rect 148824 150192 148830 150204
rect 147732 150164 148830 150192
rect 147732 150152 147738 150164
rect 148824 150152 148830 150164
rect 148882 150152 148888 150204
rect 165706 150152 165712 150204
rect 165764 150192 165770 150204
rect 166764 150192 166770 150204
rect 165764 150164 166770 150192
rect 165764 150152 165770 150164
rect 166764 150152 166770 150164
rect 166822 150152 166828 150204
rect 171134 150152 171140 150204
rect 171192 150192 171198 150204
rect 171916 150192 171922 150204
rect 171192 150164 171922 150192
rect 171192 150152 171198 150164
rect 171916 150152 171922 150164
rect 171974 150152 171980 150204
rect 172698 150152 172704 150204
rect 172756 150192 172762 150204
rect 173848 150192 173854 150204
rect 172756 150164 173854 150192
rect 172756 150152 172762 150164
rect 173848 150152 173854 150164
rect 173906 150152 173912 150204
rect 182266 150152 182272 150204
rect 182324 150192 182330 150204
rect 183416 150192 183422 150204
rect 182324 150164 183422 150192
rect 182324 150152 182330 150164
rect 183416 150152 183422 150164
rect 183474 150152 183480 150204
rect 183554 150152 183560 150204
rect 183612 150192 183618 150204
rect 184704 150192 184710 150204
rect 183612 150164 184710 150192
rect 183612 150152 183618 150164
rect 184704 150152 184710 150164
rect 184762 150152 184768 150204
rect 200298 150152 200304 150204
rect 200356 150192 200362 150204
rect 201448 150192 201454 150204
rect 200356 150164 201454 150192
rect 200356 150152 200362 150164
rect 201448 150152 201454 150164
rect 201506 150152 201512 150204
rect 219526 150152 219532 150204
rect 219584 150192 219590 150204
rect 220676 150192 220682 150204
rect 219584 150164 220682 150192
rect 219584 150152 219590 150164
rect 220676 150152 220682 150164
rect 220734 150152 220740 150204
rect 222286 150152 222292 150204
rect 222344 150192 222350 150204
rect 223252 150192 223258 150204
rect 222344 150164 223258 150192
rect 222344 150152 222350 150164
rect 223252 150152 223258 150164
rect 223310 150152 223316 150204
rect 229186 150152 229192 150204
rect 229244 150192 229250 150204
rect 230336 150192 230342 150204
rect 229244 150164 230342 150192
rect 229244 150152 229250 150164
rect 230336 150152 230342 150164
rect 230394 150152 230400 150204
rect 238938 150152 238944 150204
rect 238996 150192 239002 150204
rect 239996 150192 240002 150204
rect 238996 150164 240002 150192
rect 238996 150152 239002 150164
rect 239996 150152 240002 150164
rect 240054 150152 240060 150204
rect 253934 150152 253940 150204
rect 253992 150192 253998 150204
rect 254716 150192 254722 150204
rect 253992 150164 254722 150192
rect 253992 150152 253998 150164
rect 254716 150152 254722 150164
rect 254774 150152 254780 150204
rect 256786 150152 256792 150204
rect 256844 150192 256850 150204
rect 257936 150192 257942 150204
rect 256844 150164 257942 150192
rect 256844 150152 256850 150164
rect 257936 150152 257942 150164
rect 257994 150152 258000 150204
rect 258074 150152 258080 150204
rect 258132 150192 258138 150204
rect 259224 150192 259230 150204
rect 258132 150164 259230 150192
rect 258132 150152 258138 150164
rect 259224 150152 259230 150164
rect 259282 150152 259288 150204
rect 264376 150152 264382 150204
rect 264434 150152 264440 150204
rect 269114 150152 269120 150204
rect 269172 150192 269178 150204
rect 270172 150192 270178 150204
rect 269172 150164 270178 150192
rect 269172 150152 269178 150164
rect 270172 150152 270178 150164
rect 270230 150152 270236 150204
rect 281534 150152 281540 150204
rect 281592 150192 281598 150204
rect 282316 150192 282322 150204
rect 281592 150164 282322 150192
rect 281592 150152 281598 150164
rect 282316 150152 282322 150164
rect 282374 150152 282380 150204
rect 283098 150152 283104 150204
rect 283156 150192 283162 150204
rect 284248 150192 284254 150204
rect 283156 150164 284254 150192
rect 283156 150152 283162 150164
rect 284248 150152 284254 150164
rect 284306 150152 284312 150204
rect 284386 150152 284392 150204
rect 284444 150192 284450 150204
rect 285536 150192 285542 150204
rect 284444 150164 285542 150192
rect 284444 150152 284450 150164
rect 285536 150152 285542 150164
rect 285594 150152 285600 150204
rect 299474 150152 299480 150204
rect 299532 150192 299538 150204
rect 300348 150192 300354 150204
rect 299532 150164 300354 150192
rect 299532 150152 299538 150164
rect 300348 150152 300354 150164
rect 300406 150152 300412 150204
rect 321738 150152 321744 150204
rect 321796 150192 321802 150204
rect 322796 150192 322802 150204
rect 321796 150164 322802 150192
rect 321796 150152 321802 150164
rect 322796 150152 322802 150164
rect 322854 150152 322860 150204
rect 338390 150152 338396 150204
rect 338448 150192 338454 150204
rect 339448 150192 339454 150204
rect 338448 150164 339454 150192
rect 338448 150152 338454 150164
rect 339448 150152 339454 150164
rect 339506 150152 339512 150204
rect 345106 150152 345112 150204
rect 345164 150192 345170 150204
rect 345888 150192 345894 150204
rect 345164 150164 345894 150192
rect 345164 150152 345170 150164
rect 345888 150152 345894 150164
rect 345946 150152 345952 150204
rect 358906 150152 358912 150204
rect 358964 150192 358970 150204
rect 360056 150192 360062 150204
rect 358964 150164 360062 150192
rect 358964 150152 358970 150164
rect 360056 150152 360062 150164
rect 360114 150152 360120 150204
rect 362954 150152 362960 150204
rect 363012 150192 363018 150204
rect 363920 150192 363926 150204
rect 363012 150164 363926 150192
rect 363012 150152 363018 150164
rect 363920 150152 363926 150164
rect 363978 150152 363984 150204
rect 373994 150152 374000 150204
rect 374052 150192 374058 150204
rect 374776 150192 374782 150204
rect 374052 150164 374782 150192
rect 374052 150152 374058 150164
rect 374776 150152 374782 150164
rect 374834 150152 374840 150204
rect 378134 150152 378140 150204
rect 378192 150192 378198 150204
rect 379284 150192 379290 150204
rect 378192 150164 379290 150192
rect 378192 150152 378198 150164
rect 379284 150152 379290 150164
rect 379342 150152 379348 150204
rect 403158 150152 403164 150204
rect 403216 150192 403222 150204
rect 404308 150192 404314 150204
rect 403216 150164 404314 150192
rect 403216 150152 403222 150164
rect 404308 150152 404314 150164
rect 404366 150152 404372 150204
rect 426710 150152 426716 150204
rect 426768 150192 426774 150204
rect 428688 150192 428694 150204
rect 426768 150164 428694 150192
rect 426768 150152 426774 150164
rect 428688 150152 428694 150164
rect 428746 150152 428752 150204
rect 444466 150152 444472 150204
rect 444524 150192 444530 150204
rect 453160 150192 453166 150204
rect 444524 150164 453166 150192
rect 444524 150152 444530 150164
rect 453160 150152 453166 150164
rect 453218 150152 453224 150204
rect 477678 150152 477684 150204
rect 477736 150192 477742 150204
rect 478828 150192 478834 150204
rect 477736 150164 478834 150192
rect 477736 150152 477742 150164
rect 478828 150152 478834 150164
rect 478886 150152 478892 150204
rect 478966 150152 478972 150204
rect 479024 150192 479030 150204
rect 480116 150192 480122 150204
rect 479024 150164 480122 150192
rect 479024 150152 479030 150164
rect 480116 150152 480122 150164
rect 480174 150152 480180 150204
rect 481634 150152 481640 150204
rect 481692 150192 481698 150204
rect 482692 150192 482698 150204
rect 481692 150164 482698 150192
rect 481692 150152 481698 150164
rect 482692 150152 482698 150164
rect 482750 150152 482756 150204
rect 483198 150152 483204 150204
rect 483256 150192 483262 150204
rect 483980 150192 483986 150204
rect 483256 150164 483986 150192
rect 483256 150152 483262 150164
rect 483980 150152 483986 150164
rect 484038 150152 484044 150204
rect 505278 150152 505284 150204
rect 505336 150192 505342 150204
rect 506428 150192 506434 150204
rect 505336 150164 506434 150192
rect 505336 150152 505342 150164
rect 506428 150152 506434 150164
rect 506486 150152 506492 150204
rect 518020 150152 518026 150204
rect 518078 150192 518084 150204
rect 518802 150192 518808 150204
rect 518078 150164 518808 150192
rect 518078 150152 518084 150164
rect 518802 150152 518808 150164
rect 518860 150152 518866 150204
rect 427722 150084 427728 150136
rect 427780 150124 427786 150136
rect 434484 150124 434490 150136
rect 427780 150096 434490 150124
rect 427780 150084 427786 150096
rect 434484 150084 434490 150096
rect 434542 150084 434548 150136
rect 6362 150016 6368 150068
rect 6420 150056 6426 150068
rect 111150 150056 111156 150068
rect 6420 150028 111156 150056
rect 6420 150016 6426 150028
rect 111150 150016 111156 150028
rect 111208 150016 111214 150068
rect 23382 149948 23388 150000
rect 23440 149988 23446 150000
rect 116946 149988 116952 150000
rect 23440 149960 116952 149988
rect 23440 149948 23446 149960
rect 116946 149948 116952 149960
rect 117004 149948 117010 150000
rect 13354 149880 13360 149932
rect 13412 149920 13418 149932
rect 116670 149920 116676 149932
rect 13412 149892 116676 149920
rect 13412 149880 13418 149892
rect 116670 149880 116676 149892
rect 116728 149880 116734 149932
rect 9582 149812 9588 149864
rect 9640 149852 9646 149864
rect 116578 149852 116584 149864
rect 9640 149824 116584 149852
rect 9640 149812 9646 149824
rect 116578 149812 116584 149824
rect 116636 149812 116642 149864
rect 88978 149744 88984 149796
rect 89036 149784 89042 149796
rect 114002 149784 114008 149796
rect 89036 149756 114008 149784
rect 89036 149744 89042 149756
rect 114002 149744 114008 149756
rect 114060 149744 114066 149796
rect 85482 149676 85488 149728
rect 85540 149716 85546 149728
rect 113910 149716 113916 149728
rect 85540 149688 113916 149716
rect 85540 149676 85546 149688
rect 113910 149676 113916 149688
rect 113968 149676 113974 149728
rect 81986 149608 81992 149660
rect 82044 149648 82050 149660
rect 112346 149648 112352 149660
rect 82044 149620 112352 149648
rect 82044 149608 82050 149620
rect 112346 149608 112352 149620
rect 112404 149608 112410 149660
rect 78582 149540 78588 149592
rect 78640 149580 78646 149592
rect 113082 149580 113088 149592
rect 78640 149552 113088 149580
rect 78640 149540 78646 149552
rect 113082 149540 113088 149552
rect 113140 149540 113146 149592
rect 75178 149472 75184 149524
rect 75236 149512 75242 149524
rect 112990 149512 112996 149524
rect 75236 149484 112996 149512
rect 75236 149472 75242 149484
rect 112990 149472 112996 149484
rect 113048 149472 113054 149524
rect 71682 149404 71688 149456
rect 71740 149444 71746 149456
rect 112898 149444 112904 149456
rect 71740 149416 112904 149444
rect 71740 149404 71746 149416
rect 112898 149404 112904 149416
rect 112956 149404 112962 149456
rect 26970 149336 26976 149388
rect 27028 149376 27034 149388
rect 117038 149376 117044 149388
rect 27028 149348 117044 149376
rect 27028 149336 27034 149348
rect 117038 149336 117044 149348
rect 117096 149336 117102 149388
rect 92290 149268 92296 149320
rect 92348 149308 92354 149320
rect 92348 149280 93854 149308
rect 92348 149268 92354 149280
rect 93826 149104 93854 149280
rect 95786 149268 95792 149320
rect 95844 149268 95850 149320
rect 105262 149268 105268 149320
rect 105320 149308 105326 149320
rect 116210 149308 116216 149320
rect 105320 149280 116216 149308
rect 105320 149268 105326 149280
rect 116210 149268 116216 149280
rect 116268 149268 116274 149320
rect 95804 149240 95832 149268
rect 116486 149240 116492 149252
rect 95804 149212 101628 149240
rect 93826 149076 96614 149104
rect 96586 148696 96614 149076
rect 101600 148764 101628 149212
rect 104866 149212 116492 149240
rect 104866 148968 104894 149212
rect 116486 149200 116492 149212
rect 116544 149200 116550 149252
rect 109678 149132 109684 149184
rect 109736 149172 109742 149184
rect 116026 149172 116032 149184
rect 109736 149144 116032 149172
rect 109736 149132 109742 149144
rect 116026 149132 116032 149144
rect 116084 149132 116090 149184
rect 114094 149104 114100 149116
rect 103532 148940 104894 148968
rect 105372 149076 114100 149104
rect 103532 148764 103560 148940
rect 101600 148736 103560 148764
rect 105372 148696 105400 149076
rect 114094 149064 114100 149076
rect 114152 149064 114158 149116
rect 109586 148996 109592 149048
rect 109644 149036 109650 149048
rect 116118 149036 116124 149048
rect 109644 149008 116124 149036
rect 109644 148996 109650 149008
rect 116118 148996 116124 149008
rect 116176 148996 116182 149048
rect 96586 148668 105400 148696
rect 109770 147568 109776 147620
rect 109828 147608 109834 147620
rect 116118 147608 116124 147620
rect 109828 147580 116124 147608
rect 109828 147568 109834 147580
rect 116118 147568 116124 147580
rect 116176 147568 116182 147620
rect 114094 140700 114100 140752
rect 114152 140740 114158 140752
rect 116394 140740 116400 140752
rect 114152 140712 116400 140740
rect 114152 140700 114158 140712
rect 116394 140700 116400 140712
rect 116452 140700 116458 140752
rect 114002 137912 114008 137964
rect 114060 137952 114066 137964
rect 116210 137952 116216 137964
rect 114060 137924 116216 137952
rect 114060 137912 114066 137924
rect 116210 137912 116216 137924
rect 116268 137912 116274 137964
rect 113910 136552 113916 136604
rect 113968 136592 113974 136604
rect 116394 136592 116400 136604
rect 113968 136564 116400 136592
rect 113968 136552 113974 136564
rect 116394 136552 116400 136564
rect 116452 136552 116458 136604
rect 112346 133832 112352 133884
rect 112404 133872 112410 133884
rect 116118 133872 116124 133884
rect 112404 133844 116124 133872
rect 112404 133832 112410 133844
rect 116118 133832 116124 133844
rect 116176 133832 116182 133884
rect 113082 132404 113088 132456
rect 113140 132444 113146 132456
rect 116118 132444 116124 132456
rect 113140 132416 116124 132444
rect 113140 132404 113146 132416
rect 116118 132404 116124 132416
rect 116176 132404 116182 132456
rect 112990 131044 112996 131096
rect 113048 131084 113054 131096
rect 116118 131084 116124 131096
rect 113048 131056 116124 131084
rect 113048 131044 113054 131056
rect 116118 131044 116124 131056
rect 116176 131044 116182 131096
rect 112898 128256 112904 128308
rect 112956 128296 112962 128308
rect 116118 128296 116124 128308
rect 112956 128268 116124 128296
rect 112956 128256 112962 128268
rect 116118 128256 116124 128268
rect 116176 128256 116182 128308
rect 112806 126896 112812 126948
rect 112864 126936 112870 126948
rect 116118 126936 116124 126948
rect 112864 126908 116124 126936
rect 112864 126896 112870 126908
rect 116118 126896 116124 126908
rect 116176 126896 116182 126948
rect 112714 124108 112720 124160
rect 112772 124148 112778 124160
rect 116118 124148 116124 124160
rect 112772 124120 116124 124148
rect 112772 124108 112778 124120
rect 116118 124108 116124 124120
rect 116176 124108 116182 124160
rect 112622 122748 112628 122800
rect 112680 122788 112686 122800
rect 116118 122788 116124 122800
rect 112680 122760 116124 122788
rect 112680 122748 112686 122760
rect 116118 122748 116124 122760
rect 116176 122748 116182 122800
rect 112530 121388 112536 121440
rect 112588 121428 112594 121440
rect 116118 121428 116124 121440
rect 112588 121400 116124 121428
rect 112588 121388 112594 121400
rect 116118 121388 116124 121400
rect 116176 121388 116182 121440
rect 111610 118600 111616 118652
rect 111668 118640 111674 118652
rect 116118 118640 116124 118652
rect 111668 118612 116124 118640
rect 111668 118600 111674 118612
rect 116118 118600 116124 118612
rect 116176 118600 116182 118652
rect 112438 117240 112444 117292
rect 112496 117280 112502 117292
rect 116118 117280 116124 117292
rect 112496 117252 116124 117280
rect 112496 117240 112502 117252
rect 116118 117240 116124 117252
rect 116176 117240 116182 117292
rect 111518 114452 111524 114504
rect 111576 114492 111582 114504
rect 116118 114492 116124 114504
rect 111576 114464 116124 114492
rect 111576 114452 111582 114464
rect 116118 114452 116124 114464
rect 116176 114452 116182 114504
rect 111426 113092 111432 113144
rect 111484 113132 111490 113144
rect 116118 113132 116124 113144
rect 111484 113104 116124 113132
rect 111484 113092 111490 113104
rect 116118 113092 116124 113104
rect 116176 113092 116182 113144
rect 111334 111732 111340 111784
rect 111392 111772 111398 111784
rect 116118 111772 116124 111784
rect 111392 111744 116124 111772
rect 111392 111732 111398 111744
rect 116118 111732 116124 111744
rect 116176 111732 116182 111784
rect 111242 108944 111248 108996
rect 111300 108984 111306 108996
rect 116118 108984 116124 108996
rect 111300 108956 116124 108984
rect 111300 108944 111306 108956
rect 116118 108944 116124 108956
rect 116176 108944 116182 108996
rect 111150 92420 111156 92472
rect 111208 92460 111214 92472
rect 115934 92460 115940 92472
rect 111208 92432 115940 92460
rect 111208 92420 111214 92432
rect 115934 92420 115940 92432
rect 115992 92420 115998 92472
rect 111058 89632 111064 89684
rect 111116 89672 111122 89684
rect 116118 89672 116124 89684
rect 111116 89644 116124 89672
rect 111116 89632 111122 89644
rect 116118 89632 116124 89644
rect 116176 89632 116182 89684
rect 113818 88272 113824 88324
rect 113876 88312 113882 88324
rect 115934 88312 115940 88324
rect 113876 88284 115940 88312
rect 113876 88272 113882 88284
rect 115934 88272 115940 88284
rect 115992 88272 115998 88324
rect 114462 86980 114468 87032
rect 114520 87020 114526 87032
rect 116670 87020 116676 87032
rect 114520 86992 116676 87020
rect 114520 86980 114526 86992
rect 116670 86980 116676 86992
rect 116728 86980 116734 87032
rect 113910 86912 113916 86964
rect 113968 86952 113974 86964
rect 116026 86952 116032 86964
rect 113968 86924 116032 86952
rect 113968 86912 113974 86924
rect 116026 86912 116032 86924
rect 116084 86912 116090 86964
rect 114002 83920 114008 83972
rect 114060 83960 114066 83972
rect 116578 83960 116584 83972
rect 114060 83932 116584 83960
rect 114060 83920 114066 83932
rect 116578 83920 116584 83932
rect 116636 83920 116642 83972
rect 114094 82764 114100 82816
rect 114152 82804 114158 82816
rect 116118 82804 116124 82816
rect 114152 82776 116124 82804
rect 114152 82764 114158 82776
rect 116118 82764 116124 82776
rect 116176 82764 116182 82816
rect 114186 79976 114192 80028
rect 114244 80016 114250 80028
rect 115934 80016 115940 80028
rect 114244 79988 115940 80016
rect 114244 79976 114250 79988
rect 115934 79976 115940 79988
rect 115992 79976 115998 80028
rect 114186 71748 114192 71800
rect 114244 71788 114250 71800
rect 116026 71788 116032 71800
rect 114244 71760 116032 71788
rect 114244 71748 114250 71760
rect 116026 71748 116032 71760
rect 116084 71748 116090 71800
rect 114094 69028 114100 69080
rect 114152 69068 114158 69080
rect 116210 69068 116216 69080
rect 114152 69040 116216 69068
rect 114152 69028 114158 69040
rect 116210 69028 116216 69040
rect 116268 69028 116274 69080
rect 114002 67600 114008 67652
rect 114060 67640 114066 67652
rect 115934 67640 115940 67652
rect 114060 67612 115940 67640
rect 114060 67600 114066 67612
rect 115934 67600 115940 67612
rect 115992 67600 115998 67652
rect 113910 66240 113916 66292
rect 113968 66280 113974 66292
rect 116578 66280 116584 66292
rect 113968 66252 116584 66280
rect 113968 66240 113974 66252
rect 116578 66240 116584 66252
rect 116636 66240 116642 66292
rect 114462 64676 114468 64728
rect 114520 64716 114526 64728
rect 116578 64716 116584 64728
rect 114520 64688 116584 64716
rect 114520 64676 114526 64688
rect 116578 64676 116584 64688
rect 116636 64676 116642 64728
rect 113818 63520 113824 63572
rect 113876 63560 113882 63572
rect 116026 63560 116032 63572
rect 113876 63532 116032 63560
rect 113876 63520 113882 63532
rect 116026 63520 116032 63532
rect 116084 63520 116090 63572
rect 109678 41420 109684 41472
rect 109736 41460 109742 41472
rect 116118 41460 116124 41472
rect 109736 41432 116124 41460
rect 109736 41420 109742 41432
rect 116118 41420 116124 41432
rect 116176 41420 116182 41472
rect 114094 38632 114100 38684
rect 114152 38672 114158 38684
rect 116394 38672 116400 38684
rect 114152 38644 116400 38672
rect 114152 38632 114158 38644
rect 116394 38632 116400 38644
rect 116452 38632 116458 38684
rect 116210 38496 116216 38548
rect 116268 38536 116274 38548
rect 116394 38536 116400 38548
rect 116268 38508 116400 38536
rect 116268 38496 116274 38508
rect 116394 38496 116400 38508
rect 116452 38496 116458 38548
rect 114186 37272 114192 37324
rect 114244 37312 114250 37324
rect 115934 37312 115940 37324
rect 114244 37284 115940 37312
rect 114244 37272 114250 37284
rect 115934 37272 115940 37284
rect 115992 37272 115998 37324
rect 111058 34484 111064 34536
rect 111116 34524 111122 34536
rect 116118 34524 116124 34536
rect 111116 34496 116124 34524
rect 111116 34484 111122 34496
rect 116118 34484 116124 34496
rect 116176 34484 116182 34536
rect 112438 33124 112444 33176
rect 112496 33164 112502 33176
rect 116118 33164 116124 33176
rect 112496 33136 116124 33164
rect 112496 33124 112502 33136
rect 116118 33124 116124 33136
rect 116176 33124 116182 33176
rect 112530 31764 112536 31816
rect 112588 31804 112594 31816
rect 116118 31804 116124 31816
rect 112588 31776 116124 31804
rect 112588 31764 112594 31776
rect 116118 31764 116124 31776
rect 116176 31764 116182 31816
rect 112622 28976 112628 29028
rect 112680 29016 112686 29028
rect 116118 29016 116124 29028
rect 112680 28988 116124 29016
rect 112680 28976 112686 28988
rect 116118 28976 116124 28988
rect 116176 28976 116182 29028
rect 112714 27616 112720 27668
rect 112772 27656 112778 27668
rect 116118 27656 116124 27668
rect 112772 27628 116124 27656
rect 112772 27616 112778 27628
rect 116118 27616 116124 27628
rect 116176 27616 116182 27668
rect 112806 24828 112812 24880
rect 112864 24868 112870 24880
rect 116118 24868 116124 24880
rect 112864 24840 116124 24868
rect 112864 24828 112870 24840
rect 116118 24828 116124 24840
rect 116176 24828 116182 24880
rect 111150 23468 111156 23520
rect 111208 23508 111214 23520
rect 116118 23508 116124 23520
rect 111208 23480 116124 23508
rect 111208 23468 111214 23480
rect 116118 23468 116124 23480
rect 116176 23468 116182 23520
rect 111242 22108 111248 22160
rect 111300 22148 111306 22160
rect 116118 22148 116124 22160
rect 111300 22120 116124 22148
rect 111300 22108 111306 22120
rect 116118 22108 116124 22120
rect 116176 22108 116182 22160
rect 109770 4156 109776 4208
rect 109828 4196 109834 4208
rect 115934 4196 115940 4208
rect 109828 4168 115940 4196
rect 109828 4156 109834 4168
rect 115934 4156 115940 4168
rect 115992 4156 115998 4208
rect 111058 3924 111064 3936
rect 57946 3896 70716 3924
rect 55186 3828 56594 3856
rect 55186 3788 55214 3828
rect 49620 3760 55214 3788
rect 56566 3788 56594 3828
rect 57946 3788 57974 3896
rect 56566 3760 57974 3788
rect 58636 3828 69612 3856
rect 26206 3012 27614 3040
rect 2498 2864 2504 2916
rect 2556 2904 2562 2916
rect 26206 2904 26234 3012
rect 2556 2876 26234 2904
rect 2556 2864 2562 2876
rect 27586 2836 27614 3012
rect 27586 2808 35894 2836
rect 35866 2632 35894 2808
rect 49620 2644 49648 3760
rect 50080 3692 56594 3720
rect 50080 3448 50108 3692
rect 56566 3652 56594 3692
rect 58636 3652 58664 3828
rect 56566 3624 58664 3652
rect 54036 3556 66254 3584
rect 54036 3516 54064 3556
rect 66226 3516 66254 3556
rect 53944 3488 54064 3516
rect 58820 3488 63494 3516
rect 66226 3488 69060 3516
rect 53944 3448 53972 3488
rect 49804 3420 50108 3448
rect 53806 3420 53972 3448
rect 49804 2644 49832 3420
rect 53806 3244 53834 3420
rect 58820 3244 58848 3488
rect 63466 3448 63494 3488
rect 63466 3420 68968 3448
rect 59188 3352 68876 3380
rect 59188 3312 59216 3352
rect 49896 3216 53834 3244
rect 54036 3216 58848 3244
rect 59096 3284 59216 3312
rect 49896 2644 49924 3216
rect 54036 3176 54064 3216
rect 59096 3176 59124 3284
rect 49988 3148 54064 3176
rect 58636 3148 59124 3176
rect 59280 3216 68784 3244
rect 49988 2644 50016 3148
rect 40678 2632 40684 2644
rect 35866 2604 40684 2632
rect 40678 2592 40684 2604
rect 40736 2592 40742 2644
rect 43622 2592 43628 2644
rect 43680 2632 43686 2644
rect 45646 2632 45652 2644
rect 43680 2604 45652 2632
rect 43680 2592 43686 2604
rect 45646 2592 45652 2604
rect 45704 2592 45710 2644
rect 49602 2592 49608 2644
rect 49660 2592 49666 2644
rect 49786 2592 49792 2644
rect 49844 2592 49850 2644
rect 49878 2592 49884 2644
rect 49936 2592 49942 2644
rect 49970 2592 49976 2644
rect 50028 2592 50034 2644
rect 53926 2592 53932 2644
rect 53984 2632 53990 2644
rect 58636 2632 58664 3148
rect 59280 3108 59308 3216
rect 59004 3080 59308 3108
rect 59004 2644 59032 3080
rect 59096 2876 66116 2904
rect 53984 2604 58664 2632
rect 53984 2592 53990 2604
rect 58986 2592 58992 2644
rect 59044 2592 59050 2644
rect 32766 2524 32772 2576
rect 32824 2564 32830 2576
rect 59096 2564 59124 2876
rect 63466 2808 65840 2836
rect 63466 2700 63494 2808
rect 59740 2672 63494 2700
rect 59740 2644 59768 2672
rect 59722 2592 59728 2644
rect 59780 2592 59786 2644
rect 59814 2592 59820 2644
rect 59872 2632 59878 2644
rect 59872 2604 65656 2632
rect 59872 2592 59878 2604
rect 32824 2536 59124 2564
rect 32824 2524 32830 2536
rect 40678 2456 40684 2508
rect 40736 2496 40742 2508
rect 64874 2496 64880 2508
rect 40736 2468 53834 2496
rect 40736 2456 40742 2468
rect 39666 2388 39672 2440
rect 39724 2428 39730 2440
rect 53650 2428 53656 2440
rect 39724 2400 53656 2428
rect 39724 2388 39730 2400
rect 53650 2388 53656 2400
rect 53708 2388 53714 2440
rect 53806 2428 53834 2468
rect 59740 2468 64880 2496
rect 53806 2400 55904 2428
rect 36354 2320 36360 2372
rect 36412 2360 36418 2372
rect 43622 2360 43628 2372
rect 36412 2332 43628 2360
rect 36412 2320 36418 2332
rect 43622 2320 43628 2332
rect 43680 2320 43686 2372
rect 46290 2320 46296 2372
rect 46348 2360 46354 2372
rect 49786 2360 49792 2372
rect 46348 2332 49792 2360
rect 46348 2320 46354 2332
rect 49786 2320 49792 2332
rect 49844 2320 49850 2372
rect 55876 2360 55904 2400
rect 56226 2388 56232 2440
rect 56284 2428 56290 2440
rect 59740 2428 59768 2468
rect 64874 2456 64880 2468
rect 64932 2456 64938 2508
rect 56284 2400 59768 2428
rect 65628 2428 65656 2604
rect 65812 2496 65840 2808
rect 66088 2700 66116 2876
rect 66088 2672 66254 2700
rect 66226 2632 66254 2672
rect 67542 2632 67548 2644
rect 66226 2604 67548 2632
rect 67542 2592 67548 2604
rect 67600 2592 67606 2644
rect 68756 2564 68784 3216
rect 68848 2644 68876 3352
rect 68940 2644 68968 3420
rect 69032 2644 69060 3488
rect 69584 3312 69612 3828
rect 69584 3284 69888 3312
rect 69860 2644 69888 3284
rect 70688 2644 70716 3896
rect 77266 3896 111064 3924
rect 77266 3856 77294 3896
rect 111058 3884 111064 3896
rect 111116 3884 111122 3936
rect 112438 3856 112444 3868
rect 72436 3828 77294 3856
rect 80026 3828 112444 3856
rect 72436 2644 72464 3828
rect 80026 3788 80054 3828
rect 112438 3816 112444 3828
rect 112496 3816 112502 3868
rect 112530 3788 112536 3800
rect 72528 3760 80054 3788
rect 80256 3760 112536 3788
rect 72528 2644 72556 3760
rect 80256 3584 80284 3760
rect 112530 3748 112536 3760
rect 112588 3748 112594 3800
rect 112622 3720 112628 3732
rect 74506 3556 80284 3584
rect 80900 3692 112628 3720
rect 68830 2592 68836 2644
rect 68888 2592 68894 2644
rect 68922 2592 68928 2644
rect 68980 2592 68986 2644
rect 69014 2592 69020 2644
rect 69072 2592 69078 2644
rect 69842 2592 69848 2644
rect 69900 2592 69906 2644
rect 70670 2592 70676 2644
rect 70728 2592 70734 2644
rect 72418 2592 72424 2644
rect 72476 2592 72482 2644
rect 72510 2592 72516 2644
rect 72568 2592 72574 2644
rect 74506 2564 74534 3556
rect 80900 3244 80928 3692
rect 112622 3680 112628 3692
rect 112680 3680 112686 3732
rect 112714 3652 112720 3664
rect 75012 3216 80928 3244
rect 83844 3624 112720 3652
rect 75012 2644 75040 3216
rect 83844 3176 83872 3624
rect 112714 3612 112720 3624
rect 112772 3612 112778 3664
rect 112806 3584 112812 3596
rect 76300 3148 83872 3176
rect 84166 3556 112812 3584
rect 76300 2644 76328 3148
rect 84166 3108 84194 3556
rect 112806 3544 112812 3556
rect 112864 3544 112870 3596
rect 111150 3516 111156 3528
rect 80026 3080 84194 3108
rect 84396 3488 111156 3516
rect 74994 2592 75000 2644
rect 75052 2592 75058 2644
rect 76282 2592 76288 2644
rect 76340 2592 76346 2644
rect 76466 2592 76472 2644
rect 76524 2632 76530 2644
rect 80026 2632 80054 3080
rect 84396 3040 84424 3488
rect 111150 3476 111156 3488
rect 111208 3476 111214 3528
rect 111242 3448 111248 3460
rect 84120 3012 84424 3040
rect 84488 3420 111248 3448
rect 84120 2972 84148 3012
rect 84028 2944 84148 2972
rect 84028 2644 84056 2944
rect 84488 2644 84516 3420
rect 111242 3408 111248 3420
rect 111300 3408 111306 3460
rect 114186 3380 114192 3392
rect 84580 3352 114192 3380
rect 84580 2644 84608 3352
rect 114186 3340 114192 3352
rect 114244 3340 114250 3392
rect 114094 3312 114100 3324
rect 88306 3284 114100 3312
rect 88306 3176 88334 3284
rect 114094 3272 114100 3284
rect 114152 3272 114158 3324
rect 85132 3148 88334 3176
rect 85132 3040 85160 3148
rect 85040 3012 85160 3040
rect 88306 3080 104894 3108
rect 85040 2700 85068 3012
rect 88306 2972 88334 3080
rect 84764 2672 85068 2700
rect 85316 2944 88334 2972
rect 104866 2972 104894 3080
rect 109586 3000 109592 3052
rect 109644 3040 109650 3052
rect 117958 3040 117964 3052
rect 109644 3012 117964 3040
rect 109644 3000 109650 3012
rect 117958 3000 117964 3012
rect 118016 3000 118022 3052
rect 117682 2972 117688 2984
rect 104866 2944 117688 2972
rect 84764 2644 84792 2672
rect 85316 2644 85344 2944
rect 117682 2932 117688 2944
rect 117740 2932 117746 2984
rect 115842 2904 115848 2916
rect 85776 2876 101444 2904
rect 76524 2604 80054 2632
rect 76524 2592 76530 2604
rect 84010 2592 84016 2644
rect 84068 2592 84074 2644
rect 84470 2592 84476 2644
rect 84528 2592 84534 2644
rect 84562 2592 84568 2644
rect 84620 2592 84626 2644
rect 84746 2592 84752 2644
rect 84804 2592 84810 2644
rect 85298 2592 85304 2644
rect 85356 2592 85362 2644
rect 68756 2536 74534 2564
rect 76558 2524 76564 2576
rect 76616 2564 76622 2576
rect 85776 2564 85804 2876
rect 88306 2808 96614 2836
rect 85850 2592 85856 2644
rect 85908 2632 85914 2644
rect 88306 2632 88334 2808
rect 85908 2604 88334 2632
rect 85908 2592 85914 2604
rect 76616 2536 85804 2564
rect 96586 2564 96614 2808
rect 101416 2700 101444 2876
rect 104866 2876 115848 2904
rect 104360 2808 104572 2836
rect 104360 2700 104388 2808
rect 101416 2672 104388 2700
rect 104544 2700 104572 2808
rect 104866 2700 104894 2876
rect 115842 2864 115848 2876
rect 115900 2864 115906 2916
rect 104544 2672 104894 2700
rect 106246 2808 293954 2836
rect 98270 2592 98276 2644
rect 98328 2632 98334 2644
rect 106090 2632 106096 2644
rect 98328 2604 106096 2632
rect 98328 2592 98334 2604
rect 106090 2592 106096 2604
rect 106148 2592 106154 2644
rect 106246 2564 106274 2808
rect 96586 2536 106274 2564
rect 76616 2524 76622 2536
rect 72510 2496 72516 2508
rect 65812 2468 72516 2496
rect 72510 2456 72516 2468
rect 72568 2456 72574 2508
rect 109586 2456 109592 2508
rect 109644 2496 109650 2508
rect 116578 2496 116584 2508
rect 109644 2468 116584 2496
rect 109644 2456 109650 2468
rect 116578 2456 116584 2468
rect 116636 2456 116642 2508
rect 293926 2496 293954 2808
rect 425808 2808 443684 2836
rect 425808 2508 425836 2808
rect 443656 2508 443684 2808
rect 294782 2496 294788 2508
rect 293926 2468 294788 2496
rect 294782 2456 294788 2468
rect 294840 2456 294846 2508
rect 425790 2456 425796 2508
rect 425848 2456 425854 2508
rect 443638 2456 443644 2508
rect 443696 2456 443702 2508
rect 65628 2400 66254 2428
rect 56284 2388 56290 2400
rect 59814 2360 59820 2372
rect 55876 2332 59820 2360
rect 59814 2320 59820 2332
rect 59872 2320 59878 2372
rect 66226 2360 66254 2400
rect 68830 2388 68836 2440
rect 68888 2428 68894 2440
rect 84010 2428 84016 2440
rect 68888 2400 84016 2428
rect 68888 2388 68894 2400
rect 84010 2388 84016 2400
rect 84068 2388 84074 2440
rect 106182 2388 106188 2440
rect 106240 2428 106246 2440
rect 116670 2428 116676 2440
rect 106240 2400 116676 2428
rect 106240 2388 106246 2400
rect 116670 2388 116676 2400
rect 116728 2388 116734 2440
rect 76558 2360 76564 2372
rect 66226 2332 76564 2360
rect 76558 2320 76564 2332
rect 76616 2320 76622 2372
rect 102962 2320 102968 2372
rect 103020 2360 103026 2372
rect 116762 2360 116768 2372
rect 103020 2332 116768 2360
rect 103020 2320 103026 2332
rect 116762 2320 116768 2332
rect 116820 2320 116826 2372
rect 42978 2252 42984 2304
rect 43036 2292 43042 2304
rect 49878 2292 49884 2304
rect 43036 2264 49884 2292
rect 43036 2252 43042 2264
rect 49878 2252 49884 2264
rect 49936 2252 49942 2304
rect 52914 2252 52920 2304
rect 52972 2292 52978 2304
rect 58986 2292 58992 2304
rect 52972 2264 58992 2292
rect 52972 2252 52978 2264
rect 58986 2252 58992 2264
rect 59044 2252 59050 2304
rect 68922 2252 68928 2304
rect 68980 2292 68986 2304
rect 84470 2292 84476 2304
rect 68980 2264 84476 2292
rect 68980 2252 68986 2264
rect 84470 2252 84476 2264
rect 84528 2252 84534 2304
rect 99650 2252 99656 2304
rect 99708 2292 99714 2304
rect 116854 2292 116860 2304
rect 99708 2264 116860 2292
rect 99708 2252 99714 2264
rect 116854 2252 116860 2264
rect 116912 2252 116918 2304
rect 69658 2184 69664 2236
rect 69716 2224 69722 2236
rect 84746 2224 84752 2236
rect 69716 2196 84752 2224
rect 69716 2184 69722 2196
rect 84746 2184 84752 2196
rect 84804 2184 84810 2236
rect 96338 2184 96344 2236
rect 96396 2224 96402 2236
rect 116946 2224 116952 2236
rect 96396 2196 116952 2224
rect 96396 2184 96402 2196
rect 116946 2184 116952 2196
rect 117004 2184 117010 2236
rect 63034 2116 63040 2168
rect 63092 2156 63098 2168
rect 63092 2128 66254 2156
rect 63092 2116 63098 2128
rect 66226 2020 66254 2128
rect 69842 2116 69848 2168
rect 69900 2156 69906 2168
rect 76282 2156 76288 2168
rect 69900 2128 76288 2156
rect 69900 2116 69906 2128
rect 76282 2116 76288 2128
rect 76340 2116 76346 2168
rect 93026 2116 93032 2168
rect 93084 2156 93090 2168
rect 117038 2156 117044 2168
rect 93084 2128 117044 2156
rect 93084 2116 93090 2128
rect 117038 2116 117044 2128
rect 117096 2116 117102 2168
rect 70670 2048 70676 2100
rect 70728 2088 70734 2100
rect 74994 2088 75000 2100
rect 70728 2060 75000 2088
rect 70728 2048 70734 2060
rect 74994 2048 75000 2060
rect 75052 2048 75058 2100
rect 89622 2048 89628 2100
rect 89680 2088 89686 2100
rect 117130 2088 117136 2100
rect 89680 2060 117136 2088
rect 89680 2048 89686 2060
rect 117130 2048 117136 2060
rect 117188 2048 117194 2100
rect 72418 2020 72424 2032
rect 66226 1992 72424 2020
rect 72418 1980 72424 1992
rect 72476 1980 72482 2032
rect 86402 1980 86408 2032
rect 86460 2020 86466 2032
rect 117222 2020 117228 2032
rect 86460 1992 117228 2020
rect 86460 1980 86466 1992
rect 117222 1980 117228 1992
rect 117280 1980 117286 2032
rect 82630 1912 82636 1964
rect 82688 1952 82694 1964
rect 116486 1952 116492 1964
rect 82688 1924 116492 1952
rect 82688 1912 82694 1924
rect 116486 1912 116492 1924
rect 116544 1912 116550 1964
rect 79318 1844 79324 1896
rect 79376 1884 79382 1896
rect 116394 1884 116400 1896
rect 79376 1856 116400 1884
rect 79376 1844 79382 1856
rect 116394 1844 116400 1856
rect 116452 1844 116458 1896
rect 72694 1776 72700 1828
rect 72752 1816 72758 1828
rect 109678 1816 109684 1828
rect 72752 1788 109684 1816
rect 72752 1776 72758 1788
rect 109678 1776 109684 1788
rect 109736 1776 109742 1828
rect 76006 1708 76012 1760
rect 76064 1748 76070 1760
rect 116302 1748 116308 1760
rect 76064 1720 116308 1748
rect 76064 1708 76070 1720
rect 116302 1708 116308 1720
rect 116360 1708 116366 1760
rect 32674 1640 32680 1692
rect 32732 1680 32738 1692
rect 116210 1680 116216 1692
rect 32732 1652 116216 1680
rect 32732 1640 32738 1652
rect 116210 1640 116216 1652
rect 116268 1640 116274 1692
rect 29270 1572 29276 1624
rect 29328 1612 29334 1624
rect 116026 1612 116032 1624
rect 29328 1584 116032 1612
rect 29328 1572 29334 1584
rect 116026 1572 116032 1584
rect 116084 1572 116090 1624
rect 25958 1504 25964 1556
rect 26016 1544 26022 1556
rect 116118 1544 116124 1556
rect 26016 1516 116124 1544
rect 26016 1504 26022 1516
rect 116118 1504 116124 1516
rect 116176 1504 116182 1556
rect 22646 1436 22652 1488
rect 22704 1476 22710 1488
rect 115934 1476 115940 1488
rect 22704 1448 115940 1476
rect 22704 1436 22710 1448
rect 115934 1436 115940 1448
rect 115992 1436 115998 1488
rect 117682 1436 117688 1488
rect 117740 1476 117746 1488
rect 143626 1476 143632 1488
rect 117740 1448 143632 1476
rect 117740 1436 117746 1448
rect 143626 1436 143632 1448
rect 143684 1436 143690 1488
rect 5994 1368 6000 1420
rect 6052 1408 6058 1420
rect 109770 1408 109776 1420
rect 6052 1380 109776 1408
rect 6052 1368 6058 1380
rect 109770 1368 109776 1380
rect 109828 1368 109834 1420
rect 117958 1368 117964 1420
rect 118016 1408 118022 1420
rect 193582 1408 193588 1420
rect 118016 1380 193588 1408
rect 118016 1368 118022 1380
rect 193582 1368 193588 1380
rect 193640 1368 193646 1420
rect 294782 1368 294788 1420
rect 294840 1408 294846 1420
rect 343634 1408 343640 1420
rect 294840 1380 343640 1408
rect 294840 1368 294846 1380
rect 343634 1368 343640 1380
rect 343692 1368 343698 1420
rect 491294 1368 491300 1420
rect 491352 1408 491358 1420
rect 493594 1408 493600 1420
rect 491352 1380 493600 1408
rect 491352 1368 491358 1380
rect 493594 1368 493600 1380
rect 493652 1368 493658 1420
<< via1 >>
rect 146668 161372 146720 161424
rect 153752 161372 153804 161424
rect 136640 160080 136692 160132
rect 144276 160080 144328 160132
rect 83648 160012 83700 160064
rect 167000 160012 167052 160064
rect 170220 160012 170272 160064
rect 198924 160012 198976 160064
rect 203064 160012 203116 160064
rect 211068 160012 211120 160064
rect 211436 160012 211488 160064
rect 280344 160012 280396 160064
rect 281264 160012 281316 160064
rect 332692 160012 332744 160064
rect 335084 160012 335136 160064
rect 374000 160012 374052 160064
rect 378876 160012 378928 160064
rect 398564 160012 398616 160064
rect 25596 159944 25648 159996
rect 109868 159944 109920 159996
rect 117228 159944 117280 159996
rect 191748 159944 191800 159996
rect 198004 159944 198056 159996
rect 269120 159944 269172 159996
rect 271236 159944 271288 159996
rect 272800 159944 272852 159996
rect 275376 159944 275428 159996
rect 329104 159944 329156 159996
rect 329196 159944 329248 159996
rect 369860 159944 369912 159996
rect 372160 159944 372212 159996
rect 396172 159944 396224 159996
rect 399024 159944 399076 159996
rect 408500 159944 408552 159996
rect 476120 159944 476172 159996
rect 70124 159876 70176 159928
rect 148692 159876 148744 159928
rect 152464 159876 152516 159928
rect 160100 159876 160152 159928
rect 160192 159876 160244 159928
rect 188252 159876 188304 159928
rect 191288 159876 191340 159928
rect 264888 159876 264940 159928
rect 268660 159876 268712 159928
rect 324044 159876 324096 159928
rect 328368 159876 328420 159928
rect 369492 159876 369544 159928
rect 379704 159876 379756 159928
rect 405832 159876 405884 159928
rect 470508 159876 470560 159928
rect 471428 159876 471480 159928
rect 477684 159876 477736 159928
rect 480628 159876 480680 159928
rect 485964 159876 486016 159928
rect 56692 159808 56744 159860
rect 136548 159808 136600 159860
rect 142620 159808 142672 159860
rect 146300 159808 146352 159860
rect 153752 159808 153804 159860
rect 175004 159808 175056 159860
rect 63408 159740 63460 159792
rect 18880 159672 18932 159724
rect 107292 159672 107344 159724
rect 109684 159672 109736 159724
rect 137652 159672 137704 159724
rect 146852 159740 146904 159792
rect 148600 159740 148652 159792
rect 144276 159672 144328 159724
rect 148784 159672 148836 159724
rect 148968 159672 149020 159724
rect 150808 159740 150860 159792
rect 152556 159740 152608 159792
rect 153476 159740 153528 159792
rect 180708 159808 180760 159860
rect 184572 159808 184624 159860
rect 259552 159808 259604 159860
rect 261944 159808 261996 159860
rect 318800 159808 318852 159860
rect 320824 159808 320876 159860
rect 362960 159808 363012 159860
rect 376300 159808 376352 159860
rect 406200 159808 406252 159860
rect 409972 159808 410024 159860
rect 417424 159808 417476 159860
rect 467196 159808 467248 159860
rect 473360 159808 473412 159860
rect 177856 159740 177908 159792
rect 253940 159740 253992 159792
rect 255228 159740 255280 159792
rect 313372 159740 313424 159792
rect 314108 159740 314160 159792
rect 357992 159740 358044 159792
rect 365444 159740 365496 159792
rect 395528 159740 395580 159792
rect 396540 159740 396592 159792
rect 413192 159740 413244 159792
rect 424324 159740 424376 159792
rect 442816 159740 442868 159792
rect 472256 159740 472308 159792
rect 479432 159740 479484 159792
rect 479800 159740 479852 159792
rect 485228 159740 485280 159792
rect 164148 159672 164200 159724
rect 167736 159672 167788 159724
rect 246948 159672 247000 159724
rect 248512 159672 248564 159724
rect 301412 159672 301464 159724
rect 49976 159604 50028 159656
rect 142252 159604 142304 159656
rect 143356 159604 143408 159656
rect 148600 159604 148652 159656
rect 160100 159604 160152 159656
rect 161020 159604 161072 159656
rect 240324 159604 240376 159656
rect 241796 159604 241848 159656
rect 303528 159672 303580 159724
rect 309048 159672 309100 159724
rect 354864 159672 354916 159724
rect 357808 159672 357860 159724
rect 369216 159672 369268 159724
rect 369584 159672 369636 159724
rect 401048 159672 401100 159724
rect 403256 159672 403308 159724
rect 416596 159672 416648 159724
rect 420920 159672 420972 159724
rect 440424 159672 440476 159724
rect 302332 159604 302384 159656
rect 349252 159604 349304 159656
rect 351920 159604 351972 159656
rect 385316 159604 385368 159656
rect 389824 159604 389876 159656
rect 413836 159604 413888 159656
rect 417516 159604 417568 159656
rect 437664 159604 437716 159656
rect 448704 159604 448756 159656
rect 455880 159604 455932 159656
rect 32312 159536 32364 159588
rect 126244 159536 126296 159588
rect 127624 159536 127676 159588
rect 139860 159536 139912 159588
rect 139952 159536 140004 159588
rect 157248 159536 157300 159588
rect 157616 159536 157668 159588
rect 239312 159536 239364 159588
rect 250996 159536 251048 159588
rect 310612 159536 310664 159588
rect 315764 159536 315816 159588
rect 358912 159536 358964 159588
rect 362868 159536 362920 159588
rect 395988 159536 396040 159588
rect 407488 159536 407540 159588
rect 429936 159536 429988 159588
rect 450360 159536 450412 159588
rect 457168 159536 457220 159588
rect 458732 159536 458784 159588
rect 465080 159536 465132 159588
rect 468024 159536 468076 159588
rect 476028 159536 476080 159588
rect 478972 159536 479024 159588
rect 484584 159536 484636 159588
rect 43260 159468 43312 159520
rect 36544 159400 36596 159452
rect 135168 159400 135220 159452
rect 136548 159468 136600 159520
rect 137376 159400 137428 159452
rect 137468 159400 137520 159452
rect 144184 159468 144236 159520
rect 225236 159468 225288 159520
rect 231676 159468 231728 159520
rect 295524 159468 295576 159520
rect 295616 159468 295668 159520
rect 342444 159468 342496 159520
rect 347688 159468 347740 159520
rect 354220 159468 354272 159520
rect 356152 159468 356204 159520
rect 390560 159468 390612 159520
rect 392308 159468 392360 159520
rect 404268 159468 404320 159520
rect 410800 159468 410852 159520
rect 432512 159468 432564 159520
rect 449532 159468 449584 159520
rect 455512 159468 455564 159520
rect 457076 159468 457128 159520
rect 464344 159468 464396 159520
rect 6276 159332 6328 159384
rect 122840 159332 122892 159384
rect 123116 159332 123168 159384
rect 142620 159332 142672 159384
rect 144828 159400 144880 159452
rect 144920 159400 144972 159452
rect 146208 159400 146260 159452
rect 146300 159400 146352 159452
rect 147128 159400 147180 159452
rect 147588 159400 147640 159452
rect 149060 159400 149112 159452
rect 149152 159400 149204 159452
rect 150808 159400 150860 159452
rect 150900 159400 150952 159452
rect 234068 159400 234120 159452
rect 234988 159400 235040 159452
rect 298008 159400 298060 159452
rect 301504 159400 301556 159452
rect 349068 159400 349120 159452
rect 349344 159400 349396 159452
rect 353208 159400 353260 159452
rect 358636 159400 358688 159452
rect 392768 159400 392820 159452
rect 404084 159400 404136 159452
rect 427360 159400 427412 159452
rect 427636 159400 427688 159452
rect 445392 159400 445444 159452
rect 451188 159400 451240 159452
rect 456800 159400 456852 159452
rect 459652 159400 459704 159452
rect 466460 159400 466512 159452
rect 468852 159400 468904 159452
rect 474832 159400 474884 159452
rect 477316 159400 477368 159452
rect 483296 159400 483348 159452
rect 518808 159400 518860 159452
rect 522672 159400 522724 159452
rect 223672 159332 223724 159384
rect 224960 159332 225012 159384
rect 290648 159332 290700 159384
rect 294788 159332 294840 159384
rect 342260 159332 342312 159384
rect 342720 159332 342772 159384
rect 343640 159332 343692 159384
rect 346032 159332 346084 159384
rect 382832 159332 382884 159384
rect 383108 159332 383160 159384
rect 411352 159332 411404 159384
rect 414204 159332 414256 159384
rect 435088 159332 435140 159384
rect 447876 159332 447928 159384
rect 456892 159332 456944 159384
rect 469680 159332 469732 159384
rect 477408 159332 477460 159384
rect 478144 159332 478196 159384
rect 483204 159332 483256 159384
rect 518716 159332 518768 159384
rect 523500 159332 523552 159384
rect 76932 159264 76984 159316
rect 152464 159264 152516 159316
rect 152556 159264 152608 159316
rect 156052 159264 156104 159316
rect 163504 159264 163556 159316
rect 193588 159264 193640 159316
rect 193680 159264 193732 159316
rect 197360 159264 197412 159316
rect 201408 159264 201460 159316
rect 207388 159264 207440 159316
rect 208124 159264 208176 159316
rect 212448 159264 212500 159316
rect 214012 159264 214064 159316
rect 281540 159264 281592 159316
rect 282092 159264 282144 159316
rect 334164 159264 334216 159316
rect 334256 159264 334308 159316
rect 374092 159264 374144 159316
rect 378048 159264 378100 159316
rect 388352 159264 388404 159316
rect 395712 159264 395764 159316
rect 404728 159264 404780 159316
rect 460480 159264 460532 159316
rect 466644 159264 466696 159316
rect 93676 159196 93728 159248
rect 175832 159196 175884 159248
rect 86960 159128 87012 159180
rect 169760 159128 169812 159180
rect 173624 159128 173676 159180
rect 175924 159128 175976 159180
rect 100484 159060 100536 159112
rect 183100 159196 183152 159248
rect 187056 159196 187108 159248
rect 216772 159196 216824 159248
rect 218244 159196 218296 159248
rect 284392 159196 284444 159248
rect 287980 159196 288032 159248
rect 338764 159196 338816 159248
rect 339316 159196 339368 159248
rect 377956 159196 378008 159248
rect 385592 159196 385644 159248
rect 398840 159196 398892 159248
rect 453764 159196 453816 159248
rect 459560 159196 459612 159248
rect 462964 159196 463016 159248
rect 469220 159196 469272 159248
rect 176108 159128 176160 159180
rect 193680 159128 193732 159180
rect 193772 159128 193824 159180
rect 180340 159060 180392 159112
rect 203892 159128 203944 159180
rect 206928 159128 206980 159180
rect 220636 159128 220688 159180
rect 220728 159128 220780 159180
rect 283196 159128 283248 159180
rect 284668 159128 284720 159180
rect 285772 159128 285824 159180
rect 107200 158992 107252 159044
rect 185584 158992 185636 159044
rect 193588 158992 193640 159044
rect 196992 158992 197044 159044
rect 73528 158924 73580 158976
rect 107568 158924 107620 158976
rect 119804 158924 119856 158976
rect 127624 158924 127676 158976
rect 96252 158856 96304 158908
rect 121828 158856 121880 158908
rect 124036 158856 124088 158908
rect 192668 158924 192720 158976
rect 130752 158856 130804 158908
rect 195152 158856 195204 158908
rect 207388 159060 207440 159112
rect 212724 159060 212776 159112
rect 212816 159060 212868 159112
rect 222108 159060 222160 159112
rect 224132 159060 224184 159112
rect 288256 159128 288308 159180
rect 288900 159128 288952 159180
rect 338396 159128 338448 159180
rect 338488 159128 338540 159180
rect 340788 159128 340840 159180
rect 341892 159128 341944 159180
rect 378232 159128 378284 159180
rect 457904 159128 457956 159180
rect 463884 159128 463936 159180
rect 307392 159060 307444 159112
rect 349344 159060 349396 159112
rect 351092 159060 351144 159112
rect 382280 159060 382332 159112
rect 409144 159060 409196 159112
rect 410892 159060 410944 159112
rect 452844 159060 452896 159112
rect 459652 159060 459704 159112
rect 461308 159060 461360 159112
rect 467840 159060 467892 159112
rect 200580 158992 200632 159044
rect 197176 158924 197228 158976
rect 212632 158924 212684 158976
rect 227720 158992 227772 159044
rect 230848 158992 230900 159044
rect 295156 158992 295208 159044
rect 298100 158992 298152 159044
rect 300768 158992 300820 159044
rect 308220 158992 308272 159044
rect 347688 158992 347740 159044
rect 347780 158992 347832 159044
rect 378784 158992 378836 159044
rect 384672 158992 384724 159044
rect 388444 158992 388496 159044
rect 388996 158992 389048 159044
rect 403256 158992 403308 159044
rect 455420 158992 455472 159044
rect 463516 158992 463568 159044
rect 465540 158992 465592 159044
rect 472440 158992 472492 159044
rect 473912 158992 473964 159044
rect 480260 158992 480312 159044
rect 217324 158924 217376 158976
rect 220452 158924 220504 158976
rect 237564 158924 237616 158976
rect 299480 158924 299532 158976
rect 301412 158924 301464 158976
rect 308588 158924 308640 158976
rect 314936 158924 314988 158976
rect 357440 158924 357492 158976
rect 361212 158924 361264 158976
rect 201408 158856 201460 158908
rect 207296 158856 207348 158908
rect 231768 158856 231820 158908
rect 238392 158856 238444 158908
rect 242808 158856 242860 158908
rect 244280 158856 244332 158908
rect 305368 158856 305420 158908
rect 305644 158856 305696 158908
rect 307668 158856 307720 158908
rect 310704 158856 310756 158908
rect 311992 158856 312044 158908
rect 312452 158856 312504 158908
rect 313464 158856 313516 158908
rect 322480 158856 322532 158908
rect 365168 158856 365220 158908
rect 102968 158788 103020 158840
rect 125508 158788 125560 158840
rect 126520 158788 126572 158840
rect 154488 158788 154540 158840
rect 156788 158788 156840 158840
rect 194508 158788 194560 158840
rect 194692 158788 194744 158840
rect 203708 158788 203760 158840
rect 206928 158788 206980 158840
rect 213828 158788 213880 158840
rect 214840 158788 214892 158840
rect 221740 158788 221792 158840
rect 261116 158788 261168 158840
rect 317052 158788 317104 158840
rect 106372 158720 106424 158772
rect 127256 158720 127308 158772
rect 127348 158720 127400 158772
rect 129740 158720 129792 158772
rect 133236 158720 133288 158772
rect 158720 158720 158772 158772
rect 81072 158652 81124 158704
rect 163044 158652 163096 158704
rect 67640 158584 67692 158636
rect 163228 158652 163280 158704
rect 167644 158652 167696 158704
rect 163320 158584 163372 158636
rect 167552 158584 167604 158636
rect 171140 158720 171192 158772
rect 172612 158720 172664 158772
rect 175832 158720 175884 158772
rect 176660 158720 176712 158772
rect 180708 158720 180760 158772
rect 167828 158652 167880 158704
rect 180892 158652 180944 158704
rect 183744 158720 183796 158772
rect 204904 158720 204956 158772
rect 210608 158720 210660 158772
rect 215392 158720 215444 158772
rect 221556 158720 221608 158772
rect 223856 158720 223908 158772
rect 240876 158720 240928 158772
rect 243360 158720 243412 158772
rect 254400 158720 254452 158772
rect 255504 158720 255556 158772
rect 258540 158720 258592 158772
rect 261024 158720 261076 158772
rect 264428 158720 264480 158772
rect 266360 158720 266412 158772
rect 267832 158720 267884 158772
rect 320272 158788 320324 158840
rect 327540 158788 327592 158840
rect 330484 158788 330536 158840
rect 319168 158720 319220 158772
rect 321560 158720 321612 158772
rect 321652 158720 321704 158772
rect 181720 158652 181772 158704
rect 181996 158652 182048 158704
rect 256792 158652 256844 158704
rect 363144 158788 363196 158840
rect 369216 158924 369268 158976
rect 384948 158924 385000 158976
rect 420092 158924 420144 158976
rect 423588 158924 423640 158976
rect 446128 158924 446180 158976
rect 453856 158924 453908 158976
rect 454592 158924 454644 158976
rect 461860 158924 461912 158976
rect 464620 158924 464672 158976
rect 471244 158924 471296 158976
rect 475568 158924 475620 158976
rect 482008 158924 482060 158976
rect 367928 158856 367980 158908
rect 386236 158856 386288 158908
rect 391480 158856 391532 158908
rect 394332 158856 394384 158908
rect 412548 158856 412600 158908
rect 413100 158856 413152 158908
rect 456248 158856 456300 158908
rect 462964 158856 463016 158908
rect 466368 158856 466420 158908
rect 472348 158856 472400 158908
rect 474740 158856 474792 158908
rect 481364 158856 481416 158908
rect 481456 158856 481508 158908
rect 486516 158856 486568 158908
rect 508320 158856 508372 158908
rect 510068 158856 510120 158908
rect 385776 158788 385828 158840
rect 388076 158788 388128 158840
rect 390376 158788 390428 158840
rect 405740 158788 405792 158840
rect 409236 158788 409288 158840
rect 413376 158788 413428 158840
rect 419632 158788 419684 158840
rect 463792 158788 463844 158840
rect 471428 158788 471480 158840
rect 476396 158788 476448 158840
rect 481640 158788 481692 158840
rect 505284 158788 505336 158840
rect 507584 158788 507636 158840
rect 330668 158720 330720 158772
rect 367192 158720 367244 158772
rect 374644 158720 374696 158772
rect 384672 158720 384724 158772
rect 384764 158720 384816 158772
rect 389180 158720 389232 158772
rect 416688 158720 416740 158772
rect 419540 158720 419592 158772
rect 452016 158720 452068 158772
rect 458180 158720 458232 158772
rect 462136 158720 462188 158772
rect 467932 158720 467984 158772
rect 473084 158720 473136 158772
rect 478972 158720 479024 158772
rect 482284 158720 482336 158772
rect 487252 158720 487304 158772
rect 505744 158720 505796 158772
rect 506756 158720 506808 158772
rect 507032 158720 507084 158772
rect 508412 158720 508464 158772
rect 509424 158720 509476 158772
rect 511724 158720 511776 158772
rect 514944 158720 514996 158772
rect 518532 158720 518584 158772
rect 170312 158584 170364 158636
rect 171968 158584 172020 158636
rect 250076 158584 250128 158636
rect 74356 158516 74408 158568
rect 71044 158448 71096 158500
rect 173072 158448 173124 158500
rect 175280 158516 175332 158568
rect 252744 158516 252796 158568
rect 175372 158448 175424 158500
rect 178684 158448 178736 158500
rect 255412 158448 255464 158500
rect 64236 158380 64288 158432
rect 163320 158380 163372 158432
rect 60924 158312 60976 158364
rect 165436 158380 165488 158432
rect 168564 158380 168616 158432
rect 247132 158380 247184 158432
rect 165252 158312 165304 158364
rect 245016 158312 245068 158364
rect 54208 158244 54260 158296
rect 160284 158244 160336 158296
rect 161848 158244 161900 158296
rect 242072 158244 242124 158296
rect 50804 158176 50856 158228
rect 157708 158176 157760 158228
rect 158444 158176 158496 158228
rect 238944 158176 238996 158228
rect 256884 158176 256936 158228
rect 315028 158176 315080 158228
rect 47492 158108 47544 158160
rect 155040 158108 155092 158160
rect 155132 158108 155184 158160
rect 237380 158108 237432 158160
rect 246764 158108 246816 158160
rect 306932 158108 306984 158160
rect 37372 158040 37424 158092
rect 146392 158040 146444 158092
rect 148416 158040 148468 158092
rect 231952 158040 232004 158092
rect 233332 158040 233384 158092
rect 297088 158040 297140 158092
rect 300676 158040 300728 158092
rect 348056 158040 348108 158092
rect 388 157972 440 158024
rect 118884 157972 118936 158024
rect 127256 157972 127308 158024
rect 127900 157972 127952 158024
rect 131580 157972 131632 158024
rect 219348 157972 219400 158024
rect 240048 157972 240100 158024
rect 302240 157972 302292 158024
rect 77760 157904 77812 157956
rect 84476 157836 84528 157888
rect 175924 157836 175976 157888
rect 176200 157904 176252 157956
rect 182272 157904 182324 157956
rect 185400 157904 185452 157956
rect 260472 157904 260524 157956
rect 178040 157836 178092 157888
rect 87788 157768 87840 157820
rect 181352 157768 181404 157820
rect 91192 157700 91244 157752
rect 188528 157836 188580 157888
rect 188804 157836 188856 157888
rect 263048 157836 263100 157888
rect 94596 157632 94648 157684
rect 190644 157768 190696 157820
rect 195520 157768 195572 157820
rect 267740 157768 267792 157820
rect 181720 157700 181772 157752
rect 181628 157632 181680 157684
rect 185400 157632 185452 157684
rect 190460 157700 190512 157752
rect 263692 157700 263744 157752
rect 236184 157632 236236 157684
rect 97908 157564 97960 157616
rect 193220 157564 193272 157616
rect 197360 157564 197412 157616
rect 251456 157564 251508 157616
rect 111340 157496 111392 157548
rect 203432 157496 203484 157548
rect 204904 157496 204956 157548
rect 258080 157496 258132 157548
rect 114744 157428 114796 157480
rect 206560 157428 206612 157480
rect 141700 157360 141752 157412
rect 227076 157360 227128 157412
rect 52460 157292 52512 157344
rect 158628 157292 158680 157344
rect 158720 157292 158772 157344
rect 55864 157224 55916 157276
rect 161572 157224 161624 157276
rect 45744 157156 45796 157208
rect 153752 157156 153804 157208
rect 160100 157156 160152 157208
rect 202788 157224 202840 157276
rect 204904 157292 204956 157344
rect 270500 157292 270552 157344
rect 204996 157224 205048 157276
rect 205088 157224 205140 157276
rect 273260 157224 273312 157276
rect 283840 157224 283892 157276
rect 335544 157224 335596 157276
rect 192116 157156 192168 157208
rect 265164 157156 265216 157208
rect 280436 157156 280488 157208
rect 333060 157156 333112 157208
rect 39028 157088 39080 157140
rect 147680 157088 147732 157140
rect 166908 157088 166960 157140
rect 245844 157088 245896 157140
rect 273720 157088 273772 157140
rect 327908 157088 327960 157140
rect 35716 157020 35768 157072
rect 145472 157020 145524 157072
rect 146852 157020 146904 157072
rect 150440 157020 150492 157072
rect 151728 157020 151780 157072
rect 234804 157020 234856 157072
rect 277124 157020 277176 157072
rect 330484 157020 330536 157072
rect 24768 156952 24820 157004
rect 136916 156952 136968 157004
rect 138296 156952 138348 157004
rect 224132 156952 224184 157004
rect 270316 156952 270368 157004
rect 325332 156952 325384 157004
rect 18052 156884 18104 156936
rect 132500 156884 132552 156936
rect 134892 156884 134944 156936
rect 210516 156884 210568 156936
rect 210608 156884 210660 156936
rect 222292 156884 222344 156936
rect 226616 156884 226668 156936
rect 291936 156884 291988 156936
rect 293868 156884 293920 156936
rect 342720 156884 342772 156936
rect 21364 156816 21416 156868
rect 135260 156816 135312 156868
rect 139124 156816 139176 156868
rect 225144 156816 225196 156868
rect 230020 156816 230072 156868
rect 294052 156816 294104 156868
rect 297272 156816 297324 156868
rect 345112 156816 345164 156868
rect 128176 156748 128228 156800
rect 214104 156748 214156 156800
rect 14648 156680 14700 156732
rect 130108 156680 130160 156732
rect 132408 156680 132460 156732
rect 219900 156748 219952 156800
rect 286324 156748 286376 156800
rect 287152 156748 287204 156800
rect 338120 156748 338172 156800
rect 219992 156680 220044 156732
rect 223212 156680 223264 156732
rect 289360 156680 289412 156732
rect 290556 156680 290608 156732
rect 340696 156680 340748 156732
rect 344376 156680 344428 156732
rect 381820 156680 381872 156732
rect 2044 156612 2096 156664
rect 120448 156612 120500 156664
rect 124864 156612 124916 156664
rect 209688 156612 209740 156664
rect 209780 156612 209832 156664
rect 210700 156612 210752 156664
rect 210792 156612 210844 156664
rect 214196 156612 214248 156664
rect 214288 156612 214340 156664
rect 216404 156612 216456 156664
rect 216496 156612 216548 156664
rect 283104 156612 283156 156664
rect 337660 156612 337712 156664
rect 376668 156612 376720 156664
rect 498292 156612 498344 156664
rect 499304 156612 499356 156664
rect 59268 156544 59320 156596
rect 164148 156544 164200 156596
rect 164240 156544 164292 156596
rect 228364 156544 228416 156596
rect 72700 156476 72752 156528
rect 174452 156476 174504 156528
rect 175004 156476 175056 156528
rect 79416 156408 79468 156460
rect 179604 156408 179656 156460
rect 92848 156340 92900 156392
rect 189816 156340 189868 156392
rect 198832 156476 198884 156528
rect 204904 156476 204956 156528
rect 204996 156476 205048 156528
rect 210424 156476 210476 156528
rect 210516 156476 210568 156528
rect 221372 156476 221424 156528
rect 223580 156476 223632 156528
rect 281632 156476 281684 156528
rect 202696 156408 202748 156460
rect 205088 156408 205140 156460
rect 210700 156408 210752 156460
rect 279056 156408 279108 156460
rect 230940 156340 230992 156392
rect 101312 156272 101364 156324
rect 196256 156272 196308 156324
rect 202788 156272 202840 156324
rect 108028 156204 108080 156256
rect 200304 156204 200356 156256
rect 205916 156204 205968 156256
rect 210424 156272 210476 156324
rect 219532 156272 219584 156324
rect 222108 156272 222160 156324
rect 269488 156272 269540 156324
rect 118148 156136 118200 156188
rect 203892 156136 203944 156188
rect 210608 156204 210660 156256
rect 213184 156204 213236 156256
rect 223580 156204 223632 156256
rect 211620 156136 211672 156188
rect 220636 156136 220688 156188
rect 266912 156204 266964 156256
rect 227720 156136 227772 156188
rect 272064 156136 272116 156188
rect 121460 156068 121512 156120
rect 205732 156068 205784 156120
rect 211068 156068 211120 156120
rect 273904 156068 273956 156120
rect 11244 156000 11296 156052
rect 127532 156000 127584 156052
rect 135812 156000 135864 156052
rect 222568 156000 222620 156052
rect 145012 155932 145064 155984
rect 229652 155932 229704 155984
rect 60096 155864 60148 155916
rect 84752 155864 84804 155916
rect 88708 155864 88760 155916
rect 186780 155864 186832 155916
rect 189632 155864 189684 155916
rect 263784 155864 263836 155916
rect 299756 155864 299808 155916
rect 347872 155864 347924 155916
rect 12164 155796 12216 155848
rect 109040 155796 109092 155848
rect 112260 155796 112312 155848
rect 204352 155796 204404 155848
rect 206468 155796 206520 155848
rect 276112 155796 276164 155848
rect 296444 155796 296496 155848
rect 345204 155796 345256 155848
rect 46572 155728 46624 155780
rect 75828 155728 75880 155780
rect 81900 155728 81952 155780
rect 181444 155728 181496 155780
rect 186228 155728 186280 155780
rect 260840 155728 260892 155780
rect 293040 155728 293092 155780
rect 342352 155728 342404 155780
rect 71872 155660 71924 155712
rect 172704 155660 172756 155712
rect 176292 155660 176344 155712
rect 253388 155660 253440 155712
rect 289728 155660 289780 155712
rect 340052 155660 340104 155712
rect 33140 155592 33192 155644
rect 60004 155592 60056 155644
rect 75184 155592 75236 155644
rect 176384 155592 176436 155644
rect 177120 155592 177172 155644
rect 254032 155592 254084 155644
rect 267004 155592 267056 155644
rect 321744 155592 321796 155644
rect 39856 155524 39908 155576
rect 71780 155524 71832 155576
rect 78588 155524 78640 155576
rect 178960 155524 179012 155576
rect 179512 155524 179564 155576
rect 255872 155524 255924 155576
rect 263600 155524 263652 155576
rect 320180 155524 320232 155576
rect 340972 155524 341024 155576
rect 378140 155524 378192 155576
rect 28908 155456 28960 155508
rect 56508 155456 56560 155508
rect 62580 155456 62632 155508
rect 165712 155456 165764 155508
rect 169392 155456 169444 155508
rect 248236 155456 248288 155508
rect 260288 155456 260340 155508
rect 317604 155456 317656 155508
rect 333428 155456 333480 155508
rect 373448 155456 373500 155508
rect 7932 155388 7984 155440
rect 124680 155388 124732 155440
rect 134064 155388 134116 155440
rect 137560 155388 137612 155440
rect 149244 155388 149296 155440
rect 232872 155388 232924 155440
rect 253572 155388 253624 155440
rect 312452 155388 312504 155440
rect 330116 155388 330168 155440
rect 370872 155388 370924 155440
rect 8760 155320 8812 155372
rect 125692 155320 125744 155372
rect 145840 155320 145892 155372
rect 229192 155320 229244 155372
rect 250168 155320 250220 155372
rect 309876 155320 309928 155372
rect 316592 155320 316644 155372
rect 360660 155320 360712 155372
rect 4528 155252 4580 155304
rect 122012 155252 122064 155304
rect 142528 155252 142580 155304
rect 227812 155252 227864 155304
rect 243452 155252 243504 155304
rect 304724 155252 304776 155304
rect 306564 155252 306616 155304
rect 352472 155252 352524 155304
rect 373816 155252 373868 155304
rect 403164 155252 403216 155304
rect 5356 155184 5408 155236
rect 123024 155184 123076 155236
rect 129004 155184 129056 155236
rect 217416 155184 217468 155236
rect 236736 155184 236788 155236
rect 299664 155184 299716 155236
rect 303160 155184 303212 155236
rect 350356 155184 350408 155236
rect 367100 155184 367152 155236
rect 399024 155184 399076 155236
rect 401600 155184 401652 155236
rect 425520 155184 425572 155236
rect 53380 155116 53432 155168
rect 76932 155116 76984 155168
rect 86132 155116 86184 155168
rect 183560 155116 183612 155168
rect 186688 155116 186740 155168
rect 95424 155048 95476 155100
rect 186320 155048 186372 155100
rect 186504 155048 186556 155100
rect 191748 155048 191800 155100
rect 192944 155116 192996 155168
rect 266268 155116 266320 155168
rect 309968 155116 310020 155168
rect 355508 155116 355560 155168
rect 194968 155048 195020 155100
rect 196348 155048 196400 155100
rect 268844 155048 268896 155100
rect 98736 154980 98788 155032
rect 186228 154980 186280 155032
rect 186596 154980 186648 155032
rect 194324 154980 194376 155032
rect 199660 154980 199712 155032
rect 271420 154980 271472 155032
rect 99564 154912 99616 154964
rect 186320 154912 186372 154964
rect 188252 154912 188304 154964
rect 240692 154912 240744 154964
rect 80244 154844 80296 154896
rect 86868 154844 86920 154896
rect 122288 154844 122340 154896
rect 212264 154844 212316 154896
rect 231768 154844 231820 154896
rect 277124 154844 277176 154896
rect 125784 154776 125836 154828
rect 214840 154776 214892 154828
rect 216772 154776 216824 154828
rect 261392 154776 261444 154828
rect 107292 154708 107344 154760
rect 133328 154708 133380 154760
rect 155960 154708 156012 154760
rect 238024 154708 238076 154760
rect 110512 154640 110564 154692
rect 128360 154640 128412 154692
rect 162676 154640 162728 154692
rect 243084 154640 243136 154692
rect 146208 154572 146260 154624
rect 44180 154504 44232 154556
rect 146484 154504 146536 154556
rect 41604 154436 41656 154488
rect 150624 154504 150676 154556
rect 151820 154572 151872 154624
rect 156604 154504 156656 154556
rect 159364 154572 159416 154624
rect 240140 154572 240192 154624
rect 156788 154504 156840 154556
rect 157340 154504 157392 154556
rect 225788 154504 225840 154556
rect 231860 154504 231912 154556
rect 296444 154504 296496 154556
rect 353668 154504 353720 154556
rect 388904 154504 388956 154556
rect 34520 154368 34572 154420
rect 145380 154368 145432 154420
rect 37924 154300 37976 154352
rect 145104 154300 145156 154352
rect 30380 154232 30432 154284
rect 137100 154232 137152 154284
rect 185124 154436 185176 154488
rect 191288 154436 191340 154488
rect 200120 154436 200172 154488
rect 218336 154436 218388 154488
rect 285588 154436 285640 154488
rect 285680 154436 285732 154488
rect 337476 154436 337528 154488
rect 356244 154436 356296 154488
rect 391480 154436 391532 154488
rect 400312 154436 400364 154488
rect 424876 154436 424928 154488
rect 23480 154164 23532 154216
rect 137008 154164 137060 154216
rect 13820 154096 13872 154148
rect 126796 154096 126848 154148
rect 188436 154368 188488 154420
rect 191472 154368 191524 154420
rect 202696 154368 202748 154420
rect 208400 154368 208452 154420
rect 278412 154368 278464 154420
rect 278872 154368 278924 154420
rect 332416 154368 332468 154420
rect 349528 154368 349580 154420
rect 386328 154368 386380 154420
rect 397460 154368 397512 154420
rect 423036 154368 423088 154420
rect 146944 154300 146996 154352
rect 191288 154300 191340 154352
rect 191380 154300 191432 154352
rect 202052 154300 202104 154352
rect 204812 154300 204864 154352
rect 275836 154300 275888 154352
rect 276204 154300 276256 154352
rect 329932 154300 329984 154352
rect 346400 154300 346452 154352
rect 383752 154300 383804 154352
rect 390652 154300 390704 154352
rect 417148 154300 417200 154352
rect 9680 154028 9732 154080
rect 126888 154028 126940 154080
rect 7104 153960 7156 154012
rect 117964 153960 118016 154012
rect 2964 153892 3016 153944
rect 121736 153960 121788 154012
rect 121828 153960 121880 154012
rect 118148 153892 118200 153944
rect 124312 153892 124364 153944
rect 125508 153892 125560 153944
rect 127900 153960 127952 154012
rect 146852 154096 146904 154148
rect 137468 154028 137520 154080
rect 137652 154028 137704 154080
rect 185216 154232 185268 154284
rect 185308 154232 185360 154284
rect 258540 154232 258592 154284
rect 262220 154232 262272 154284
rect 319536 154232 319588 154284
rect 336832 154232 336884 154284
rect 376024 154232 376076 154284
rect 393320 154232 393372 154284
rect 419724 154232 419776 154284
rect 147128 154164 147180 154216
rect 152740 154164 152792 154216
rect 153292 154164 153344 154216
rect 163504 154164 163556 154216
rect 165068 154164 165120 154216
rect 168656 154164 168708 154216
rect 172520 154164 172572 154216
rect 250812 154164 250864 154216
rect 255320 154164 255372 154216
rect 314384 154164 314436 154216
rect 342812 154164 342864 154216
rect 381176 154164 381228 154216
rect 386512 154164 386564 154216
rect 414572 154164 414624 154216
rect 147036 154096 147088 154148
rect 142344 153960 142396 154012
rect 145104 153960 145156 154012
rect 148140 154028 148192 154080
rect 150072 154096 150124 154148
rect 152648 154028 152700 154080
rect 155776 154028 155828 154080
rect 153200 153960 153252 154012
rect 156880 154096 156932 154148
rect 166264 154096 166316 154148
rect 166356 154096 166408 154148
rect 245660 154096 245712 154148
rect 248604 154096 248656 154148
rect 309232 154096 309284 154148
rect 326712 154096 326764 154148
rect 368296 154096 368348 154148
rect 383660 154096 383712 154148
rect 411996 154096 412048 154148
rect 156788 154028 156840 154080
rect 235448 154028 235500 154080
rect 241888 154028 241940 154080
rect 304080 154028 304132 154080
rect 323308 154028 323360 154080
rect 365812 154028 365864 154080
rect 376852 154028 376904 154080
rect 406844 154028 406896 154080
rect 233516 153960 233568 154012
rect 235080 153960 235132 154012
rect 299020 153960 299072 154012
rect 319260 153960 319312 154012
rect 363236 153960 363288 154012
rect 369952 153960 370004 154012
rect 401600 153960 401652 154012
rect 127164 153892 127216 153944
rect 129464 153892 129516 153944
rect 129924 153892 129976 153944
rect 218060 153892 218112 153944
rect 225052 153892 225104 153944
rect 291384 153892 291436 153944
rect 313280 153892 313332 153944
rect 357808 153892 357860 153944
rect 360384 153892 360436 153944
rect 394056 153892 394108 153944
rect 397368 153892 397420 153944
rect 422484 153892 422536 153944
rect 480 153824 532 153876
rect 119804 153824 119856 153876
rect 119896 153824 119948 153876
rect 209780 153824 209832 153876
rect 215300 153824 215352 153876
rect 283656 153824 283708 153876
rect 285680 153824 285732 153876
rect 286140 153824 286192 153876
rect 286232 153824 286284 153876
rect 334900 153824 334952 153876
rect 339500 153824 339552 153876
rect 378600 153824 378652 153876
rect 380164 153824 380216 153876
rect 409420 153824 409472 153876
rect 48320 153756 48372 153808
rect 152648 153756 152700 153808
rect 152740 153756 152792 153808
rect 212908 153756 212960 153808
rect 222384 153756 222436 153808
rect 288716 153756 288768 153808
rect 363052 153756 363104 153808
rect 396540 153756 396592 153808
rect 426440 153756 426492 153808
rect 432420 153756 432472 153808
rect 57980 153688 58032 153740
rect 153292 153688 153344 153740
rect 154488 153688 154540 153740
rect 156512 153688 156564 153740
rect 156604 153688 156656 153740
rect 210424 153688 210476 153740
rect 229100 153688 229152 153740
rect 293868 153688 293920 153740
rect 64880 153620 64932 153672
rect 165068 153620 165120 153672
rect 166264 153620 166316 153672
rect 215484 153620 215536 153672
rect 238852 153620 238904 153672
rect 301596 153620 301648 153672
rect 82820 153552 82872 153604
rect 182088 153552 182140 153604
rect 182180 153552 182232 153604
rect 185032 153552 185084 153604
rect 185124 153552 185176 153604
rect 188344 153552 188396 153604
rect 188436 153552 188488 153604
rect 197544 153552 197596 153604
rect 102140 153484 102192 153536
rect 196900 153484 196952 153536
rect 196992 153484 197044 153536
rect 243728 153552 243780 153604
rect 245936 153552 245988 153604
rect 306656 153552 306708 153604
rect 198924 153484 198976 153536
rect 248880 153484 248932 153536
rect 252652 153484 252704 153536
rect 311808 153484 311860 153536
rect 331220 153484 331272 153536
rect 337016 153484 337068 153536
rect 104900 153416 104952 153468
rect 199476 153416 199528 153468
rect 201408 153416 201460 153468
rect 256608 153416 256660 153468
rect 265440 153416 265492 153468
rect 322204 153416 322256 153468
rect 108304 153348 108356 153400
rect 191380 153348 191432 153400
rect 194508 153348 194560 153400
rect 238668 153348 238720 153400
rect 259460 153348 259512 153400
rect 316960 153348 317012 153400
rect 437572 153348 437624 153400
rect 114836 153280 114888 153332
rect 118608 153280 118660 153332
rect 118792 153280 118844 153332
rect 119896 153280 119948 153332
rect 119988 153280 120040 153332
rect 207204 153280 207256 153332
rect 272892 153280 272944 153332
rect 327264 153280 327316 153332
rect 425980 153280 426032 153332
rect 431316 153280 431368 153332
rect 115940 153212 115992 153264
rect 207848 153212 207900 153264
rect 269212 153212 269264 153264
rect 324688 153212 324740 153264
rect 120080 153144 120132 153196
rect 205916 153144 205968 153196
rect 223856 153144 223908 153196
rect 288072 153144 288124 153196
rect 288256 153144 288308 153196
rect 290004 153144 290056 153196
rect 303712 153144 303764 153196
rect 351000 153144 351052 153196
rect 352012 153144 352064 153196
rect 388260 153144 388312 153196
rect 389180 153144 389232 153196
rect 412640 153144 412692 153196
rect 413100 153144 413152 153196
rect 428096 153212 428148 153264
rect 431868 153212 431920 153264
rect 427912 153144 427964 153196
rect 432696 153144 432748 153196
rect 433800 153144 433852 153196
rect 434352 153144 434404 153196
rect 86868 153076 86920 153128
rect 180248 153076 180300 153128
rect 180800 153076 180852 153128
rect 257252 153076 257304 153128
rect 264980 153076 265032 153128
rect 321468 153076 321520 153128
rect 324228 153076 324280 153128
rect 366364 153076 366416 153128
rect 368480 153076 368532 153128
rect 400404 153076 400456 153128
rect 403256 153076 403308 153128
rect 415860 153076 415912 153128
rect 419264 153076 419316 153128
rect 432788 153076 432840 153128
rect 436100 153076 436152 153128
rect 437572 153076 437624 153128
rect 437848 153144 437900 153196
rect 438400 153144 438452 153196
rect 440240 153144 440292 153196
rect 440516 153144 440568 153196
rect 441988 153212 442040 153264
rect 442172 153144 442224 153196
rect 449256 153144 449308 153196
rect 453856 153144 453908 153196
rect 459468 153144 459520 153196
rect 461860 153144 461912 153196
rect 465908 153144 465960 153196
rect 466460 153144 466512 153196
rect 469772 153144 469824 153196
rect 471428 153144 471480 153196
rect 472992 153144 473044 153196
rect 473360 153144 473412 153196
rect 475568 153144 475620 153196
rect 476120 153144 476172 153196
rect 478144 153144 478196 153196
rect 485688 153144 485740 153196
rect 489644 153144 489696 153196
rect 490748 153144 490800 153196
rect 493508 153144 493560 153196
rect 494060 153144 494112 153196
rect 496084 153144 496136 153196
rect 496636 153144 496688 153196
rect 498016 153144 498068 153196
rect 512920 153144 512972 153196
rect 515220 153144 515272 153196
rect 103520 153008 103572 153060
rect 198188 153008 198240 153060
rect 215392 153008 215444 153060
rect 279700 153008 279752 153060
rect 291476 153008 291528 153060
rect 335728 153008 335780 153060
rect 96620 152940 96672 152992
rect 193036 152940 193088 152992
rect 203708 152940 203760 152992
rect 267556 152940 267608 152992
rect 272156 152940 272208 152992
rect 320732 152940 320784 152992
rect 330944 152940 330996 152992
rect 336096 153008 336148 153060
rect 347136 153008 347188 153060
rect 349160 153008 349212 153060
rect 385592 153008 385644 153060
rect 386236 153008 386288 153060
rect 399760 153008 399812 153060
rect 406660 153008 406712 153060
rect 429292 153008 429344 153060
rect 371516 152940 371568 152992
rect 372620 152940 372672 152992
rect 403624 152940 403676 152992
rect 404360 152940 404412 152992
rect 427636 152940 427688 152992
rect 428096 152940 428148 152992
rect 431868 153008 431920 153060
rect 431960 153008 432012 153060
rect 441988 153008 442040 153060
rect 442540 153076 442592 153128
rect 443552 153076 443604 153128
rect 444472 153076 444524 153128
rect 458272 153076 458324 153128
rect 462964 153076 463016 153128
rect 467288 153076 467340 153128
rect 471244 153076 471296 153128
rect 473636 153076 473688 153128
rect 474832 153076 474884 153128
rect 476948 153076 477000 153128
rect 484032 153076 484084 153128
rect 488448 153076 488500 153128
rect 489920 153076 489972 153128
rect 492864 153076 492916 153128
rect 494152 153076 494204 153128
rect 496728 153076 496780 153128
rect 496820 153076 496872 153128
rect 498660 153076 498712 153128
rect 510988 153076 511040 153128
rect 513472 153076 513524 153128
rect 514208 153076 514260 153128
rect 517428 153076 517480 153128
rect 442264 153008 442316 153060
rect 430580 152940 430632 152992
rect 442356 152940 442408 152992
rect 89812 152872 89864 152924
rect 187884 152872 187936 152924
rect 191656 152872 191708 152924
rect 208492 152872 208544 152924
rect 212448 152872 212500 152924
rect 277768 152872 277820 152924
rect 285496 152872 285548 152924
rect 335820 152872 335872 152924
rect 335912 152872 335964 152924
rect 341340 152872 341392 152924
rect 341432 152872 341484 152924
rect 377312 152872 377364 152924
rect 378232 152872 378284 152924
rect 379888 152872 379940 152924
rect 380900 152872 380952 152924
rect 410064 152872 410116 152924
rect 411260 152872 411312 152924
rect 433156 152872 433208 152924
rect 433524 152872 433576 152924
rect 449900 153008 449952 153060
rect 456892 153008 456944 153060
rect 460756 153008 460808 153060
rect 463516 153008 463568 153060
rect 466552 153008 466604 153060
rect 466644 153008 466696 153060
rect 470416 153008 470468 153060
rect 472348 153008 472400 153060
rect 474924 153008 474976 153060
rect 484492 153008 484544 153060
rect 489000 153008 489052 153060
rect 492680 153008 492732 153060
rect 495440 153008 495492 153060
rect 495532 153008 495584 153060
rect 497372 153008 497424 153060
rect 442540 152940 442592 152992
rect 447968 152940 448020 152992
rect 463884 152940 463936 152992
rect 468392 152940 468444 152992
rect 472440 152940 472492 152992
rect 474280 152940 474332 152992
rect 483112 152940 483164 152992
rect 487804 152940 487856 152992
rect 491668 152940 491720 152992
rect 494796 152940 494848 152992
rect 512276 152940 512328 152992
rect 514760 152940 514812 152992
rect 443184 152872 443236 152924
rect 451188 152872 451240 152924
rect 459652 152872 459704 152924
rect 464620 152872 464672 152924
rect 465080 152872 465132 152924
rect 469128 152872 469180 152924
rect 491300 152872 491352 152924
rect 494152 152872 494204 152924
rect 513564 152872 513616 152924
rect 516140 152872 516192 152924
rect 66260 152804 66312 152856
rect 169944 152804 169996 152856
rect 173900 152804 173952 152856
rect 252100 152804 252152 152856
rect 257712 152804 257764 152856
rect 315672 152804 315724 152856
rect 317052 152804 317104 152856
rect 318248 152804 318300 152856
rect 318340 152804 318392 152856
rect 361948 152804 362000 152856
rect 365720 152804 365772 152856
rect 367008 152804 367060 152856
rect 367192 152804 367244 152856
rect 368940 152804 368992 152856
rect 369032 152804 369084 152856
rect 397184 152804 397236 152856
rect 401692 152804 401744 152856
rect 426164 152804 426216 152856
rect 426348 152804 426400 152856
rect 26424 152736 26476 152788
rect 139124 152736 139176 152788
rect 139400 152736 139452 152788
rect 141700 152736 141752 152788
rect 22192 152668 22244 152720
rect 135904 152668 135956 152720
rect 146852 152736 146904 152788
rect 149060 152736 149112 152788
rect 231584 152736 231636 152788
rect 240324 152736 240376 152788
rect 241888 152736 241940 152788
rect 244372 152736 244424 152788
rect 306012 152736 306064 152788
rect 307668 152736 307720 152788
rect 352288 152736 352340 152788
rect 357440 152736 357492 152788
rect 359372 152736 359424 152788
rect 359464 152736 359516 152788
rect 390192 152736 390244 152788
rect 15200 152600 15252 152652
rect 130752 152600 130804 152652
rect 135168 152600 135220 152652
rect 141884 152668 141936 152720
rect 151912 152668 151964 152720
rect 153568 152668 153620 152720
rect 236736 152668 236788 152720
rect 247040 152668 247092 152720
rect 307944 152668 307996 152720
rect 311532 152668 311584 152720
rect 356796 152668 356848 152720
rect 358820 152668 358872 152720
rect 393412 152668 393464 152720
rect 136916 152600 136968 152652
rect 137192 152600 137244 152652
rect 19340 152532 19392 152584
rect 133972 152532 134024 152584
rect 2872 152464 2924 152516
rect 121092 152464 121144 152516
rect 129740 152464 129792 152516
rect 216128 152600 216180 152652
rect 220452 152600 220504 152652
rect 284852 152600 284904 152652
rect 285772 152600 285824 152652
rect 291844 152600 291896 152652
rect 292212 152600 292264 152652
rect 341984 152600 342036 152652
rect 342260 152600 342312 152652
rect 343916 152600 343968 152652
rect 345296 152600 345348 152652
rect 382464 152600 382516 152652
rect 386420 152600 386472 152652
rect 140780 152532 140832 152584
rect 137560 152464 137612 152516
rect 141148 152464 141200 152516
rect 146944 152532 146996 152584
rect 221280 152532 221332 152584
rect 225236 152532 225288 152584
rect 229008 152532 229060 152584
rect 234160 152532 234212 152584
rect 297732 152532 297784 152584
rect 304816 152532 304868 152584
rect 351644 152532 351696 152584
rect 354496 152532 354548 152584
rect 389548 152532 389600 152584
rect 390376 152600 390428 152652
rect 415216 152736 415268 152788
rect 415400 152736 415452 152788
rect 427820 152736 427872 152788
rect 395528 152668 395580 152720
rect 397828 152668 397880 152720
rect 399116 152668 399168 152720
rect 424232 152668 424284 152720
rect 413928 152600 413980 152652
rect 414388 152600 414440 152652
rect 430028 152736 430080 152788
rect 430212 152804 430264 152856
rect 447324 152804 447376 152856
rect 510344 152804 510396 152856
rect 512000 152804 512052 152856
rect 434536 152736 434588 152788
rect 434720 152736 434772 152788
rect 428188 152668 428240 152720
rect 438860 152736 438912 152788
rect 454408 152736 454460 152788
rect 511632 152736 511684 152788
rect 513748 152736 513800 152788
rect 394884 152532 394936 152584
rect 420368 152532 420420 152584
rect 423404 152532 423456 152584
rect 437112 152600 437164 152652
rect 440240 152668 440292 152720
rect 440332 152668 440384 152720
rect 445484 152668 445536 152720
rect 441436 152600 441488 152652
rect 441620 152600 441672 152652
rect 444748 152600 444800 152652
rect 459560 152600 459612 152652
rect 465264 152600 465316 152652
rect 429844 152532 429896 152584
rect 441528 152532 441580 152584
rect 442080 152532 442132 152584
rect 444656 152532 444708 152584
rect 445576 152532 445628 152584
rect 456984 152532 457036 152584
rect 458180 152532 458232 152584
rect 463976 152532 464028 152584
rect 226432 152464 226484 152516
rect 227904 152464 227956 152516
rect 293224 152464 293276 152516
rect 298652 152464 298704 152516
rect 335912 152464 335964 152516
rect 336004 152464 336056 152516
rect 346492 152464 346544 152516
rect 347964 152464 348016 152516
rect 385040 152464 385092 152516
rect 385316 152464 385368 152516
rect 387616 152464 387668 152516
rect 393136 152464 393188 152516
rect 419080 152464 419132 152516
rect 421196 152464 421248 152516
rect 432604 152464 432656 152516
rect 432696 152464 432748 152516
rect 60004 152396 60056 152448
rect 144276 152396 144328 152448
rect 144828 152396 144880 152448
rect 162216 152396 162268 152448
rect 164332 152396 164384 152448
rect 244372 152396 244424 152448
rect 251180 152396 251232 152448
rect 311164 152396 311216 152448
rect 311992 152396 312044 152448
rect 356152 152396 356204 152448
rect 361580 152396 361632 152448
rect 395344 152396 395396 152448
rect 398840 152396 398892 152448
rect 413284 152396 413336 152448
rect 413836 152396 413888 152448
rect 416504 152396 416556 152448
rect 418436 152396 418488 152448
rect 113180 152328 113232 152380
rect 120080 152328 120132 152380
rect 120172 152328 120224 152380
rect 211068 152328 211120 152380
rect 221740 152328 221792 152380
rect 282920 152328 282972 152380
rect 283196 152328 283248 152380
rect 287428 152328 287480 152380
rect 291844 152328 291896 152380
rect 336188 152328 336240 152380
rect 343640 152328 343692 152380
rect 380532 152328 380584 152380
rect 381452 152328 381504 152380
rect 410708 152328 410760 152380
rect 413192 152328 413244 152380
rect 421656 152328 421708 152380
rect 425152 152328 425204 152380
rect 430028 152396 430080 152448
rect 435732 152396 435784 152448
rect 436192 152464 436244 152516
rect 444564 152464 444616 152516
rect 445484 152464 445536 152516
rect 455696 152464 455748 152516
rect 436376 152396 436428 152448
rect 437480 152396 437532 152448
rect 444472 152396 444524 152448
rect 56508 152260 56560 152312
rect 141056 152260 141108 152312
rect 141148 152260 141200 152312
rect 146944 152260 146996 152312
rect 150440 152260 150492 152312
rect 167368 152260 167420 152312
rect 172612 152260 172664 152312
rect 249524 152260 249576 152312
rect 255504 152260 255556 152312
rect 313096 152260 313148 152312
rect 320272 152260 320324 152312
rect 323124 152260 323176 152312
rect 76932 152192 76984 152244
rect 159640 152192 159692 152244
rect 160192 152192 160244 152244
rect 177672 152192 177724 152244
rect 187976 152192 188028 152244
rect 262404 152192 262456 152244
rect 266360 152192 266412 152244
rect 320824 152192 320876 152244
rect 320916 152192 320968 152244
rect 361304 152260 361356 152312
rect 364524 152260 364576 152312
rect 369032 152260 369084 152312
rect 324320 152192 324372 152244
rect 367008 152192 367060 152244
rect 367100 152192 367152 152244
rect 398472 152260 398524 152312
rect 398564 152260 398616 152312
rect 408132 152260 408184 152312
rect 410892 152260 410944 152312
rect 438308 152328 438360 152380
rect 438400 152328 438452 152380
rect 453764 152396 453816 152448
rect 445116 152328 445168 152380
rect 456340 152328 456392 152380
rect 371332 152192 371384 152244
rect 402336 152192 402388 152244
rect 405832 152192 405884 152244
rect 408776 152192 408828 152244
rect 409236 152192 409288 152244
rect 426716 152192 426768 152244
rect 84752 152124 84804 152176
rect 164792 152124 164844 152176
rect 167000 152124 167052 152176
rect 182732 152124 182784 152176
rect 192668 152124 192720 152176
rect 213552 152124 213604 152176
rect 213828 152124 213880 152176
rect 274548 152124 274600 152176
rect 278780 152124 278832 152176
rect 331772 152124 331824 152176
rect 335820 152124 335872 152176
rect 336832 152124 336884 152176
rect 336924 152124 336976 152176
rect 372804 152124 372856 152176
rect 384948 152124 385000 152176
rect 392124 152124 392176 152176
rect 394332 152124 394384 152176
rect 417792 152124 417844 152176
rect 419632 152124 419684 152176
rect 427728 152124 427780 152176
rect 432696 152260 432748 152312
rect 432788 152260 432840 152312
rect 438952 152260 439004 152312
rect 440516 152260 440568 152312
rect 455052 152260 455104 152312
rect 455512 152260 455564 152312
rect 462044 152260 462096 152312
rect 429384 152192 429436 152244
rect 446680 152192 446732 152244
rect 456800 152192 456852 152244
rect 463332 152192 463384 152244
rect 431224 152124 431276 152176
rect 431316 152124 431368 152176
rect 444104 152124 444156 152176
rect 75828 152056 75880 152108
rect 154488 152056 154540 152108
rect 156052 152056 156104 152108
rect 172520 152056 172572 152108
rect 185584 152056 185636 152108
rect 200764 152056 200816 152108
rect 71780 151988 71832 152040
rect 149428 151988 149480 152040
rect 169760 151988 169812 152040
rect 185308 151988 185360 152040
rect 195152 151988 195204 152040
rect 218704 151988 218756 152040
rect 109040 151920 109092 151972
rect 128176 151920 128228 151972
rect 128360 151920 128412 151972
rect 203340 151920 203392 151972
rect 212724 151920 212776 151972
rect 272708 152056 272760 152108
rect 272800 152056 272852 152108
rect 325976 152056 326028 152108
rect 335360 152056 335412 152108
rect 375380 152056 375432 152108
rect 382280 152056 382332 152108
rect 386972 152056 387024 152108
rect 388352 152056 388404 152108
rect 407488 152056 407540 152108
rect 408500 152056 408552 152108
rect 423588 152056 423640 152108
rect 423680 152056 423732 152108
rect 426348 152056 426400 152108
rect 432420 152056 432472 152108
rect 444748 152056 444800 152108
rect 242808 151988 242860 152040
rect 300952 151988 301004 152040
rect 301044 151988 301096 152040
rect 336004 151988 336056 152040
rect 243360 151920 243412 151972
rect 302884 151920 302936 151972
rect 317420 151920 317472 151972
rect 320916 151920 320968 151972
rect 321560 151920 321612 151972
rect 325608 151920 325660 151972
rect 325884 151920 325936 151972
rect 342444 151988 342496 152040
rect 344560 151988 344612 152040
rect 354680 151988 354732 152040
rect 359464 151988 359516 152040
rect 378784 151988 378836 152040
rect 384396 151988 384448 152040
rect 385776 151988 385828 152040
rect 394700 151988 394752 152040
rect 404728 151988 404780 152040
rect 421012 151988 421064 152040
rect 367652 151920 367704 151972
rect 375472 151920 375524 151972
rect 405556 151920 405608 151972
rect 416596 151920 416648 151972
rect 426808 151988 426860 152040
rect 432696 151988 432748 152040
rect 443460 151988 443512 152040
rect 443552 151988 443604 152040
rect 450544 152124 450596 152176
rect 455880 152124 455932 152176
rect 461400 152124 461452 152176
rect 446312 152056 446364 152108
rect 460112 152056 460164 152108
rect 445300 151988 445352 152040
rect 458824 151988 458876 152040
rect 485780 151988 485832 152040
rect 490288 151988 490340 152040
rect 516692 151988 516744 152040
rect 520280 151988 520332 152040
rect 422576 151920 422628 151972
rect 429844 151920 429896 151972
rect 434536 151920 434588 151972
rect 439596 151920 439648 151972
rect 440240 151920 440292 151972
rect 451096 151920 451148 151972
rect 451188 151920 451240 151972
rect 457628 151920 457680 151972
rect 469220 151920 469272 151972
rect 472348 151920 472400 151972
rect 487344 151920 487396 151972
rect 490932 151920 490984 151972
rect 509056 151920 509108 151972
rect 510896 151920 510948 151972
rect 515496 151920 515548 151972
rect 518992 151920 519044 151972
rect 30196 151852 30248 151904
rect 74540 151852 74592 151904
rect 107568 151852 107620 151904
rect 175096 151852 175148 151904
rect 176660 151852 176712 151904
rect 190460 151852 190512 151904
rect 261024 151852 261076 151904
rect 316316 151852 316368 151904
rect 320732 151852 320784 151904
rect 326620 151852 326672 151904
rect 33600 151784 33652 151836
rect 84200 151784 84252 151836
rect 105820 151784 105872 151836
rect 109776 151784 109828 151836
rect 109868 151784 109920 151836
rect 138480 151784 138532 151836
rect 138572 151784 138624 151836
rect 141884 151784 141936 151836
rect 142252 151784 142304 151836
rect 157064 151784 157116 151836
rect 183100 151784 183152 151836
rect 195612 151784 195664 151836
rect 277400 151784 277452 151836
rect 331128 151852 331180 151904
rect 332600 151852 332652 151904
rect 336924 151852 336976 151904
rect 337016 151852 337068 151904
rect 372160 151852 372212 151904
rect 396172 151852 396224 151904
rect 402980 151852 403032 151904
rect 404268 151852 404320 151904
rect 418436 151852 418488 151904
rect 419540 151852 419592 151904
rect 437020 151852 437072 151904
rect 437112 151852 437164 151904
rect 442172 151852 442224 151904
rect 442264 151852 442316 151904
rect 325608 151716 325660 151768
rect 362592 151784 362644 151836
rect 363144 151784 363196 151836
rect 364524 151784 364576 151836
rect 388444 151784 388496 151836
rect 404912 151784 404964 151836
rect 417424 151784 417476 151836
rect 431868 151784 431920 151836
rect 432604 151784 432656 151836
rect 440884 151784 440936 151836
rect 441436 151784 441488 151836
rect 444840 151852 444892 151904
rect 452476 151852 452528 151904
rect 467840 151852 467892 151904
rect 471060 151852 471112 151904
rect 488540 151852 488592 151904
rect 492220 151852 492272 151904
rect 507768 151852 507820 151904
rect 509516 151852 509568 151904
rect 516048 151852 516100 151904
rect 519912 151852 519964 151904
rect 451832 151784 451884 151836
rect 457168 151784 457220 151836
rect 462688 151784 462740 151836
rect 464344 151784 464396 151836
rect 467748 151784 467800 151836
rect 467932 151784 467984 151836
rect 471704 151784 471756 151836
rect 488172 151784 488224 151836
rect 491576 151784 491628 151836
rect 499120 151784 499172 151836
rect 499948 151784 500000 151836
rect 517428 151784 517480 151836
rect 521568 151784 521620 151836
rect 446036 151648 446088 151700
rect 84200 151376 84252 151428
rect 117228 151376 117280 151428
rect 74540 151308 74592 151360
rect 117136 151308 117188 151360
rect 68008 151240 68060 151292
rect 112812 151240 112864 151292
rect 64512 151172 64564 151224
rect 112720 151172 112772 151224
rect 61108 151104 61160 151156
rect 112628 151104 112680 151156
rect 57704 151036 57756 151088
rect 112536 151036 112588 151088
rect 54208 150968 54260 151020
rect 111616 150968 111668 151020
rect 50804 150900 50856 150952
rect 112444 150900 112496 150952
rect 47308 150832 47360 150884
rect 111524 150832 111576 150884
rect 43904 150764 43956 150816
rect 111432 150764 111484 150816
rect 40500 150696 40552 150748
rect 111340 150696 111392 150748
rect 37004 150628 37056 150680
rect 111248 150628 111300 150680
rect 19800 150560 19852 150612
rect 116860 150560 116912 150612
rect 16396 150492 16448 150544
rect 116768 150492 116820 150544
rect 2688 150424 2740 150476
rect 111064 150424 111116 150476
rect 263692 150288 263744 150340
rect 122840 150152 122892 150204
rect 123714 150152 123766 150204
rect 146392 150152 146444 150204
rect 147542 150152 147594 150204
rect 147680 150152 147732 150204
rect 148830 150152 148882 150204
rect 165712 150152 165764 150204
rect 166770 150152 166822 150204
rect 171140 150152 171192 150204
rect 171922 150152 171974 150204
rect 172704 150152 172756 150204
rect 173854 150152 173906 150204
rect 182272 150152 182324 150204
rect 183422 150152 183474 150204
rect 183560 150152 183612 150204
rect 184710 150152 184762 150204
rect 200304 150152 200356 150204
rect 201454 150152 201506 150204
rect 219532 150152 219584 150204
rect 220682 150152 220734 150204
rect 222292 150152 222344 150204
rect 223258 150152 223310 150204
rect 229192 150152 229244 150204
rect 230342 150152 230394 150204
rect 238944 150152 238996 150204
rect 240002 150152 240054 150204
rect 253940 150152 253992 150204
rect 254722 150152 254774 150204
rect 256792 150152 256844 150204
rect 257942 150152 257994 150204
rect 258080 150152 258132 150204
rect 259230 150152 259282 150204
rect 264382 150152 264434 150204
rect 269120 150152 269172 150204
rect 270178 150152 270230 150204
rect 281540 150152 281592 150204
rect 282322 150152 282374 150204
rect 283104 150152 283156 150204
rect 284254 150152 284306 150204
rect 284392 150152 284444 150204
rect 285542 150152 285594 150204
rect 299480 150152 299532 150204
rect 300354 150152 300406 150204
rect 321744 150152 321796 150204
rect 322802 150152 322854 150204
rect 338396 150152 338448 150204
rect 339454 150152 339506 150204
rect 345112 150152 345164 150204
rect 345894 150152 345946 150204
rect 358912 150152 358964 150204
rect 360062 150152 360114 150204
rect 362960 150152 363012 150204
rect 363926 150152 363978 150204
rect 374000 150152 374052 150204
rect 374782 150152 374834 150204
rect 378140 150152 378192 150204
rect 379290 150152 379342 150204
rect 403164 150152 403216 150204
rect 404314 150152 404366 150204
rect 426716 150152 426768 150204
rect 428694 150152 428746 150204
rect 444472 150152 444524 150204
rect 453166 150152 453218 150204
rect 477684 150152 477736 150204
rect 478834 150152 478886 150204
rect 478972 150152 479024 150204
rect 480122 150152 480174 150204
rect 481640 150152 481692 150204
rect 482698 150152 482750 150204
rect 483204 150152 483256 150204
rect 483986 150152 484038 150204
rect 505284 150152 505336 150204
rect 506434 150152 506486 150204
rect 518026 150152 518078 150204
rect 518808 150152 518860 150204
rect 427728 150084 427780 150136
rect 434490 150084 434542 150136
rect 6368 150016 6420 150068
rect 111156 150016 111208 150068
rect 23388 149948 23440 150000
rect 116952 149948 117004 150000
rect 13360 149880 13412 149932
rect 116676 149880 116728 149932
rect 9588 149812 9640 149864
rect 116584 149812 116636 149864
rect 88984 149744 89036 149796
rect 114008 149744 114060 149796
rect 85488 149676 85540 149728
rect 113916 149676 113968 149728
rect 81992 149608 82044 149660
rect 112352 149608 112404 149660
rect 78588 149540 78640 149592
rect 113088 149540 113140 149592
rect 75184 149472 75236 149524
rect 112996 149472 113048 149524
rect 71688 149404 71740 149456
rect 112904 149404 112956 149456
rect 26976 149336 27028 149388
rect 117044 149336 117096 149388
rect 92296 149268 92348 149320
rect 95792 149268 95844 149320
rect 105268 149268 105320 149320
rect 116216 149268 116268 149320
rect 116492 149200 116544 149252
rect 109684 149132 109736 149184
rect 116032 149132 116084 149184
rect 114100 149064 114152 149116
rect 109592 148996 109644 149048
rect 116124 148996 116176 149048
rect 109776 147568 109828 147620
rect 116124 147568 116176 147620
rect 114100 140700 114152 140752
rect 116400 140700 116452 140752
rect 114008 137912 114060 137964
rect 116216 137912 116268 137964
rect 113916 136552 113968 136604
rect 116400 136552 116452 136604
rect 112352 133832 112404 133884
rect 116124 133832 116176 133884
rect 113088 132404 113140 132456
rect 116124 132404 116176 132456
rect 112996 131044 113048 131096
rect 116124 131044 116176 131096
rect 112904 128256 112956 128308
rect 116124 128256 116176 128308
rect 112812 126896 112864 126948
rect 116124 126896 116176 126948
rect 112720 124108 112772 124160
rect 116124 124108 116176 124160
rect 112628 122748 112680 122800
rect 116124 122748 116176 122800
rect 112536 121388 112588 121440
rect 116124 121388 116176 121440
rect 111616 118600 111668 118652
rect 116124 118600 116176 118652
rect 112444 117240 112496 117292
rect 116124 117240 116176 117292
rect 111524 114452 111576 114504
rect 116124 114452 116176 114504
rect 111432 113092 111484 113144
rect 116124 113092 116176 113144
rect 111340 111732 111392 111784
rect 116124 111732 116176 111784
rect 111248 108944 111300 108996
rect 116124 108944 116176 108996
rect 111156 92420 111208 92472
rect 115940 92420 115992 92472
rect 111064 89632 111116 89684
rect 116124 89632 116176 89684
rect 113824 88272 113876 88324
rect 115940 88272 115992 88324
rect 114468 86980 114520 87032
rect 116676 86980 116728 87032
rect 113916 86912 113968 86964
rect 116032 86912 116084 86964
rect 114008 83920 114060 83972
rect 116584 83920 116636 83972
rect 114100 82764 114152 82816
rect 116124 82764 116176 82816
rect 114192 79976 114244 80028
rect 115940 79976 115992 80028
rect 114192 71748 114244 71800
rect 116032 71748 116084 71800
rect 114100 69028 114152 69080
rect 116216 69028 116268 69080
rect 114008 67600 114060 67652
rect 115940 67600 115992 67652
rect 113916 66240 113968 66292
rect 116584 66240 116636 66292
rect 114468 64676 114520 64728
rect 116584 64676 116636 64728
rect 113824 63520 113876 63572
rect 116032 63520 116084 63572
rect 109684 41420 109736 41472
rect 116124 41420 116176 41472
rect 114100 38632 114152 38684
rect 116400 38632 116452 38684
rect 116216 38496 116268 38548
rect 116400 38496 116452 38548
rect 114192 37272 114244 37324
rect 115940 37272 115992 37324
rect 111064 34484 111116 34536
rect 116124 34484 116176 34536
rect 112444 33124 112496 33176
rect 116124 33124 116176 33176
rect 112536 31764 112588 31816
rect 116124 31764 116176 31816
rect 112628 28976 112680 29028
rect 116124 28976 116176 29028
rect 112720 27616 112772 27668
rect 116124 27616 116176 27668
rect 112812 24828 112864 24880
rect 116124 24828 116176 24880
rect 111156 23468 111208 23520
rect 116124 23468 116176 23520
rect 111248 22108 111300 22160
rect 116124 22108 116176 22160
rect 109776 4156 109828 4208
rect 115940 4156 115992 4208
rect 2504 2864 2556 2916
rect 40684 2592 40736 2644
rect 43628 2592 43680 2644
rect 45652 2592 45704 2644
rect 49608 2592 49660 2644
rect 49792 2592 49844 2644
rect 49884 2592 49936 2644
rect 49976 2592 50028 2644
rect 53932 2592 53984 2644
rect 58992 2592 59044 2644
rect 32772 2524 32824 2576
rect 59728 2592 59780 2644
rect 59820 2592 59872 2644
rect 40684 2456 40736 2508
rect 39672 2388 39724 2440
rect 53656 2388 53708 2440
rect 36360 2320 36412 2372
rect 43628 2320 43680 2372
rect 46296 2320 46348 2372
rect 49792 2320 49844 2372
rect 56232 2388 56284 2440
rect 64880 2456 64932 2508
rect 67548 2592 67600 2644
rect 111064 3884 111116 3936
rect 112444 3816 112496 3868
rect 112536 3748 112588 3800
rect 68836 2592 68888 2644
rect 68928 2592 68980 2644
rect 69020 2592 69072 2644
rect 69848 2592 69900 2644
rect 70676 2592 70728 2644
rect 72424 2592 72476 2644
rect 72516 2592 72568 2644
rect 112628 3680 112680 3732
rect 112720 3612 112772 3664
rect 112812 3544 112864 3596
rect 75000 2592 75052 2644
rect 76288 2592 76340 2644
rect 76472 2592 76524 2644
rect 111156 3476 111208 3528
rect 111248 3408 111300 3460
rect 114192 3340 114244 3392
rect 114100 3272 114152 3324
rect 109592 3000 109644 3052
rect 117964 3000 118016 3052
rect 117688 2932 117740 2984
rect 84016 2592 84068 2644
rect 84476 2592 84528 2644
rect 84568 2592 84620 2644
rect 84752 2592 84804 2644
rect 85304 2592 85356 2644
rect 76564 2524 76616 2576
rect 85856 2592 85908 2644
rect 115848 2864 115900 2916
rect 98276 2592 98328 2644
rect 106096 2592 106148 2644
rect 72516 2456 72568 2508
rect 109592 2456 109644 2508
rect 116584 2456 116636 2508
rect 294788 2456 294840 2508
rect 425796 2456 425848 2508
rect 443644 2456 443696 2508
rect 59820 2320 59872 2372
rect 68836 2388 68888 2440
rect 84016 2388 84068 2440
rect 106188 2388 106240 2440
rect 116676 2388 116728 2440
rect 76564 2320 76616 2372
rect 102968 2320 103020 2372
rect 116768 2320 116820 2372
rect 42984 2252 43036 2304
rect 49884 2252 49936 2304
rect 52920 2252 52972 2304
rect 58992 2252 59044 2304
rect 68928 2252 68980 2304
rect 84476 2252 84528 2304
rect 99656 2252 99708 2304
rect 116860 2252 116912 2304
rect 69664 2184 69716 2236
rect 84752 2184 84804 2236
rect 96344 2184 96396 2236
rect 116952 2184 117004 2236
rect 63040 2116 63092 2168
rect 69848 2116 69900 2168
rect 76288 2116 76340 2168
rect 93032 2116 93084 2168
rect 117044 2116 117096 2168
rect 70676 2048 70728 2100
rect 75000 2048 75052 2100
rect 89628 2048 89680 2100
rect 117136 2048 117188 2100
rect 72424 1980 72476 2032
rect 86408 1980 86460 2032
rect 117228 1980 117280 2032
rect 82636 1912 82688 1964
rect 116492 1912 116544 1964
rect 79324 1844 79376 1896
rect 116400 1844 116452 1896
rect 72700 1776 72752 1828
rect 109684 1776 109736 1828
rect 76012 1708 76064 1760
rect 116308 1708 116360 1760
rect 32680 1640 32732 1692
rect 116216 1640 116268 1692
rect 29276 1572 29328 1624
rect 116032 1572 116084 1624
rect 25964 1504 26016 1556
rect 116124 1504 116176 1556
rect 22652 1436 22704 1488
rect 115940 1436 115992 1488
rect 117688 1436 117740 1488
rect 143632 1436 143684 1488
rect 6000 1368 6052 1420
rect 109776 1368 109828 1420
rect 117964 1368 118016 1420
rect 193588 1368 193640 1420
rect 294788 1368 294840 1420
rect 343640 1368 343692 1420
rect 491300 1368 491352 1420
rect 493600 1368 493652 1420
<< metal2 >>
rect 386 163200 442 164400
rect 492 163254 1164 163282
rect 400 158030 428 163200
rect 388 158024 440 158030
rect 388 157966 440 157972
rect 492 153882 520 163254
rect 1136 163146 1164 163254
rect 1214 163200 1270 164400
rect 2042 163200 2098 164400
rect 2870 163200 2926 164400
rect 2976 163254 3648 163282
rect 1228 163146 1256 163200
rect 1136 163118 1256 163146
rect 2056 156670 2084 163200
rect 2044 156664 2096 156670
rect 2044 156606 2096 156612
rect 480 153876 532 153882
rect 480 153818 532 153824
rect 2884 152522 2912 163200
rect 2976 153950 3004 163254
rect 3620 163146 3648 163254
rect 3698 163200 3754 164400
rect 4526 163200 4582 164400
rect 5354 163200 5410 164400
rect 6274 163200 6330 164400
rect 7102 163200 7158 164400
rect 7930 163200 7986 164400
rect 8758 163200 8814 164400
rect 8864 163254 9536 163282
rect 3712 163146 3740 163200
rect 3620 163118 3740 163146
rect 4540 155310 4568 163200
rect 4528 155304 4580 155310
rect 4528 155246 4580 155252
rect 5368 155242 5396 163200
rect 6288 159390 6316 163200
rect 6276 159384 6328 159390
rect 6276 159326 6328 159332
rect 5356 155236 5408 155242
rect 5356 155178 5408 155184
rect 7116 154018 7144 163200
rect 7944 155446 7972 163200
rect 7932 155440 7984 155446
rect 7932 155382 7984 155388
rect 8772 155378 8800 163200
rect 8760 155372 8812 155378
rect 8760 155314 8812 155320
rect 7104 154012 7156 154018
rect 7104 153954 7156 153960
rect 2964 153944 3016 153950
rect 2964 153886 3016 153892
rect 2872 152516 2924 152522
rect 2872 152458 2924 152464
rect 8864 152425 8892 163254
rect 9508 163146 9536 163254
rect 9586 163200 9642 164400
rect 9692 163254 10364 163282
rect 9600 163146 9628 163200
rect 9508 163118 9628 163146
rect 9692 154086 9720 163254
rect 10336 163146 10364 163254
rect 10414 163200 10470 164400
rect 11242 163200 11298 164400
rect 12162 163200 12218 164400
rect 12452 163254 12940 163282
rect 10428 163146 10456 163200
rect 10336 163118 10456 163146
rect 11256 156058 11284 163200
rect 11244 156052 11296 156058
rect 11244 155994 11296 156000
rect 12176 155854 12204 163200
rect 12164 155848 12216 155854
rect 12164 155790 12216 155796
rect 9680 154080 9732 154086
rect 9680 154022 9732 154028
rect 12452 152561 12480 163254
rect 12912 163146 12940 163254
rect 12990 163200 13046 164400
rect 13818 163200 13874 164400
rect 14646 163200 14702 164400
rect 15212 163254 15424 163282
rect 13004 163146 13032 163200
rect 12912 163118 13032 163146
rect 13832 154154 13860 163200
rect 14660 156738 14688 163200
rect 14648 156732 14700 156738
rect 14648 156674 14700 156680
rect 13820 154148 13872 154154
rect 13820 154090 13872 154096
rect 15212 152658 15240 163254
rect 15396 163146 15424 163254
rect 15474 163200 15530 164400
rect 16302 163200 16358 164400
rect 16592 163254 17080 163282
rect 15488 163146 15516 163200
rect 15396 163118 15516 163146
rect 16316 159497 16344 163200
rect 16302 159488 16358 159497
rect 16302 159423 16358 159432
rect 16592 153785 16620 163254
rect 17052 163146 17080 163254
rect 17130 163200 17186 164400
rect 18050 163200 18106 164400
rect 18878 163200 18934 164400
rect 19352 163254 19656 163282
rect 17144 163146 17172 163200
rect 17052 163118 17172 163146
rect 18064 156942 18092 163200
rect 18892 159730 18920 163200
rect 18880 159724 18932 159730
rect 18880 159666 18932 159672
rect 18052 156936 18104 156942
rect 18052 156878 18104 156884
rect 16578 153776 16634 153785
rect 16578 153711 16634 153720
rect 15200 152652 15252 152658
rect 15200 152594 15252 152600
rect 19352 152590 19380 163254
rect 19628 163146 19656 163254
rect 19706 163200 19762 164400
rect 19904 163254 20484 163282
rect 19720 163146 19748 163200
rect 19628 163118 19748 163146
rect 19904 153921 19932 163254
rect 20456 163146 20484 163254
rect 20534 163200 20590 164400
rect 21362 163200 21418 164400
rect 22190 163200 22246 164400
rect 23018 163200 23074 164400
rect 23492 163254 23888 163282
rect 20548 163146 20576 163200
rect 20456 163118 20576 163146
rect 21376 156874 21404 163200
rect 21364 156868 21416 156874
rect 21364 156810 21416 156816
rect 19890 153912 19946 153921
rect 19890 153847 19946 153856
rect 22204 152726 22232 163200
rect 23032 159361 23060 163200
rect 23018 159352 23074 159361
rect 23018 159287 23074 159296
rect 23492 154222 23520 163254
rect 23860 163146 23888 163254
rect 23938 163200 23994 164400
rect 24766 163200 24822 164400
rect 25594 163200 25650 164400
rect 26422 163200 26478 164400
rect 27250 163200 27306 164400
rect 28078 163200 28134 164400
rect 28906 163200 28962 164400
rect 29826 163200 29882 164400
rect 30392 163254 30604 163282
rect 23952 163146 23980 163200
rect 23860 163118 23980 163146
rect 24780 157010 24808 163200
rect 25608 160002 25636 163200
rect 25596 159996 25648 160002
rect 25596 159938 25648 159944
rect 24768 157004 24820 157010
rect 24768 156946 24820 156952
rect 23480 154216 23532 154222
rect 23480 154158 23532 154164
rect 26436 152794 26464 163200
rect 27264 154057 27292 163200
rect 28092 156641 28120 163200
rect 28078 156632 28134 156641
rect 28078 156567 28134 156576
rect 28920 155514 28948 163200
rect 29840 159633 29868 163200
rect 29826 159624 29882 159633
rect 29826 159559 29882 159568
rect 28908 155508 28960 155514
rect 28908 155450 28960 155456
rect 30392 154290 30420 163254
rect 30576 163146 30604 163254
rect 30654 163200 30710 164400
rect 31482 163200 31538 164400
rect 32310 163200 32366 164400
rect 33138 163200 33194 164400
rect 33966 163200 34022 164400
rect 34532 163254 34744 163282
rect 30668 163146 30696 163200
rect 30576 163118 30696 163146
rect 31496 156777 31524 163200
rect 32324 159594 32352 163200
rect 32312 159588 32364 159594
rect 32312 159530 32364 159536
rect 31482 156768 31538 156777
rect 31482 156703 31538 156712
rect 33152 155650 33180 163200
rect 33980 158001 34008 163200
rect 33966 157992 34022 158001
rect 33966 157927 34022 157936
rect 33140 155644 33192 155650
rect 33140 155586 33192 155592
rect 34532 154426 34560 163254
rect 34716 163146 34744 163254
rect 34794 163200 34850 164400
rect 35714 163200 35770 164400
rect 36542 163200 36598 164400
rect 37370 163200 37426 164400
rect 37936 163254 38148 163282
rect 34808 163146 34836 163200
rect 34716 163118 34836 163146
rect 35728 157078 35756 163200
rect 36556 159458 36584 163200
rect 36544 159452 36596 159458
rect 36544 159394 36596 159400
rect 37384 158098 37412 163200
rect 37372 158092 37424 158098
rect 37372 158034 37424 158040
rect 35716 157072 35768 157078
rect 35716 157014 35768 157020
rect 34520 154420 34572 154426
rect 34520 154362 34572 154368
rect 37936 154358 37964 163254
rect 38120 163146 38148 163254
rect 38198 163200 38254 164400
rect 39026 163200 39082 164400
rect 39854 163200 39910 164400
rect 40682 163200 40738 164400
rect 41602 163200 41658 164400
rect 42430 163200 42486 164400
rect 43258 163200 43314 164400
rect 44086 163200 44142 164400
rect 44192 163254 44864 163282
rect 38212 163146 38240 163200
rect 38120 163118 38240 163146
rect 39040 157146 39068 163200
rect 39028 157140 39080 157146
rect 39028 157082 39080 157088
rect 39868 155582 39896 163200
rect 40696 158137 40724 163200
rect 40682 158128 40738 158137
rect 40682 158063 40738 158072
rect 39856 155576 39908 155582
rect 39856 155518 39908 155524
rect 41616 154494 41644 163200
rect 42444 156913 42472 163200
rect 43272 159526 43300 163200
rect 43260 159520 43312 159526
rect 43260 159462 43312 159468
rect 44100 158273 44128 163200
rect 44086 158264 44142 158273
rect 44086 158199 44142 158208
rect 42430 156904 42486 156913
rect 42430 156839 42486 156848
rect 44192 154562 44220 163254
rect 44836 163146 44864 163254
rect 44914 163200 44970 164400
rect 45742 163200 45798 164400
rect 46570 163200 46626 164400
rect 47490 163200 47546 164400
rect 48318 163200 48374 164400
rect 49146 163200 49202 164400
rect 49974 163200 50030 164400
rect 50802 163200 50858 164400
rect 51092 163254 51580 163282
rect 44928 163146 44956 163200
rect 44836 163118 44956 163146
rect 45756 157214 45784 163200
rect 45744 157208 45796 157214
rect 45744 157150 45796 157156
rect 46584 155786 46612 163200
rect 47504 158166 47532 163200
rect 47492 158160 47544 158166
rect 47492 158102 47544 158108
rect 46572 155780 46624 155786
rect 46572 155722 46624 155728
rect 44180 154556 44232 154562
rect 44180 154498 44232 154504
rect 41604 154488 41656 154494
rect 41604 154430 41656 154436
rect 37924 154352 37976 154358
rect 37924 154294 37976 154300
rect 30380 154284 30432 154290
rect 30380 154226 30432 154232
rect 27250 154048 27306 154057
rect 27250 153983 27306 153992
rect 48332 153814 48360 163200
rect 49160 157049 49188 163200
rect 49988 159662 50016 163200
rect 49976 159656 50028 159662
rect 49976 159598 50028 159604
rect 50816 158234 50844 163200
rect 50804 158228 50856 158234
rect 50804 158170 50856 158176
rect 49146 157040 49202 157049
rect 49146 156975 49202 156984
rect 51092 154193 51120 163254
rect 51552 163146 51580 163254
rect 51630 163200 51686 164400
rect 52458 163200 52514 164400
rect 53378 163200 53434 164400
rect 54206 163200 54262 164400
rect 54312 163254 54984 163282
rect 51644 163146 51672 163200
rect 51552 163118 51672 163146
rect 52472 157350 52500 163200
rect 52460 157344 52512 157350
rect 52460 157286 52512 157292
rect 53392 155174 53420 163200
rect 54220 158302 54248 163200
rect 54208 158296 54260 158302
rect 54208 158238 54260 158244
rect 53380 155168 53432 155174
rect 53380 155110 53432 155116
rect 54312 154329 54340 163254
rect 54956 163146 54984 163254
rect 55034 163200 55090 164400
rect 55862 163200 55918 164400
rect 56690 163200 56746 164400
rect 57518 163200 57574 164400
rect 57992 163254 58296 163282
rect 55048 163146 55076 163200
rect 54956 163118 55076 163146
rect 55876 157282 55904 163200
rect 56704 159866 56732 163200
rect 56692 159860 56744 159866
rect 56692 159802 56744 159808
rect 57532 158409 57560 163200
rect 57518 158400 57574 158409
rect 57518 158335 57574 158344
rect 55864 157276 55916 157282
rect 55864 157218 55916 157224
rect 56508 155508 56560 155514
rect 56508 155450 56560 155456
rect 54298 154320 54354 154329
rect 54298 154255 54354 154264
rect 51078 154184 51134 154193
rect 51078 154119 51134 154128
rect 48320 153808 48372 153814
rect 48320 153750 48372 153756
rect 26424 152788 26476 152794
rect 26424 152730 26476 152736
rect 22192 152720 22244 152726
rect 22192 152662 22244 152668
rect 19340 152584 19392 152590
rect 12438 152552 12494 152561
rect 19340 152526 19392 152532
rect 12438 152487 12494 152496
rect 8850 152416 8906 152425
rect 8850 152351 8906 152360
rect 56520 152318 56548 155450
rect 57992 153746 58020 163254
rect 58268 163146 58296 163254
rect 58346 163200 58402 164400
rect 59266 163200 59322 164400
rect 60094 163200 60150 164400
rect 60922 163200 60978 164400
rect 61750 163200 61806 164400
rect 62578 163200 62634 164400
rect 63406 163200 63462 164400
rect 64234 163200 64290 164400
rect 64892 163254 65104 163282
rect 58360 163146 58388 163200
rect 58268 163118 58388 163146
rect 59280 156602 59308 163200
rect 59268 156596 59320 156602
rect 59268 156538 59320 156544
rect 60108 155922 60136 163200
rect 60936 158370 60964 163200
rect 60924 158364 60976 158370
rect 60924 158306 60976 158312
rect 60096 155916 60148 155922
rect 60096 155858 60148 155864
rect 60004 155644 60056 155650
rect 60004 155586 60056 155592
rect 57980 153740 58032 153746
rect 57980 153682 58032 153688
rect 60016 152454 60044 155586
rect 61764 155281 61792 163200
rect 62592 155514 62620 163200
rect 63420 159798 63448 163200
rect 63408 159792 63460 159798
rect 63408 159734 63460 159740
rect 64248 158438 64276 163200
rect 64236 158432 64288 158438
rect 64236 158374 64288 158380
rect 62580 155508 62632 155514
rect 62580 155450 62632 155456
rect 61750 155272 61806 155281
rect 61750 155207 61806 155216
rect 64892 153678 64920 163254
rect 65076 163146 65104 163254
rect 65154 163200 65210 164400
rect 65982 163200 66038 164400
rect 66272 163254 66760 163282
rect 65168 163146 65196 163200
rect 65076 163118 65196 163146
rect 65996 157185 66024 163200
rect 65982 157176 66038 157185
rect 65982 157111 66038 157120
rect 64880 153672 64932 153678
rect 64880 153614 64932 153620
rect 66272 152862 66300 163254
rect 66732 163146 66760 163254
rect 66810 163200 66866 164400
rect 67638 163200 67694 164400
rect 68466 163200 68522 164400
rect 69294 163200 69350 164400
rect 70122 163200 70178 164400
rect 71042 163200 71098 164400
rect 71870 163200 71926 164400
rect 72698 163200 72754 164400
rect 73526 163200 73582 164400
rect 74354 163200 74410 164400
rect 75182 163200 75238 164400
rect 76010 163200 76066 164400
rect 76930 163200 76986 164400
rect 77758 163200 77814 164400
rect 78586 163200 78642 164400
rect 79414 163200 79470 164400
rect 80242 163200 80298 164400
rect 81070 163200 81126 164400
rect 81898 163200 81954 164400
rect 82818 163200 82874 164400
rect 83646 163200 83702 164400
rect 84474 163200 84530 164400
rect 85302 163200 85358 164400
rect 86130 163200 86186 164400
rect 86958 163200 87014 164400
rect 87786 163200 87842 164400
rect 88706 163200 88762 164400
rect 89534 163200 89590 164400
rect 89824 163254 90312 163282
rect 66824 163146 66852 163200
rect 66732 163118 66852 163146
rect 67652 158642 67680 163200
rect 67640 158636 67692 158642
rect 67640 158578 67692 158584
rect 68480 155417 68508 163200
rect 69308 155553 69336 163200
rect 70136 159934 70164 163200
rect 70124 159928 70176 159934
rect 70124 159870 70176 159876
rect 71056 158506 71084 163200
rect 71044 158500 71096 158506
rect 71044 158442 71096 158448
rect 71884 155718 71912 163200
rect 72712 156534 72740 163200
rect 73540 158982 73568 163200
rect 73528 158976 73580 158982
rect 73528 158918 73580 158924
rect 74368 158574 74396 163200
rect 74356 158568 74408 158574
rect 74356 158510 74408 158516
rect 72700 156528 72752 156534
rect 72700 156470 72752 156476
rect 71872 155712 71924 155718
rect 71872 155654 71924 155660
rect 75196 155650 75224 163200
rect 75828 155780 75880 155786
rect 75828 155722 75880 155728
rect 75184 155644 75236 155650
rect 75184 155586 75236 155592
rect 71780 155576 71832 155582
rect 69294 155544 69350 155553
rect 71780 155518 71832 155524
rect 69294 155479 69350 155488
rect 68466 155408 68522 155417
rect 68466 155343 68522 155352
rect 66260 152856 66312 152862
rect 66260 152798 66312 152804
rect 60004 152448 60056 152454
rect 60004 152390 60056 152396
rect 56508 152312 56560 152318
rect 56508 152254 56560 152260
rect 71792 152046 71820 155518
rect 75840 152114 75868 155722
rect 76024 155689 76052 163200
rect 76944 159322 76972 163200
rect 76932 159316 76984 159322
rect 76932 159258 76984 159264
rect 77772 157962 77800 163200
rect 77760 157956 77812 157962
rect 77760 157898 77812 157904
rect 76010 155680 76066 155689
rect 76010 155615 76066 155624
rect 78600 155582 78628 163200
rect 79428 156466 79456 163200
rect 79416 156460 79468 156466
rect 79416 156402 79468 156408
rect 78588 155576 78640 155582
rect 78588 155518 78640 155524
rect 76932 155168 76984 155174
rect 76932 155110 76984 155116
rect 76944 152250 76972 155110
rect 80256 154902 80284 163200
rect 81084 158710 81112 163200
rect 81072 158704 81124 158710
rect 81072 158646 81124 158652
rect 81912 155786 81940 163200
rect 81900 155780 81952 155786
rect 81900 155722 81952 155728
rect 80244 154896 80296 154902
rect 80244 154838 80296 154844
rect 82832 153610 82860 163200
rect 83660 160070 83688 163200
rect 83648 160064 83700 160070
rect 83648 160006 83700 160012
rect 84488 157894 84516 163200
rect 84476 157888 84528 157894
rect 84476 157830 84528 157836
rect 84752 155916 84804 155922
rect 84752 155858 84804 155864
rect 82820 153604 82872 153610
rect 82820 153546 82872 153552
rect 76932 152244 76984 152250
rect 76932 152186 76984 152192
rect 84764 152182 84792 155858
rect 85316 155825 85344 163200
rect 85302 155816 85358 155825
rect 85302 155751 85358 155760
rect 86144 155174 86172 163200
rect 86972 159186 87000 163200
rect 86960 159180 87012 159186
rect 86960 159122 87012 159128
rect 87800 157826 87828 163200
rect 87788 157820 87840 157826
rect 87788 157762 87840 157768
rect 88720 155922 88748 163200
rect 89548 158794 89576 163200
rect 89548 158766 89760 158794
rect 88708 155916 88760 155922
rect 88708 155858 88760 155864
rect 86132 155168 86184 155174
rect 86132 155110 86184 155116
rect 86868 154896 86920 154902
rect 86868 154838 86920 154844
rect 86880 153134 86908 154838
rect 89732 154465 89760 158766
rect 89718 154456 89774 154465
rect 89718 154391 89774 154400
rect 86868 153128 86920 153134
rect 86868 153070 86920 153076
rect 89824 152930 89852 163254
rect 90284 163146 90312 163254
rect 90362 163200 90418 164400
rect 91190 163200 91246 164400
rect 92018 163200 92074 164400
rect 92846 163200 92902 164400
rect 93674 163200 93730 164400
rect 94594 163200 94650 164400
rect 95422 163200 95478 164400
rect 96250 163200 96306 164400
rect 96632 163254 97028 163282
rect 90376 163146 90404 163200
rect 90284 163118 90404 163146
rect 91204 157758 91232 163200
rect 91192 157752 91244 157758
rect 91192 157694 91244 157700
rect 92032 155961 92060 163200
rect 92860 156398 92888 163200
rect 93688 159254 93716 163200
rect 93676 159248 93728 159254
rect 93676 159190 93728 159196
rect 94608 157690 94636 163200
rect 94596 157684 94648 157690
rect 94596 157626 94648 157632
rect 92848 156392 92900 156398
rect 92848 156334 92900 156340
rect 92018 155952 92074 155961
rect 92018 155887 92074 155896
rect 95436 155106 95464 163200
rect 96264 158914 96292 163200
rect 96252 158908 96304 158914
rect 96252 158850 96304 158856
rect 95424 155100 95476 155106
rect 95424 155042 95476 155048
rect 96632 152998 96660 163254
rect 97000 163146 97028 163254
rect 97078 163200 97134 164400
rect 97906 163200 97962 164400
rect 98734 163200 98790 164400
rect 99562 163200 99618 164400
rect 100482 163200 100538 164400
rect 101310 163200 101366 164400
rect 102138 163200 102194 164400
rect 102966 163200 103022 164400
rect 103532 163254 103744 163282
rect 97092 163146 97120 163200
rect 97000 163118 97120 163146
rect 97920 157622 97948 163200
rect 97908 157616 97960 157622
rect 97908 157558 97960 157564
rect 98748 155038 98776 163200
rect 98736 155032 98788 155038
rect 98736 154974 98788 154980
rect 99576 154970 99604 163200
rect 100496 159118 100524 163200
rect 100484 159112 100536 159118
rect 100484 159054 100536 159060
rect 101324 156330 101352 163200
rect 101312 156324 101364 156330
rect 101312 156266 101364 156272
rect 99564 154964 99616 154970
rect 99564 154906 99616 154912
rect 102152 153542 102180 163200
rect 102980 158846 103008 163200
rect 102968 158840 103020 158846
rect 102968 158782 103020 158788
rect 102140 153536 102192 153542
rect 102140 153478 102192 153484
rect 103532 153066 103560 163254
rect 103716 163146 103744 163254
rect 103794 163200 103850 164400
rect 104622 163200 104678 164400
rect 104912 163254 105400 163282
rect 103808 163146 103836 163200
rect 103716 163118 103836 163146
rect 104636 158545 104664 163200
rect 104622 158536 104678 158545
rect 104622 158471 104678 158480
rect 104912 153474 104940 163254
rect 105372 163146 105400 163254
rect 105450 163200 105506 164400
rect 106370 163200 106426 164400
rect 107198 163200 107254 164400
rect 108026 163200 108082 164400
rect 108316 163254 108804 163282
rect 105464 163146 105492 163200
rect 105372 163118 105492 163146
rect 106384 158778 106412 163200
rect 107212 159050 107240 163200
rect 107292 159724 107344 159730
rect 107292 159666 107344 159672
rect 107200 159044 107252 159050
rect 107200 158986 107252 158992
rect 106372 158772 106424 158778
rect 106372 158714 106424 158720
rect 107304 154766 107332 159666
rect 107568 158976 107620 158982
rect 107568 158918 107620 158924
rect 107292 154760 107344 154766
rect 107292 154702 107344 154708
rect 104900 153468 104952 153474
rect 104900 153410 104952 153416
rect 103520 153060 103572 153066
rect 103520 153002 103572 153008
rect 96620 152992 96672 152998
rect 96620 152934 96672 152940
rect 89812 152924 89864 152930
rect 89812 152866 89864 152872
rect 84752 152176 84804 152182
rect 84752 152118 84804 152124
rect 75828 152108 75880 152114
rect 75828 152050 75880 152056
rect 71780 152040 71832 152046
rect 71780 151982 71832 151988
rect 107580 151910 107608 158918
rect 108040 156262 108068 163200
rect 108028 156256 108080 156262
rect 108028 156198 108080 156204
rect 108316 153406 108344 163254
rect 108776 163146 108804 163254
rect 108854 163200 108910 164400
rect 109682 163200 109738 164400
rect 110510 163200 110566 164400
rect 111338 163200 111394 164400
rect 112258 163200 112314 164400
rect 113086 163200 113142 164400
rect 113192 163254 113864 163282
rect 108868 163146 108896 163200
rect 108776 163118 108896 163146
rect 109696 159730 109724 163200
rect 109868 159996 109920 160002
rect 109868 159938 109920 159944
rect 109684 159724 109736 159730
rect 109684 159666 109736 159672
rect 109040 155848 109092 155854
rect 109040 155790 109092 155796
rect 108304 153400 108356 153406
rect 108304 153342 108356 153348
rect 109052 151978 109080 155790
rect 109040 151972 109092 151978
rect 109040 151914 109092 151920
rect 30196 151904 30248 151910
rect 30196 151846 30248 151852
rect 74540 151904 74592 151910
rect 74540 151846 74592 151852
rect 107568 151904 107620 151910
rect 107568 151846 107620 151852
rect 19800 150612 19852 150618
rect 19800 150554 19852 150560
rect 16396 150544 16448 150550
rect 16396 150486 16448 150492
rect 2688 150476 2740 150482
rect 2688 150418 2740 150424
rect 2700 149940 2728 150418
rect 6368 150068 6420 150074
rect 6368 150010 6420 150016
rect 6380 149954 6408 150010
rect 6118 149926 6408 149954
rect 13018 149938 13400 149954
rect 16408 149940 16436 150486
rect 19812 149940 19840 150554
rect 23388 150000 23440 150006
rect 23322 149948 23388 149954
rect 23322 149942 23440 149948
rect 13018 149932 13412 149938
rect 13018 149926 13360 149932
rect 23322 149926 23428 149942
rect 30208 149940 30236 151846
rect 33600 151836 33652 151842
rect 33600 151778 33652 151784
rect 33612 149940 33640 151778
rect 74552 151366 74580 151846
rect 109880 151842 109908 159938
rect 110524 154698 110552 163200
rect 111352 157554 111380 163200
rect 111340 157548 111392 157554
rect 111340 157490 111392 157496
rect 112272 155854 112300 163200
rect 113100 157321 113128 163200
rect 113086 157312 113142 157321
rect 113086 157247 113142 157256
rect 112260 155848 112312 155854
rect 112260 155790 112312 155796
rect 110512 154692 110564 154698
rect 110512 154634 110564 154640
rect 113192 152386 113220 163254
rect 113836 163146 113864 163254
rect 113914 163200 113970 164400
rect 114742 163200 114798 164400
rect 114848 163254 115520 163282
rect 113928 163146 113956 163200
rect 113836 163118 113956 163146
rect 114756 157486 114784 163200
rect 114744 157480 114796 157486
rect 114744 157422 114796 157428
rect 114848 153338 114876 163254
rect 115492 163146 115520 163254
rect 115570 163200 115626 164400
rect 115952 163254 116348 163282
rect 115584 163146 115612 163200
rect 115492 163118 115612 163146
rect 114836 153332 114888 153338
rect 114836 153274 114888 153280
rect 115952 153270 115980 163254
rect 116320 163146 116348 163254
rect 116398 163200 116454 164400
rect 117226 163200 117282 164400
rect 118146 163200 118202 164400
rect 118974 163200 119030 164400
rect 119802 163200 119858 164400
rect 120184 163254 120580 163282
rect 116412 163146 116440 163200
rect 116320 163118 116440 163146
rect 117240 160002 117268 163200
rect 117228 159996 117280 160002
rect 117228 159938 117280 159944
rect 118160 156194 118188 163200
rect 118988 161474 119016 163200
rect 118804 161446 119016 161474
rect 118148 156188 118200 156194
rect 118148 156130 118200 156136
rect 117964 154012 118016 154018
rect 117964 153954 118016 153960
rect 117976 153898 118004 153954
rect 118148 153944 118200 153950
rect 117976 153892 118148 153898
rect 117976 153886 118200 153892
rect 117976 153870 118188 153886
rect 118606 153368 118662 153377
rect 118804 153338 118832 161446
rect 119816 158982 119844 163200
rect 119804 158976 119856 158982
rect 119804 158918 119856 158924
rect 118884 158024 118936 158030
rect 118884 157966 118936 157972
rect 118606 153303 118608 153312
rect 118660 153303 118662 153312
rect 118792 153332 118844 153338
rect 118608 153274 118660 153280
rect 118792 153274 118844 153280
rect 115940 153264 115992 153270
rect 115940 153206 115992 153212
rect 113180 152380 113232 152386
rect 113180 152322 113232 152328
rect 84200 151836 84252 151842
rect 84200 151778 84252 151784
rect 105820 151836 105872 151842
rect 105820 151778 105872 151784
rect 109776 151836 109828 151842
rect 109776 151778 109828 151784
rect 109868 151836 109920 151842
rect 109868 151778 109920 151784
rect 84212 151434 84240 151778
rect 84200 151428 84252 151434
rect 84200 151370 84252 151376
rect 74540 151360 74592 151366
rect 74540 151302 74592 151308
rect 68008 151292 68060 151298
rect 68008 151234 68060 151240
rect 64512 151224 64564 151230
rect 64512 151166 64564 151172
rect 61108 151156 61160 151162
rect 61108 151098 61160 151104
rect 57704 151088 57756 151094
rect 57704 151030 57756 151036
rect 54208 151020 54260 151026
rect 54208 150962 54260 150968
rect 50804 150952 50856 150958
rect 50804 150894 50856 150900
rect 47308 150884 47360 150890
rect 47308 150826 47360 150832
rect 43904 150816 43956 150822
rect 43904 150758 43956 150764
rect 40500 150748 40552 150754
rect 40500 150690 40552 150696
rect 37004 150680 37056 150686
rect 37004 150622 37056 150628
rect 37016 149940 37044 150622
rect 40512 149940 40540 150690
rect 43916 149940 43944 150758
rect 47320 149940 47348 150826
rect 50816 149940 50844 150894
rect 54220 149940 54248 150962
rect 57716 149940 57744 151030
rect 61120 149940 61148 151098
rect 64524 149940 64552 151166
rect 68020 149940 68048 151234
rect 105832 149940 105860 151778
rect 13360 149874 13412 149880
rect 9588 149864 9640 149870
rect 9522 149812 9588 149818
rect 9522 149806 9640 149812
rect 9522 149790 9628 149806
rect 88642 149802 89024 149818
rect 88642 149796 89036 149802
rect 88642 149790 88984 149796
rect 88984 149738 89036 149744
rect 85488 149728 85540 149734
rect 81742 149666 82032 149682
rect 85238 149676 85488 149682
rect 85238 149670 85540 149676
rect 81742 149660 82044 149666
rect 81742 149654 81992 149660
rect 85238 149654 85528 149670
rect 81992 149602 82044 149608
rect 78588 149592 78640 149598
rect 74842 149530 75224 149546
rect 78338 149540 78588 149546
rect 102598 149560 102654 149569
rect 78338 149534 78640 149540
rect 74842 149524 75236 149530
rect 74842 149518 75184 149524
rect 78338 149518 78628 149534
rect 102350 149518 102598 149546
rect 102598 149495 102654 149504
rect 109682 149560 109738 149569
rect 109682 149495 109738 149504
rect 75184 149466 75236 149472
rect 71688 149456 71740 149462
rect 26726 149394 27016 149410
rect 71438 149404 71688 149410
rect 99286 149424 99342 149433
rect 71438 149398 71740 149404
rect 26726 149388 27028 149394
rect 26726 149382 26976 149388
rect 71438 149382 71728 149398
rect 92046 149382 92336 149410
rect 95542 149382 95832 149410
rect 98946 149382 99286 149410
rect 26976 149330 27028 149336
rect 92308 149326 92336 149382
rect 95804 149326 95832 149382
rect 99286 149359 99342 149368
rect 105266 149424 105322 149433
rect 109250 149382 109632 149410
rect 105266 149359 105322 149368
rect 105280 149326 105308 149359
rect 92296 149320 92348 149326
rect 92296 149262 92348 149268
rect 95792 149320 95844 149326
rect 95792 149262 95844 149268
rect 105268 149320 105320 149326
rect 105268 149262 105320 149268
rect 109604 149054 109632 149382
rect 109696 149190 109724 149495
rect 109684 149184 109736 149190
rect 109684 149126 109736 149132
rect 109592 149048 109644 149054
rect 109592 148990 109644 148996
rect 109788 147626 109816 151778
rect 117228 151428 117280 151434
rect 117228 151370 117280 151376
rect 117136 151360 117188 151366
rect 117136 151302 117188 151308
rect 112812 151292 112864 151298
rect 112812 151234 112864 151240
rect 112720 151224 112772 151230
rect 112720 151166 112772 151172
rect 112628 151156 112680 151162
rect 112628 151098 112680 151104
rect 112536 151088 112588 151094
rect 112536 151030 112588 151036
rect 111616 151020 111668 151026
rect 111616 150962 111668 150968
rect 111524 150884 111576 150890
rect 111524 150826 111576 150832
rect 111432 150816 111484 150822
rect 111432 150758 111484 150764
rect 111340 150748 111392 150754
rect 111340 150690 111392 150696
rect 111248 150680 111300 150686
rect 111248 150622 111300 150628
rect 111064 150476 111116 150482
rect 111064 150418 111116 150424
rect 109776 147620 109828 147626
rect 109776 147562 109828 147568
rect 111076 89690 111104 150418
rect 111156 150068 111208 150074
rect 111156 150010 111208 150016
rect 111168 92478 111196 150010
rect 111260 109002 111288 150622
rect 111352 111790 111380 150690
rect 111444 113150 111472 150758
rect 111536 114510 111564 150826
rect 111628 118658 111656 150962
rect 112444 150952 112496 150958
rect 112444 150894 112496 150900
rect 112352 149660 112404 149666
rect 112352 149602 112404 149608
rect 112364 133890 112392 149602
rect 112352 133884 112404 133890
rect 112352 133826 112404 133832
rect 111616 118652 111668 118658
rect 111616 118594 111668 118600
rect 112456 117298 112484 150894
rect 112548 121446 112576 151030
rect 112640 122806 112668 151098
rect 112732 124166 112760 151166
rect 112824 126954 112852 151234
rect 116860 150612 116912 150618
rect 116860 150554 116912 150560
rect 116768 150544 116820 150550
rect 116768 150486 116820 150492
rect 116676 149932 116728 149938
rect 116676 149874 116728 149880
rect 116584 149864 116636 149870
rect 116584 149806 116636 149812
rect 114008 149796 114060 149802
rect 114008 149738 114060 149744
rect 113916 149728 113968 149734
rect 113916 149670 113968 149676
rect 113088 149592 113140 149598
rect 113088 149534 113140 149540
rect 112996 149524 113048 149530
rect 112996 149466 113048 149472
rect 112904 149456 112956 149462
rect 112904 149398 112956 149404
rect 112916 128314 112944 149398
rect 113008 131102 113036 149466
rect 113100 132462 113128 149534
rect 113822 143712 113878 143721
rect 113822 143647 113878 143656
rect 113088 132456 113140 132462
rect 113088 132398 113140 132404
rect 112996 131096 113048 131102
rect 112996 131038 113048 131044
rect 112904 128308 112956 128314
rect 112904 128250 112956 128256
rect 112812 126948 112864 126954
rect 112812 126890 112864 126896
rect 112720 124160 112772 124166
rect 112720 124102 112772 124108
rect 112628 122800 112680 122806
rect 112628 122742 112680 122748
rect 112536 121440 112588 121446
rect 112536 121382 112588 121388
rect 112444 117292 112496 117298
rect 112444 117234 112496 117240
rect 111524 114504 111576 114510
rect 111524 114446 111576 114452
rect 111432 113144 111484 113150
rect 111432 113086 111484 113092
rect 111340 111784 111392 111790
rect 111340 111726 111392 111732
rect 111248 108996 111300 109002
rect 111248 108938 111300 108944
rect 111156 92472 111208 92478
rect 111156 92414 111208 92420
rect 111064 89684 111116 89690
rect 111064 89626 111116 89632
rect 113836 88330 113864 143647
rect 113928 136610 113956 149670
rect 114020 137970 114048 149738
rect 116216 149320 116268 149326
rect 116216 149262 116268 149268
rect 116032 149184 116084 149190
rect 116032 149126 116084 149132
rect 114100 149116 114152 149122
rect 114100 149058 114152 149064
rect 114112 140758 114140 149058
rect 116044 145761 116072 149126
rect 116124 149048 116176 149054
rect 116124 148990 116176 148996
rect 116136 148753 116164 148990
rect 116122 148744 116178 148753
rect 116122 148679 116178 148688
rect 116124 147620 116176 147626
rect 116124 147562 116176 147568
rect 116136 147393 116164 147562
rect 116122 147384 116178 147393
rect 116122 147319 116178 147328
rect 116030 145752 116086 145761
rect 116030 145687 116086 145696
rect 116228 143449 116256 149262
rect 116492 149252 116544 149258
rect 116492 149194 116544 149200
rect 116214 143440 116270 143449
rect 116214 143375 116270 143384
rect 116504 141817 116532 149194
rect 116490 141808 116546 141817
rect 116490 141743 116546 141752
rect 114100 140752 114152 140758
rect 114100 140694 114152 140700
rect 116400 140752 116452 140758
rect 116400 140694 116452 140700
rect 116412 140049 116440 140694
rect 116398 140040 116454 140049
rect 116398 139975 116454 139984
rect 114008 137964 114060 137970
rect 114008 137906 114060 137912
rect 116216 137964 116268 137970
rect 116216 137906 116268 137912
rect 116228 137873 116256 137906
rect 116214 137864 116270 137873
rect 116214 137799 116270 137808
rect 113916 136604 113968 136610
rect 113916 136546 113968 136552
rect 116400 136604 116452 136610
rect 116400 136546 116452 136552
rect 116412 136105 116440 136546
rect 116398 136096 116454 136105
rect 116398 136031 116454 136040
rect 116124 133884 116176 133890
rect 116124 133826 116176 133832
rect 116136 133793 116164 133826
rect 116122 133784 116178 133793
rect 116122 133719 116178 133728
rect 113914 132560 113970 132569
rect 113914 132495 113970 132504
rect 113824 88324 113876 88330
rect 113824 88266 113876 88272
rect 113928 86970 113956 132495
rect 116124 132456 116176 132462
rect 116124 132398 116176 132404
rect 116136 132297 116164 132398
rect 116122 132288 116178 132297
rect 116122 132223 116178 132232
rect 116124 131096 116176 131102
rect 116124 131038 116176 131044
rect 116136 130393 116164 131038
rect 116122 130384 116178 130393
rect 116122 130319 116178 130328
rect 116124 128308 116176 128314
rect 116124 128250 116176 128256
rect 116136 128081 116164 128250
rect 116122 128072 116178 128081
rect 116122 128007 116178 128016
rect 116124 126948 116176 126954
rect 116124 126890 116176 126896
rect 116136 126449 116164 126890
rect 116122 126440 116178 126449
rect 116122 126375 116178 126384
rect 116124 124160 116176 124166
rect 116124 124102 116176 124108
rect 116136 123865 116164 124102
rect 116122 123856 116178 123865
rect 116122 123791 116178 123800
rect 116124 122800 116176 122806
rect 116124 122742 116176 122748
rect 116136 122641 116164 122742
rect 116122 122632 116178 122641
rect 116122 122567 116178 122576
rect 116124 121440 116176 121446
rect 116124 121382 116176 121388
rect 114006 120864 114062 120873
rect 114006 120799 114062 120808
rect 113916 86964 113968 86970
rect 113916 86906 113968 86912
rect 114020 83978 114048 120799
rect 116136 120737 116164 121382
rect 116122 120728 116178 120737
rect 116122 120663 116178 120672
rect 116124 118652 116176 118658
rect 116124 118594 116176 118600
rect 116136 118425 116164 118594
rect 116122 118416 116178 118425
rect 116122 118351 116178 118360
rect 116124 117292 116176 117298
rect 116124 117234 116176 117240
rect 116136 116793 116164 117234
rect 116122 116784 116178 116793
rect 116122 116719 116178 116728
rect 116124 114504 116176 114510
rect 116124 114446 116176 114452
rect 116136 114209 116164 114446
rect 116122 114200 116178 114209
rect 116122 114135 116178 114144
rect 116124 113144 116176 113150
rect 116124 113086 116176 113092
rect 116136 112985 116164 113086
rect 116122 112976 116178 112985
rect 116122 112911 116178 112920
rect 116124 111784 116176 111790
rect 116124 111726 116176 111732
rect 116136 111217 116164 111726
rect 116122 111208 116178 111217
rect 116122 111143 116178 111152
rect 114098 109576 114154 109585
rect 114098 109511 114154 109520
rect 114008 83972 114060 83978
rect 114008 83914 114060 83920
rect 114112 82822 114140 109511
rect 116124 108996 116176 109002
rect 116124 108938 116176 108944
rect 116136 108905 116164 108938
rect 116122 108896 116178 108905
rect 116122 108831 116178 108840
rect 114190 98152 114246 98161
rect 114190 98087 114246 98096
rect 114100 82816 114152 82822
rect 114100 82758 114152 82764
rect 114204 80034 114232 98087
rect 116596 93673 116624 149806
rect 116688 95849 116716 149874
rect 116780 97753 116808 150486
rect 116872 99385 116900 150554
rect 116952 150000 117004 150006
rect 116952 149942 117004 149948
rect 116964 101561 116992 149942
rect 117044 149388 117096 149394
rect 117044 149330 117096 149336
rect 117056 103193 117084 149330
rect 117148 104553 117176 151302
rect 117240 113234 117268 151370
rect 118896 149954 118924 157966
rect 119804 153876 119856 153882
rect 119804 153818 119856 153824
rect 119896 153876 119948 153882
rect 119896 153818 119948 153824
rect 119816 150226 119844 153818
rect 119908 153338 119936 153818
rect 119986 153368 120042 153377
rect 119896 153332 119948 153338
rect 119986 153303 119988 153312
rect 119896 153274 119948 153280
rect 120040 153303 120042 153312
rect 119988 153274 120040 153280
rect 120080 153196 120132 153202
rect 120080 153138 120132 153144
rect 120092 152386 120120 153138
rect 120184 152386 120212 163254
rect 120552 163146 120580 163254
rect 120630 163200 120686 164400
rect 121458 163200 121514 164400
rect 122286 163200 122342 164400
rect 123114 163200 123170 164400
rect 124034 163200 124090 164400
rect 124862 163200 124918 164400
rect 125690 163200 125746 164400
rect 126518 163200 126574 164400
rect 127346 163200 127402 164400
rect 128174 163200 128230 164400
rect 129002 163200 129058 164400
rect 129922 163200 129978 164400
rect 130750 163200 130806 164400
rect 131578 163200 131634 164400
rect 132406 163200 132462 164400
rect 133234 163200 133290 164400
rect 134062 163200 134118 164400
rect 134890 163200 134946 164400
rect 135810 163200 135866 164400
rect 136638 163200 136694 164400
rect 137466 163200 137522 164400
rect 138294 163200 138350 164400
rect 139122 163200 139178 164400
rect 139950 163200 140006 164400
rect 140778 163200 140834 164400
rect 141698 163200 141754 164400
rect 142526 163200 142582 164400
rect 143354 163200 143410 164400
rect 144182 163200 144238 164400
rect 145010 163200 145066 164400
rect 145838 163200 145894 164400
rect 146666 163200 146722 164400
rect 147586 163200 147642 164400
rect 148414 163200 148470 164400
rect 149242 163200 149298 164400
rect 150070 163200 150126 164400
rect 150898 163200 150954 164400
rect 151726 163200 151782 164400
rect 151832 163254 152504 163282
rect 120644 163146 120672 163200
rect 120552 163118 120672 163146
rect 120448 156664 120500 156670
rect 120448 156606 120500 156612
rect 120080 152380 120132 152386
rect 120080 152322 120132 152328
rect 120172 152380 120224 152386
rect 120172 152322 120224 152328
rect 120460 150226 120488 156606
rect 121472 156126 121500 163200
rect 121828 158908 121880 158914
rect 121828 158850 121880 158856
rect 121460 156120 121512 156126
rect 121460 156062 121512 156068
rect 121840 154018 121868 158850
rect 122012 155304 122064 155310
rect 122012 155246 122064 155252
rect 121736 154012 121788 154018
rect 121736 153954 121788 153960
rect 121828 154012 121880 154018
rect 121828 153954 121880 153960
rect 121092 152516 121144 152522
rect 121092 152458 121144 152464
rect 121104 150226 121132 152458
rect 121748 150226 121776 153954
rect 122024 151814 122052 155246
rect 122300 154902 122328 163200
rect 123128 159390 123156 163200
rect 122840 159384 122892 159390
rect 122840 159326 122892 159332
rect 123116 159384 123168 159390
rect 123116 159326 123168 159332
rect 122288 154896 122340 154902
rect 122288 154838 122340 154844
rect 122024 151786 122420 151814
rect 122392 150226 122420 151786
rect 119816 150198 119890 150226
rect 120460 150198 120534 150226
rect 121104 150198 121178 150226
rect 121748 150198 121822 150226
rect 122392 150198 122466 150226
rect 122852 150210 122880 159326
rect 124048 158914 124076 163200
rect 124036 158908 124088 158914
rect 124036 158850 124088 158856
rect 124876 156670 124904 163200
rect 125704 161474 125732 163200
rect 125704 161446 125824 161474
rect 125508 158840 125560 158846
rect 125508 158782 125560 158788
rect 124864 156664 124916 156670
rect 124864 156606 124916 156612
rect 124680 155440 124732 155446
rect 124680 155382 124732 155388
rect 123024 155236 123076 155242
rect 123024 155178 123076 155184
rect 123036 150226 123064 155178
rect 124312 153944 124364 153950
rect 124312 153886 124364 153892
rect 124324 150226 124352 153886
rect 124692 151814 124720 155382
rect 125520 153950 125548 158782
rect 125692 155372 125744 155378
rect 125692 155314 125744 155320
rect 125508 153944 125560 153950
rect 125508 153886 125560 153892
rect 124692 151786 124996 151814
rect 124968 150226 124996 151786
rect 125704 150226 125732 155314
rect 125796 154834 125824 161446
rect 126244 159588 126296 159594
rect 126244 159530 126296 159536
rect 125784 154828 125836 154834
rect 125784 154770 125836 154776
rect 126256 152697 126284 159530
rect 126532 158846 126560 163200
rect 126520 158840 126572 158846
rect 126520 158782 126572 158788
rect 127360 158778 127388 163200
rect 127624 159588 127676 159594
rect 127624 159530 127676 159536
rect 127636 158982 127664 159530
rect 127806 159488 127862 159497
rect 127806 159423 127862 159432
rect 127624 158976 127676 158982
rect 127624 158918 127676 158924
rect 127256 158772 127308 158778
rect 127256 158714 127308 158720
rect 127348 158772 127400 158778
rect 127348 158714 127400 158720
rect 127268 158030 127296 158714
rect 127256 158024 127308 158030
rect 127256 157966 127308 157972
rect 127532 156052 127584 156058
rect 127532 155994 127584 156000
rect 126808 154154 127020 154170
rect 126796 154148 127020 154154
rect 126848 154142 127020 154148
rect 126796 154090 126848 154096
rect 126888 154080 126940 154086
rect 126888 154022 126940 154028
rect 126992 154034 127020 154142
rect 126242 152688 126298 152697
rect 126242 152623 126298 152632
rect 126242 152416 126298 152425
rect 126242 152351 126298 152360
rect 118896 149926 119324 149954
rect 119862 149940 119890 150198
rect 120506 149940 120534 150198
rect 121150 149940 121178 150198
rect 121794 149940 121822 150198
rect 122438 149940 122466 150198
rect 122840 150204 122892 150210
rect 123036 150198 123110 150226
rect 122840 150146 122892 150152
rect 123082 149940 123110 150198
rect 123714 150204 123766 150210
rect 124324 150198 124398 150226
rect 124968 150198 125042 150226
rect 123714 150146 123766 150152
rect 123726 149940 123754 150146
rect 124370 149940 124398 150198
rect 125014 149940 125042 150198
rect 125658 150198 125732 150226
rect 126256 150226 126284 152351
rect 126900 150226 126928 154022
rect 126992 154006 127204 154034
rect 127176 153950 127204 154006
rect 127164 153944 127216 153950
rect 127164 153886 127216 153892
rect 127544 150226 127572 155994
rect 127820 153105 127848 159423
rect 127900 158024 127952 158030
rect 127900 157966 127952 157972
rect 127912 154018 127940 157966
rect 128188 156806 128216 163200
rect 128176 156800 128228 156806
rect 128176 156742 128228 156748
rect 129016 155242 129044 163200
rect 129740 158772 129792 158778
rect 129740 158714 129792 158720
rect 129004 155236 129056 155242
rect 129004 155178 129056 155184
rect 128360 154692 128412 154698
rect 128360 154634 128412 154640
rect 127900 154012 127952 154018
rect 127900 153954 127952 153960
rect 127806 153096 127862 153105
rect 127806 153031 127862 153040
rect 128372 151978 128400 154634
rect 129464 153944 129516 153950
rect 129464 153886 129516 153892
rect 128818 152552 128874 152561
rect 128818 152487 128874 152496
rect 128176 151972 128228 151978
rect 128176 151914 128228 151920
rect 128360 151972 128412 151978
rect 128360 151914 128412 151920
rect 128188 150226 128216 151914
rect 128832 150226 128860 152487
rect 129476 150226 129504 153886
rect 129752 152522 129780 158714
rect 129936 153950 129964 163200
rect 130764 158914 130792 163200
rect 130752 158908 130804 158914
rect 130752 158850 130804 158856
rect 131592 158030 131620 163200
rect 131580 158024 131632 158030
rect 131580 157966 131632 157972
rect 132420 156738 132448 163200
rect 133248 158778 133276 163200
rect 133236 158772 133288 158778
rect 133236 158714 133288 158720
rect 132500 156936 132552 156942
rect 132500 156878 132552 156884
rect 130108 156732 130160 156738
rect 130108 156674 130160 156680
rect 132408 156732 132460 156738
rect 132408 156674 132460 156680
rect 129924 153944 129976 153950
rect 129924 153886 129976 153892
rect 129740 152516 129792 152522
rect 129740 152458 129792 152464
rect 130120 150226 130148 156674
rect 132038 153776 132094 153785
rect 132038 153711 132094 153720
rect 131394 153096 131450 153105
rect 131394 153031 131450 153040
rect 130752 152652 130804 152658
rect 130752 152594 130804 152600
rect 130764 150226 130792 152594
rect 131408 150226 131436 153031
rect 132052 150226 132080 153711
rect 132512 151814 132540 156878
rect 134076 155446 134104 163200
rect 134904 156942 134932 163200
rect 135168 159452 135220 159458
rect 135168 159394 135220 159400
rect 134892 156936 134944 156942
rect 134892 156878 134944 156884
rect 134064 155440 134116 155446
rect 134064 155382 134116 155388
rect 133328 154760 133380 154766
rect 133328 154702 133380 154708
rect 132512 151786 132724 151814
rect 132696 150226 132724 151786
rect 133340 150226 133368 154702
rect 134614 153912 134670 153921
rect 134614 153847 134670 153856
rect 133972 152584 134024 152590
rect 133972 152526 134024 152532
rect 133984 150226 134012 152526
rect 134628 150226 134656 153847
rect 135180 152658 135208 159394
rect 135260 156868 135312 156874
rect 135260 156810 135312 156816
rect 135168 152652 135220 152658
rect 135168 152594 135220 152600
rect 135272 150226 135300 156810
rect 135824 156058 135852 163200
rect 136652 160138 136680 163200
rect 136640 160132 136692 160138
rect 136640 160074 136692 160080
rect 136548 159860 136600 159866
rect 136548 159802 136600 159808
rect 136560 159526 136588 159802
rect 136548 159520 136600 159526
rect 136548 159462 136600 159468
rect 137374 159488 137430 159497
rect 137480 159458 137508 163200
rect 137652 159724 137704 159730
rect 137652 159666 137704 159672
rect 137374 159423 137376 159432
rect 137428 159423 137430 159432
rect 137468 159452 137520 159458
rect 137376 159394 137428 159400
rect 137468 159394 137520 159400
rect 136546 159352 136602 159361
rect 136546 159287 136602 159296
rect 135812 156052 135864 156058
rect 135812 155994 135864 156000
rect 135904 152720 135956 152726
rect 135904 152662 135956 152668
rect 135916 150226 135944 152662
rect 136560 150226 136588 159287
rect 136916 157004 136968 157010
rect 136916 156946 136968 156952
rect 136928 152658 136956 156946
rect 137560 155440 137612 155446
rect 137560 155382 137612 155388
rect 137100 154284 137152 154290
rect 137100 154226 137152 154232
rect 137008 154216 137060 154222
rect 137008 154158 137060 154164
rect 136916 152652 136968 152658
rect 136916 152594 136968 152600
rect 137020 151814 137048 154158
rect 137112 154034 137140 154226
rect 137468 154080 137520 154086
rect 137112 154028 137468 154034
rect 137112 154022 137520 154028
rect 137112 154006 137508 154022
rect 137192 152652 137244 152658
rect 137192 152594 137244 152600
rect 137204 151814 137232 152594
rect 137572 152522 137600 155382
rect 137664 154086 137692 159666
rect 138308 157010 138336 163200
rect 138570 159488 138626 159497
rect 138570 159423 138626 159432
rect 138296 157004 138348 157010
rect 138296 156946 138348 156952
rect 137652 154080 137704 154086
rect 137652 154022 137704 154028
rect 137560 152516 137612 152522
rect 137560 152458 137612 152464
rect 138584 151842 138612 159423
rect 139136 156874 139164 163200
rect 139398 159624 139454 159633
rect 139398 159559 139454 159568
rect 139858 159624 139914 159633
rect 139964 159594 139992 163200
rect 139858 159559 139860 159568
rect 139124 156868 139176 156874
rect 139124 156810 139176 156816
rect 139412 152794 139440 159559
rect 139912 159559 139914 159568
rect 139952 159588 140004 159594
rect 139860 159530 139912 159536
rect 139952 159530 140004 159536
rect 139950 156632 140006 156641
rect 139950 156567 140006 156576
rect 139766 154048 139822 154057
rect 139766 153983 139822 153992
rect 139124 152788 139176 152794
rect 139124 152730 139176 152736
rect 139400 152788 139452 152794
rect 139400 152730 139452 152736
rect 138480 151836 138532 151842
rect 137020 151786 137140 151814
rect 137204 151786 137876 151814
rect 137112 150226 137140 151786
rect 137848 150226 137876 151786
rect 138480 151778 138532 151784
rect 138572 151836 138624 151842
rect 138572 151778 138624 151784
rect 138492 150226 138520 151778
rect 139136 150226 139164 152730
rect 139780 150226 139808 153983
rect 139964 151814 139992 156567
rect 140792 152590 140820 163200
rect 141712 157418 141740 163200
rect 142252 159656 142304 159662
rect 142252 159598 142304 159604
rect 141700 157412 141752 157418
rect 141700 157354 141752 157360
rect 141700 152788 141752 152794
rect 141700 152730 141752 152736
rect 140780 152584 140832 152590
rect 140780 152526 140832 152532
rect 141148 152516 141200 152522
rect 141148 152458 141200 152464
rect 141160 152318 141188 152458
rect 141056 152312 141108 152318
rect 141056 152254 141108 152260
rect 141148 152312 141200 152318
rect 141148 152254 141200 152260
rect 139964 151786 140452 151814
rect 140424 150226 140452 151786
rect 141068 150226 141096 152254
rect 141712 150226 141740 152730
rect 141884 152720 141936 152726
rect 141884 152662 141936 152668
rect 141896 151842 141924 152662
rect 142264 151842 142292 159598
rect 142540 155310 142568 163200
rect 142620 159860 142672 159866
rect 142620 159802 142672 159808
rect 142632 159390 142660 159802
rect 143368 159662 143396 163200
rect 143356 159656 143408 159662
rect 143356 159598 143408 159604
rect 144196 159526 144224 163200
rect 144276 160132 144328 160138
rect 144276 160074 144328 160080
rect 144288 159730 144316 160074
rect 144276 159724 144328 159730
rect 144276 159666 144328 159672
rect 144918 159624 144974 159633
rect 144918 159559 144974 159568
rect 144184 159520 144236 159526
rect 144184 159462 144236 159468
rect 144932 159458 144960 159559
rect 144828 159452 144880 159458
rect 144828 159394 144880 159400
rect 144920 159452 144972 159458
rect 144920 159394 144972 159400
rect 142620 159384 142672 159390
rect 142620 159326 142672 159332
rect 142710 156768 142766 156777
rect 142710 156703 142766 156712
rect 142528 155304 142580 155310
rect 142528 155246 142580 155252
rect 142344 154012 142396 154018
rect 142344 153954 142396 153960
rect 141884 151836 141936 151842
rect 141884 151778 141936 151784
rect 142252 151836 142304 151842
rect 142252 151778 142304 151784
rect 142356 150226 142384 153954
rect 142724 151814 142752 156703
rect 143630 152688 143686 152697
rect 143630 152623 143686 152632
rect 142724 151786 143028 151814
rect 143000 150226 143028 151786
rect 143644 150226 143672 152623
rect 144840 152454 144868 159394
rect 144918 157992 144974 158001
rect 144918 157927 144974 157936
rect 144276 152448 144328 152454
rect 144276 152390 144328 152396
rect 144828 152448 144880 152454
rect 144828 152390 144880 152396
rect 144288 150226 144316 152390
rect 144932 150226 144960 157927
rect 145024 155990 145052 163200
rect 145472 157072 145524 157078
rect 145472 157014 145524 157020
rect 145012 155984 145064 155990
rect 145012 155926 145064 155932
rect 145380 154420 145432 154426
rect 145380 154362 145432 154368
rect 145104 154352 145156 154358
rect 145104 154294 145156 154300
rect 145116 154018 145144 154294
rect 145104 154012 145156 154018
rect 145104 153954 145156 153960
rect 145392 150498 145420 154362
rect 145484 151814 145512 157014
rect 145852 155378 145880 163200
rect 146680 161430 146708 163200
rect 146668 161424 146720 161430
rect 146668 161366 146720 161372
rect 146300 159860 146352 159866
rect 146300 159802 146352 159808
rect 146312 159458 146340 159802
rect 146852 159792 146904 159798
rect 146852 159734 146904 159740
rect 146208 159452 146260 159458
rect 146208 159394 146260 159400
rect 146300 159452 146352 159458
rect 146300 159394 146352 159400
rect 145840 155372 145892 155378
rect 145840 155314 145892 155320
rect 146220 154630 146248 159394
rect 146392 158092 146444 158098
rect 146392 158034 146444 158040
rect 146208 154624 146260 154630
rect 146208 154566 146260 154572
rect 145484 151786 146248 151814
rect 145392 150470 145604 150498
rect 145576 150226 145604 150470
rect 146220 150226 146248 151786
rect 126256 150198 126330 150226
rect 126900 150198 126974 150226
rect 127544 150198 127618 150226
rect 128188 150198 128262 150226
rect 128832 150198 128906 150226
rect 129476 150198 129550 150226
rect 130120 150198 130194 150226
rect 130764 150198 130838 150226
rect 131408 150198 131482 150226
rect 132052 150198 132126 150226
rect 132696 150198 132770 150226
rect 133340 150198 133414 150226
rect 133984 150198 134058 150226
rect 134628 150198 134702 150226
rect 135272 150198 135346 150226
rect 135916 150198 135990 150226
rect 136560 150198 136634 150226
rect 137112 150198 137278 150226
rect 137848 150198 137922 150226
rect 138492 150198 138566 150226
rect 139136 150198 139210 150226
rect 139780 150198 139854 150226
rect 140424 150198 140498 150226
rect 141068 150198 141142 150226
rect 141712 150198 141786 150226
rect 142356 150198 142430 150226
rect 143000 150198 143074 150226
rect 143644 150198 143718 150226
rect 144288 150198 144362 150226
rect 144932 150198 145006 150226
rect 145576 150198 145650 150226
rect 146220 150198 146294 150226
rect 146404 150210 146432 158034
rect 146864 157078 146892 159734
rect 147600 159458 147628 163200
rect 147128 159452 147180 159458
rect 147128 159394 147180 159400
rect 147588 159452 147640 159458
rect 147588 159394 147640 159400
rect 146852 157072 146904 157078
rect 146852 157014 146904 157020
rect 146484 154556 146536 154562
rect 146484 154498 146536 154504
rect 146496 154442 146524 154498
rect 146496 154414 147076 154442
rect 146944 154352 146996 154358
rect 146944 154294 146996 154300
rect 146956 154170 146984 154294
rect 146864 154154 146984 154170
rect 147048 154154 147076 154414
rect 147140 154222 147168 159394
rect 148428 158098 148456 163200
rect 148692 159928 148744 159934
rect 148692 159870 148744 159876
rect 148600 159792 148652 159798
rect 148600 159734 148652 159740
rect 148612 159662 148640 159734
rect 148600 159656 148652 159662
rect 148600 159598 148652 159604
rect 148704 159576 148732 159870
rect 148796 159730 149008 159746
rect 148784 159724 149020 159730
rect 148836 159718 148968 159724
rect 148784 159666 148836 159672
rect 148968 159666 149020 159672
rect 148704 159548 149192 159576
rect 149164 159458 149192 159548
rect 149060 159452 149112 159458
rect 149060 159394 149112 159400
rect 149152 159452 149204 159458
rect 149152 159394 149204 159400
rect 148416 158092 148468 158098
rect 148416 158034 148468 158040
rect 147680 157140 147732 157146
rect 147680 157082 147732 157088
rect 147128 154216 147180 154222
rect 147128 154158 147180 154164
rect 146852 154148 146984 154154
rect 146904 154142 146984 154148
rect 147036 154148 147088 154154
rect 146852 154090 146904 154096
rect 147036 154090 147088 154096
rect 146852 152788 146904 152794
rect 146852 152730 146904 152736
rect 146864 150226 146892 152730
rect 146944 152584 146996 152590
rect 146944 152526 146996 152532
rect 146956 152318 146984 152526
rect 146944 152312 146996 152318
rect 146944 152254 146996 152260
rect 125658 149940 125686 150198
rect 126302 149940 126330 150198
rect 126946 149940 126974 150198
rect 127590 149940 127618 150198
rect 128234 149940 128262 150198
rect 128878 149940 128906 150198
rect 129522 149940 129550 150198
rect 130166 149940 130194 150198
rect 130810 149940 130838 150198
rect 131454 149940 131482 150198
rect 132098 149940 132126 150198
rect 132742 149940 132770 150198
rect 133386 149940 133414 150198
rect 134030 149940 134058 150198
rect 134674 149940 134702 150198
rect 135318 149940 135346 150198
rect 135962 149940 135990 150198
rect 136606 149940 136634 150198
rect 137250 149940 137278 150198
rect 137894 149940 137922 150198
rect 138538 149940 138566 150198
rect 139182 149940 139210 150198
rect 139826 149940 139854 150198
rect 140470 149940 140498 150198
rect 141114 149940 141142 150198
rect 141758 149940 141786 150198
rect 142402 149940 142430 150198
rect 143046 149940 143074 150198
rect 143690 149940 143718 150198
rect 144334 149940 144362 150198
rect 144978 149940 145006 150198
rect 145622 149940 145650 150198
rect 146266 149940 146294 150198
rect 146392 150204 146444 150210
rect 146864 150198 146938 150226
rect 147692 150210 147720 157082
rect 148140 154080 148192 154086
rect 148140 154022 148192 154028
rect 148152 150226 148180 154022
rect 149072 152794 149100 159394
rect 149256 155446 149284 163200
rect 149610 158128 149666 158137
rect 149610 158063 149666 158072
rect 149244 155440 149296 155446
rect 149244 155382 149296 155388
rect 149060 152788 149112 152794
rect 149060 152730 149112 152736
rect 149428 152040 149480 152046
rect 149428 151982 149480 151988
rect 149440 150226 149468 151982
rect 149624 151814 149652 158063
rect 150084 154154 150112 163200
rect 150808 159792 150860 159798
rect 150808 159734 150860 159740
rect 150820 159458 150848 159734
rect 150912 159458 150940 163200
rect 150808 159452 150860 159458
rect 150808 159394 150860 159400
rect 150900 159452 150952 159458
rect 150900 159394 150952 159400
rect 151740 157078 151768 163200
rect 150440 157072 150492 157078
rect 150440 157014 150492 157020
rect 151728 157072 151780 157078
rect 151728 157014 151780 157020
rect 150072 154148 150124 154154
rect 150072 154090 150124 154096
rect 150452 152318 150480 157014
rect 150990 156904 151046 156913
rect 150990 156839 151046 156848
rect 150624 154556 150676 154562
rect 150624 154498 150676 154504
rect 150440 152312 150492 152318
rect 150440 152254 150492 152260
rect 149624 151786 150020 151814
rect 149992 150226 150020 151786
rect 150636 150226 150664 154498
rect 151004 151814 151032 156839
rect 151832 154630 151860 163254
rect 152476 163146 152504 163254
rect 152554 163200 152610 164400
rect 153474 163200 153530 164400
rect 153580 163254 154252 163282
rect 152568 163146 152596 163200
rect 152476 163118 152596 163146
rect 152464 159928 152516 159934
rect 152464 159870 152516 159876
rect 152476 159322 152504 159870
rect 153488 159798 153516 163200
rect 152556 159792 152608 159798
rect 152556 159734 152608 159740
rect 153476 159792 153528 159798
rect 153476 159734 153528 159740
rect 152568 159322 152596 159734
rect 152464 159316 152516 159322
rect 152464 159258 152516 159264
rect 152556 159316 152608 159322
rect 152556 159258 152608 159264
rect 152554 158264 152610 158273
rect 152554 158199 152610 158208
rect 151820 154624 151872 154630
rect 151820 154566 151872 154572
rect 151912 152720 151964 152726
rect 151912 152662 151964 152668
rect 151004 151786 151308 151814
rect 151280 150226 151308 151786
rect 151924 150226 151952 152662
rect 152568 150226 152596 158199
rect 152740 154216 152792 154222
rect 152740 154158 152792 154164
rect 153292 154216 153344 154222
rect 153292 154158 153344 154164
rect 152648 154080 152700 154086
rect 152648 154022 152700 154028
rect 152660 153814 152688 154022
rect 152752 153814 152780 154158
rect 153200 154012 153252 154018
rect 153200 153954 153252 153960
rect 152648 153808 152700 153814
rect 152648 153750 152700 153756
rect 152740 153808 152792 153814
rect 152740 153750 152792 153756
rect 153212 150226 153240 153954
rect 153304 153746 153332 154158
rect 153292 153740 153344 153746
rect 153292 153682 153344 153688
rect 153580 152726 153608 163254
rect 154224 163146 154252 163254
rect 154302 163200 154358 164400
rect 155130 163200 155186 164400
rect 155958 163200 156014 164400
rect 156786 163200 156842 164400
rect 157614 163200 157670 164400
rect 158442 163200 158498 164400
rect 159362 163200 159418 164400
rect 160190 163200 160246 164400
rect 161018 163200 161074 164400
rect 161846 163200 161902 164400
rect 162674 163200 162730 164400
rect 163502 163200 163558 164400
rect 164330 163200 164386 164400
rect 165250 163200 165306 164400
rect 166078 163200 166134 164400
rect 166184 163254 166396 163282
rect 154316 163146 154344 163200
rect 154224 163118 154344 163146
rect 153752 161424 153804 161430
rect 153752 161366 153804 161372
rect 153764 159866 153792 161366
rect 153752 159860 153804 159866
rect 153752 159802 153804 159808
rect 154488 158840 154540 158846
rect 154488 158782 154540 158788
rect 153752 157208 153804 157214
rect 153752 157150 153804 157156
rect 153568 152720 153620 152726
rect 153568 152662 153620 152668
rect 153764 151814 153792 157150
rect 154500 153746 154528 158782
rect 155144 158166 155172 163200
rect 155040 158160 155092 158166
rect 155040 158102 155092 158108
rect 155132 158160 155184 158166
rect 155132 158102 155184 158108
rect 154488 153740 154540 153746
rect 154488 153682 154540 153688
rect 154488 152108 154540 152114
rect 154488 152050 154540 152056
rect 153764 151786 153884 151814
rect 153856 150226 153884 151786
rect 154500 150226 154528 152050
rect 155052 151814 155080 158102
rect 155972 154766 156000 163200
rect 156052 159316 156104 159322
rect 156052 159258 156104 159264
rect 155960 154760 156012 154766
rect 155960 154702 156012 154708
rect 155776 154080 155828 154086
rect 155776 154022 155828 154028
rect 155052 151786 155172 151814
rect 155144 150226 155172 151786
rect 155788 150226 155816 154022
rect 156064 152114 156092 159258
rect 156800 158846 156828 163200
rect 157246 159624 157302 159633
rect 157628 159594 157656 163200
rect 157246 159559 157248 159568
rect 157300 159559 157302 159568
rect 157616 159588 157668 159594
rect 157248 159530 157300 159536
rect 157616 159530 157668 159536
rect 157338 159488 157394 159497
rect 157338 159423 157394 159432
rect 156788 158840 156840 158846
rect 156788 158782 156840 158788
rect 156418 157040 156474 157049
rect 156418 156975 156474 156984
rect 156052 152108 156104 152114
rect 156052 152050 156104 152056
rect 156432 150226 156460 156975
rect 157352 154562 157380 159423
rect 158456 158234 158484 163200
rect 158720 158772 158772 158778
rect 158720 158714 158772 158720
rect 157708 158228 157760 158234
rect 157708 158170 157760 158176
rect 158444 158228 158496 158234
rect 158444 158170 158496 158176
rect 156604 154556 156656 154562
rect 156604 154498 156656 154504
rect 156788 154556 156840 154562
rect 156788 154498 156840 154504
rect 157340 154556 157392 154562
rect 157340 154498 157392 154504
rect 156616 153746 156644 154498
rect 156800 154086 156828 154498
rect 156880 154148 156932 154154
rect 156880 154090 156932 154096
rect 156788 154080 156840 154086
rect 156788 154022 156840 154028
rect 156892 153898 156920 154090
rect 156708 153870 156920 153898
rect 156512 153740 156564 153746
rect 156512 153682 156564 153688
rect 156604 153740 156656 153746
rect 156604 153682 156656 153688
rect 156524 153626 156552 153682
rect 156708 153626 156736 153870
rect 156524 153598 156736 153626
rect 157064 151836 157116 151842
rect 157064 151778 157116 151784
rect 157076 150226 157104 151778
rect 157720 150226 157748 158170
rect 158732 157350 158760 158714
rect 158628 157344 158680 157350
rect 158628 157286 158680 157292
rect 158720 157344 158772 157350
rect 158720 157286 158772 157292
rect 158640 157162 158668 157286
rect 158640 157134 158760 157162
rect 158350 154184 158406 154193
rect 158350 154119 158406 154128
rect 158364 150226 158392 154119
rect 158732 151814 158760 157134
rect 159376 154630 159404 163200
rect 160204 159934 160232 163200
rect 160100 159928 160152 159934
rect 160100 159870 160152 159876
rect 160192 159928 160244 159934
rect 160192 159870 160244 159876
rect 160112 159746 160140 159870
rect 160112 159718 160232 159746
rect 160100 159656 160152 159662
rect 160100 159598 160152 159604
rect 160112 157214 160140 159598
rect 160100 157208 160152 157214
rect 160100 157150 160152 157156
rect 159364 154624 159416 154630
rect 159364 154566 159416 154572
rect 160204 152250 160232 159718
rect 161032 159662 161060 163200
rect 161020 159656 161072 159662
rect 161020 159598 161072 159604
rect 161860 158302 161888 163200
rect 160284 158296 160336 158302
rect 160284 158238 160336 158244
rect 161848 158296 161900 158302
rect 161848 158238 161900 158244
rect 159640 152244 159692 152250
rect 159640 152186 159692 152192
rect 160192 152244 160244 152250
rect 160192 152186 160244 152192
rect 158732 151786 159036 151814
rect 159008 150226 159036 151786
rect 159652 150226 159680 152186
rect 160296 150226 160324 158238
rect 161572 157276 161624 157282
rect 161572 157218 161624 157224
rect 160926 154320 160982 154329
rect 160926 154255 160982 154264
rect 160940 150226 160968 154255
rect 161584 150226 161612 157218
rect 162688 154698 162716 163200
rect 163516 159322 163544 163200
rect 164148 159724 164200 159730
rect 164148 159666 164200 159672
rect 163504 159316 163556 159322
rect 163504 159258 163556 159264
rect 163044 158704 163096 158710
rect 163228 158704 163280 158710
rect 163096 158652 163228 158658
rect 163044 158646 163280 158652
rect 163056 158630 163268 158646
rect 163320 158636 163372 158642
rect 163320 158578 163372 158584
rect 163332 158438 163360 158578
rect 163320 158432 163372 158438
rect 162858 158400 162914 158409
rect 163320 158374 163372 158380
rect 162858 158335 162914 158344
rect 162676 154692 162728 154698
rect 162676 154634 162728 154640
rect 162216 152448 162268 152454
rect 162216 152390 162268 152396
rect 162228 150226 162256 152390
rect 162872 150226 162900 158335
rect 164160 156754 164188 159666
rect 164160 156726 164280 156754
rect 164252 156602 164280 156726
rect 164148 156596 164200 156602
rect 164148 156538 164200 156544
rect 164240 156596 164292 156602
rect 164240 156538 164292 156544
rect 163504 154216 163556 154222
rect 163504 154158 163556 154164
rect 163516 150226 163544 154158
rect 164160 150226 164188 156538
rect 164344 152454 164372 163200
rect 165264 158370 165292 163200
rect 166092 163146 166120 163200
rect 166184 163146 166212 163254
rect 166092 163118 166212 163146
rect 165436 158432 165488 158438
rect 165436 158374 165488 158380
rect 165252 158364 165304 158370
rect 165252 158306 165304 158312
rect 165068 154216 165120 154222
rect 165068 154158 165120 154164
rect 165080 153678 165108 154158
rect 165068 153672 165120 153678
rect 165068 153614 165120 153620
rect 164332 152448 164384 152454
rect 164332 152390 164384 152396
rect 164792 152176 164844 152182
rect 164792 152118 164844 152124
rect 164804 150226 164832 152118
rect 165448 150226 165476 158374
rect 165712 155508 165764 155514
rect 165712 155450 165764 155456
rect 146392 150146 146444 150152
rect 146910 149940 146938 150198
rect 147542 150204 147594 150210
rect 147542 150146 147594 150152
rect 147680 150204 147732 150210
rect 148152 150198 148226 150226
rect 147680 150146 147732 150152
rect 147554 149940 147582 150146
rect 148198 149940 148226 150198
rect 148830 150204 148882 150210
rect 149440 150198 149514 150226
rect 149992 150198 150066 150226
rect 150636 150198 150710 150226
rect 151280 150198 151354 150226
rect 151924 150198 151998 150226
rect 152568 150198 152642 150226
rect 153212 150198 153286 150226
rect 153856 150198 153930 150226
rect 154500 150198 154574 150226
rect 155144 150198 155218 150226
rect 155788 150198 155862 150226
rect 156432 150198 156506 150226
rect 157076 150198 157150 150226
rect 157720 150198 157794 150226
rect 158364 150198 158438 150226
rect 159008 150198 159082 150226
rect 159652 150198 159726 150226
rect 160296 150198 160370 150226
rect 160940 150198 161014 150226
rect 161584 150198 161658 150226
rect 162228 150198 162302 150226
rect 162872 150198 162946 150226
rect 163516 150198 163590 150226
rect 164160 150198 164234 150226
rect 164804 150198 164878 150226
rect 165448 150198 165522 150226
rect 165724 150210 165752 155450
rect 166078 155272 166134 155281
rect 166078 155207 166134 155216
rect 166092 150226 166120 155207
rect 166368 154154 166396 163254
rect 166906 163200 166962 164400
rect 167734 163200 167790 164400
rect 168562 163200 168618 164400
rect 169390 163200 169446 164400
rect 170218 163200 170274 164400
rect 171138 163200 171194 164400
rect 171966 163200 172022 164400
rect 172532 163254 172744 163282
rect 166920 157146 166948 163200
rect 167000 160064 167052 160070
rect 167000 160006 167052 160012
rect 166908 157140 166960 157146
rect 166908 157082 166960 157088
rect 166264 154148 166316 154154
rect 166264 154090 166316 154096
rect 166356 154148 166408 154154
rect 166356 154090 166408 154096
rect 166276 153678 166304 154090
rect 166264 153672 166316 153678
rect 166264 153614 166316 153620
rect 167012 152182 167040 160006
rect 167748 159730 167776 163200
rect 167736 159724 167788 159730
rect 167736 159666 167788 159672
rect 167644 158704 167696 158710
rect 167828 158704 167880 158710
rect 167696 158652 167828 158658
rect 167644 158646 167880 158652
rect 167552 158636 167604 158642
rect 167656 158630 167868 158646
rect 167552 158578 167604 158584
rect 167368 152312 167420 152318
rect 167368 152254 167420 152260
rect 167000 152176 167052 152182
rect 167000 152118 167052 152124
rect 167380 150226 167408 152254
rect 167564 151814 167592 158578
rect 168576 158438 168604 163200
rect 168564 158432 168616 158438
rect 168564 158374 168616 158380
rect 169298 157176 169354 157185
rect 169298 157111 169354 157120
rect 168656 154216 168708 154222
rect 168656 154158 168708 154164
rect 167564 151786 168052 151814
rect 168024 150226 168052 151786
rect 168668 150226 168696 154158
rect 169312 150226 169340 157111
rect 169404 155514 169432 163200
rect 170232 160070 170260 163200
rect 170220 160064 170272 160070
rect 170220 160006 170272 160012
rect 169760 159180 169812 159186
rect 169760 159122 169812 159128
rect 169392 155508 169444 155514
rect 169392 155450 169444 155456
rect 169772 152046 169800 159122
rect 171152 158778 171180 163200
rect 171140 158772 171192 158778
rect 171140 158714 171192 158720
rect 171980 158642 172008 163200
rect 170312 158636 170364 158642
rect 170312 158578 170364 158584
rect 171968 158636 172020 158642
rect 171968 158578 172020 158584
rect 169944 152856 169996 152862
rect 169944 152798 169996 152804
rect 169760 152040 169812 152046
rect 169760 151982 169812 151988
rect 169956 150226 169984 152798
rect 170324 151814 170352 158578
rect 171138 155544 171194 155553
rect 171138 155479 171194 155488
rect 170324 151786 170628 151814
rect 170600 150226 170628 151786
rect 148830 150146 148882 150152
rect 148842 149940 148870 150146
rect 149486 149940 149514 150198
rect 150038 149940 150066 150198
rect 150682 149940 150710 150198
rect 151326 149940 151354 150198
rect 151970 149940 151998 150198
rect 152614 149940 152642 150198
rect 153258 149940 153286 150198
rect 153902 149940 153930 150198
rect 154546 149940 154574 150198
rect 155190 149940 155218 150198
rect 155834 149940 155862 150198
rect 156478 149940 156506 150198
rect 157122 149940 157150 150198
rect 157766 149940 157794 150198
rect 158410 149940 158438 150198
rect 159054 149940 159082 150198
rect 159698 149940 159726 150198
rect 160342 149940 160370 150198
rect 160986 149940 161014 150198
rect 161630 149940 161658 150198
rect 162274 149940 162302 150198
rect 162918 149940 162946 150198
rect 163562 149940 163590 150198
rect 164206 149940 164234 150198
rect 164850 149940 164878 150198
rect 165494 149940 165522 150198
rect 165712 150204 165764 150210
rect 166092 150198 166166 150226
rect 165712 150146 165764 150152
rect 166138 149940 166166 150198
rect 166770 150204 166822 150210
rect 167380 150198 167454 150226
rect 168024 150198 168098 150226
rect 168668 150198 168742 150226
rect 169312 150198 169386 150226
rect 169956 150198 170030 150226
rect 170600 150198 170674 150226
rect 171152 150210 171180 155479
rect 171230 155408 171286 155417
rect 171230 155343 171286 155352
rect 171244 150226 171272 155343
rect 172532 154222 172560 163254
rect 172716 163146 172744 163254
rect 172794 163200 172850 164400
rect 173622 163200 173678 164400
rect 173912 163254 174400 163282
rect 172808 163146 172836 163200
rect 172716 163118 172836 163146
rect 173636 159186 173664 163200
rect 173624 159180 173676 159186
rect 173624 159122 173676 159128
rect 172612 158772 172664 158778
rect 172612 158714 172664 158720
rect 172520 154216 172572 154222
rect 172520 154158 172572 154164
rect 172624 152318 172652 158714
rect 173072 158500 173124 158506
rect 173072 158442 173124 158448
rect 172704 155712 172756 155718
rect 172704 155654 172756 155660
rect 172612 152312 172664 152318
rect 172612 152254 172664 152260
rect 172520 152108 172572 152114
rect 172520 152050 172572 152056
rect 172532 150226 172560 152050
rect 166770 150146 166822 150152
rect 166782 149940 166810 150146
rect 167426 149940 167454 150198
rect 168070 149940 168098 150198
rect 168714 149940 168742 150198
rect 169358 149940 169386 150198
rect 170002 149940 170030 150198
rect 170646 149940 170674 150198
rect 171140 150204 171192 150210
rect 171244 150198 171318 150226
rect 171140 150146 171192 150152
rect 171290 149940 171318 150198
rect 171922 150204 171974 150210
rect 172532 150198 172606 150226
rect 172716 150210 172744 155654
rect 173084 151814 173112 158442
rect 173912 152862 173940 163254
rect 174372 163146 174400 163254
rect 174450 163200 174506 164400
rect 175278 163200 175334 164400
rect 176106 163200 176162 164400
rect 177026 163200 177082 164400
rect 177854 163200 177910 164400
rect 178682 163200 178738 164400
rect 179510 163200 179566 164400
rect 180338 163200 180394 164400
rect 180812 163254 181116 163282
rect 174464 163146 174492 163200
rect 174372 163118 174492 163146
rect 175004 159860 175056 159866
rect 175004 159802 175056 159808
rect 175016 156534 175044 159802
rect 175292 158574 175320 163200
rect 176120 161474 176148 163200
rect 176120 161446 176332 161474
rect 175832 159248 175884 159254
rect 175832 159190 175884 159196
rect 175844 158778 175872 159190
rect 175936 159186 176148 159202
rect 175924 159180 176160 159186
rect 175976 159174 176108 159180
rect 175924 159122 175976 159128
rect 176108 159122 176160 159128
rect 175832 158772 175884 158778
rect 175832 158714 175884 158720
rect 175280 158568 175332 158574
rect 175280 158510 175332 158516
rect 175372 158500 175424 158506
rect 175372 158442 175424 158448
rect 174452 156528 174504 156534
rect 174452 156470 174504 156476
rect 175004 156528 175056 156534
rect 175004 156470 175056 156476
rect 173900 152856 173952 152862
rect 173900 152798 173952 152804
rect 173084 151786 173204 151814
rect 173176 150226 173204 151786
rect 174464 150226 174492 156470
rect 175096 151904 175148 151910
rect 175096 151846 175148 151852
rect 175108 150226 175136 151846
rect 175384 151814 175412 158442
rect 176200 157956 176252 157962
rect 176200 157898 176252 157904
rect 175924 157888 175976 157894
rect 176212 157842 176240 157898
rect 175976 157836 176240 157842
rect 175924 157830 176240 157836
rect 175936 157814 176240 157830
rect 176304 155718 176332 161446
rect 176660 158772 176712 158778
rect 176660 158714 176712 158720
rect 176292 155712 176344 155718
rect 176292 155654 176344 155660
rect 176384 155644 176436 155650
rect 176384 155586 176436 155592
rect 175384 151786 175780 151814
rect 175752 150226 175780 151786
rect 176396 150226 176424 155586
rect 176672 151910 176700 158714
rect 177040 157334 177068 163200
rect 177868 159798 177896 163200
rect 177856 159792 177908 159798
rect 177856 159734 177908 159740
rect 178696 158506 178724 163200
rect 178684 158500 178736 158506
rect 178684 158442 178736 158448
rect 178040 157888 178092 157894
rect 178040 157830 178092 157836
rect 177040 157306 177160 157334
rect 177026 155680 177082 155689
rect 177132 155650 177160 157306
rect 177026 155615 177082 155624
rect 177120 155644 177172 155650
rect 176660 151904 176712 151910
rect 176660 151846 176712 151852
rect 177040 150226 177068 155615
rect 177120 155586 177172 155592
rect 177672 152244 177724 152250
rect 177672 152186 177724 152192
rect 177684 150226 177712 152186
rect 178052 151814 178080 157830
rect 179524 155582 179552 163200
rect 180352 159118 180380 163200
rect 180708 159860 180760 159866
rect 180708 159802 180760 159808
rect 180340 159112 180392 159118
rect 180340 159054 180392 159060
rect 180720 158778 180748 159802
rect 180708 158772 180760 158778
rect 180708 158714 180760 158720
rect 179604 156460 179656 156466
rect 179604 156402 179656 156408
rect 178960 155576 179012 155582
rect 178960 155518 179012 155524
rect 179512 155576 179564 155582
rect 179512 155518 179564 155524
rect 178052 151786 178356 151814
rect 178328 150226 178356 151786
rect 178972 150226 179000 155518
rect 179616 150226 179644 156402
rect 180812 153134 180840 163254
rect 181088 163146 181116 163254
rect 181166 163200 181222 164400
rect 181994 163200 182050 164400
rect 182192 163254 182864 163282
rect 181180 163146 181208 163200
rect 181088 163118 181208 163146
rect 182008 158710 182036 163200
rect 180892 158704 180944 158710
rect 180892 158646 180944 158652
rect 181720 158704 181772 158710
rect 181720 158646 181772 158652
rect 181996 158704 182048 158710
rect 181996 158646 182048 158652
rect 180248 153128 180300 153134
rect 180248 153070 180300 153076
rect 180800 153128 180852 153134
rect 180800 153070 180852 153076
rect 180260 150226 180288 153070
rect 180904 150226 180932 158646
rect 181352 157820 181404 157826
rect 181352 157762 181404 157768
rect 181364 157706 181392 157762
rect 181732 157758 181760 158646
rect 181720 157752 181772 157758
rect 181364 157690 181668 157706
rect 181720 157694 181772 157700
rect 181364 157684 181680 157690
rect 181364 157678 181628 157684
rect 181628 157626 181680 157632
rect 181444 155780 181496 155786
rect 181444 155722 181496 155728
rect 171922 150146 171974 150152
rect 171934 149940 171962 150146
rect 172578 149940 172606 150198
rect 172704 150204 172756 150210
rect 173176 150198 173250 150226
rect 172704 150146 172756 150152
rect 173222 149940 173250 150198
rect 173854 150204 173906 150210
rect 174464 150198 174538 150226
rect 175108 150198 175182 150226
rect 175752 150198 175826 150226
rect 176396 150198 176470 150226
rect 177040 150198 177114 150226
rect 177684 150198 177758 150226
rect 178328 150198 178402 150226
rect 178972 150198 179046 150226
rect 179616 150198 179690 150226
rect 180260 150198 180334 150226
rect 173854 150146 173906 150152
rect 173866 149940 173894 150146
rect 174510 149940 174538 150198
rect 175154 149940 175182 150198
rect 175798 149940 175826 150198
rect 176442 149940 176470 150198
rect 177086 149940 177114 150198
rect 177730 149940 177758 150198
rect 178374 149940 178402 150198
rect 179018 149940 179046 150198
rect 179662 149940 179690 150198
rect 180306 149940 180334 150198
rect 180858 150198 180932 150226
rect 181456 150226 181484 155722
rect 182192 153610 182220 163254
rect 182836 163146 182864 163254
rect 182914 163200 182970 164400
rect 183742 163200 183798 164400
rect 184570 163200 184626 164400
rect 185398 163200 185454 164400
rect 186226 163200 186282 164400
rect 187054 163200 187110 164400
rect 187882 163200 187938 164400
rect 188802 163200 188858 164400
rect 189630 163200 189686 164400
rect 190458 163200 190514 164400
rect 191286 163200 191342 164400
rect 192114 163200 192170 164400
rect 192942 163200 192998 164400
rect 193770 163200 193826 164400
rect 194690 163200 194746 164400
rect 195518 163200 195574 164400
rect 196346 163200 196402 164400
rect 197174 163200 197230 164400
rect 198002 163200 198058 164400
rect 198830 163200 198886 164400
rect 199658 163200 199714 164400
rect 200578 163200 200634 164400
rect 201406 163200 201462 164400
rect 202234 163200 202290 164400
rect 202340 163254 202736 163282
rect 182928 163146 182956 163200
rect 182836 163118 182956 163146
rect 183100 159248 183152 159254
rect 183100 159190 183152 159196
rect 182272 157956 182324 157962
rect 182272 157898 182324 157904
rect 182088 153604 182140 153610
rect 182088 153546 182140 153552
rect 182180 153604 182232 153610
rect 182180 153546 182232 153552
rect 182100 150226 182128 153546
rect 181456 150198 181530 150226
rect 182100 150198 182174 150226
rect 182284 150210 182312 157898
rect 182732 152176 182784 152182
rect 182732 152118 182784 152124
rect 182744 150226 182772 152118
rect 183112 151842 183140 159190
rect 183756 158778 183784 163200
rect 184584 159866 184612 163200
rect 184572 159860 184624 159866
rect 184572 159802 184624 159808
rect 183744 158772 183796 158778
rect 183744 158714 183796 158720
rect 185412 157962 185440 163200
rect 185584 159044 185636 159050
rect 185584 158986 185636 158992
rect 185400 157956 185452 157962
rect 185400 157898 185452 157904
rect 185400 157684 185452 157690
rect 185400 157626 185452 157632
rect 184018 155816 184074 155825
rect 184018 155751 184074 155760
rect 183560 155168 183612 155174
rect 183560 155110 183612 155116
rect 183100 151836 183152 151842
rect 183100 151778 183152 151784
rect 180858 149940 180886 150198
rect 181502 149940 181530 150198
rect 182146 149940 182174 150198
rect 182272 150204 182324 150210
rect 182744 150198 182818 150226
rect 183572 150210 183600 155110
rect 184032 150226 184060 155751
rect 185124 154488 185176 154494
rect 185124 154430 185176 154436
rect 185136 153610 185164 154430
rect 185214 154320 185270 154329
rect 185214 154255 185216 154264
rect 185268 154255 185270 154264
rect 185308 154284 185360 154290
rect 185216 154226 185268 154232
rect 185308 154226 185360 154232
rect 185032 153604 185084 153610
rect 185032 153546 185084 153552
rect 185124 153604 185176 153610
rect 185124 153546 185176 153552
rect 185044 153490 185072 153546
rect 185320 153490 185348 154226
rect 185044 153462 185348 153490
rect 185308 152040 185360 152046
rect 185308 151982 185360 151988
rect 185320 150226 185348 151982
rect 185412 151814 185440 157626
rect 185596 152114 185624 158986
rect 186240 155786 186268 163200
rect 187068 159254 187096 163200
rect 187896 161474 187924 163200
rect 187896 161446 188016 161474
rect 187056 159248 187108 159254
rect 187056 159190 187108 159196
rect 186780 155916 186832 155922
rect 186780 155858 186832 155864
rect 186228 155780 186280 155786
rect 186228 155722 186280 155728
rect 186688 155168 186740 155174
rect 186688 155110 186740 155116
rect 186320 155100 186372 155106
rect 186504 155100 186556 155106
rect 186372 155060 186504 155088
rect 186320 155042 186372 155048
rect 186504 155042 186556 155048
rect 186228 155032 186280 155038
rect 186226 155000 186228 155009
rect 186596 155032 186648 155038
rect 186280 155000 186282 155009
rect 186594 155000 186596 155009
rect 186648 155000 186650 155009
rect 186226 154935 186282 154944
rect 186320 154964 186372 154970
rect 186594 154935 186650 154944
rect 186320 154906 186372 154912
rect 186332 154850 186360 154906
rect 186700 154850 186728 155110
rect 186332 154822 186728 154850
rect 185584 152108 185636 152114
rect 185584 152050 185636 152056
rect 185412 151786 185992 151814
rect 185964 150226 185992 151786
rect 186792 150226 186820 155858
rect 187238 154456 187294 154465
rect 187238 154391 187294 154400
rect 182272 150146 182324 150152
rect 182790 149940 182818 150198
rect 183422 150204 183474 150210
rect 183422 150146 183474 150152
rect 183560 150204 183612 150210
rect 184032 150198 184106 150226
rect 183560 150146 183612 150152
rect 183434 149940 183462 150146
rect 184078 149940 184106 150198
rect 184710 150204 184762 150210
rect 185320 150198 185394 150226
rect 185964 150198 186038 150226
rect 184710 150146 184762 150152
rect 184722 149940 184750 150146
rect 185366 149940 185394 150198
rect 186010 149940 186038 150198
rect 186654 150198 186820 150226
rect 186654 149940 186682 150198
rect 187252 150090 187280 154391
rect 187884 152924 187936 152930
rect 187884 152866 187936 152872
rect 187896 150090 187924 152866
rect 187988 152250 188016 161446
rect 188252 159928 188304 159934
rect 188252 159870 188304 159876
rect 188264 154970 188292 159870
rect 188816 157894 188844 163200
rect 188528 157888 188580 157894
rect 188528 157830 188580 157836
rect 188804 157888 188856 157894
rect 188804 157830 188856 157836
rect 188252 154964 188304 154970
rect 188252 154906 188304 154912
rect 188436 154420 188488 154426
rect 188436 154362 188488 154368
rect 188448 153610 188476 154362
rect 188344 153604 188396 153610
rect 188344 153546 188396 153552
rect 188436 153604 188488 153610
rect 188436 153546 188488 153552
rect 188356 153513 188384 153546
rect 188342 153504 188398 153513
rect 188342 153439 188398 153448
rect 187976 152244 188028 152250
rect 187976 152186 188028 152192
rect 188540 150226 188568 157830
rect 189170 155952 189226 155961
rect 189644 155922 189672 163200
rect 190472 157758 190500 163200
rect 191300 159934 191328 163200
rect 191748 159996 191800 160002
rect 191748 159938 191800 159944
rect 191288 159928 191340 159934
rect 191288 159870 191340 159876
rect 190644 157820 190696 157826
rect 190644 157762 190696 157768
rect 190460 157752 190512 157758
rect 190460 157694 190512 157700
rect 190656 157334 190684 157762
rect 191760 157334 191788 159938
rect 190656 157306 191144 157334
rect 189816 156392 189868 156398
rect 189816 156334 189868 156340
rect 189170 155887 189226 155896
rect 189632 155916 189684 155922
rect 188540 150198 188614 150226
rect 187252 150062 187326 150090
rect 187896 150062 187970 150090
rect 187298 149940 187326 150062
rect 187942 149940 187970 150062
rect 188586 149940 188614 150198
rect 189184 150090 189212 155887
rect 189632 155858 189684 155864
rect 189828 150090 189856 156334
rect 190460 151904 190512 151910
rect 190460 151846 190512 151852
rect 190472 150090 190500 151846
rect 191116 150226 191144 157306
rect 191668 157306 191788 157334
rect 191288 154488 191340 154494
rect 191288 154430 191340 154436
rect 191300 154358 191328 154430
rect 191472 154420 191524 154426
rect 191472 154362 191524 154368
rect 191288 154352 191340 154358
rect 191288 154294 191340 154300
rect 191380 154352 191432 154358
rect 191484 154329 191512 154362
rect 191380 154294 191432 154300
rect 191470 154320 191526 154329
rect 191392 153406 191420 154294
rect 191470 154255 191526 154264
rect 191380 153400 191432 153406
rect 191380 153342 191432 153348
rect 191668 152930 191696 157306
rect 192128 157214 192156 163200
rect 192668 158976 192720 158982
rect 192668 158918 192720 158924
rect 192116 157208 192168 157214
rect 192116 157150 192168 157156
rect 191748 155100 191800 155106
rect 191748 155042 191800 155048
rect 191656 152924 191708 152930
rect 191656 152866 191708 152872
rect 191116 150198 191190 150226
rect 189184 150062 189258 150090
rect 189828 150062 189902 150090
rect 190472 150062 190546 150090
rect 189230 149940 189258 150062
rect 189874 149940 189902 150062
rect 190518 149940 190546 150062
rect 191162 149940 191190 150198
rect 191760 150090 191788 155042
rect 192390 153504 192446 153513
rect 192390 153439 192446 153448
rect 192404 150090 192432 153439
rect 192680 152182 192708 158918
rect 192956 155174 192984 163200
rect 193588 159316 193640 159322
rect 193588 159258 193640 159264
rect 193680 159316 193732 159322
rect 193680 159258 193732 159264
rect 193600 159050 193628 159258
rect 193692 159186 193720 159258
rect 193784 159186 193812 163200
rect 193680 159180 193732 159186
rect 193680 159122 193732 159128
rect 193772 159180 193824 159186
rect 193772 159122 193824 159128
rect 193588 159044 193640 159050
rect 193588 158986 193640 158992
rect 194704 158846 194732 163200
rect 195152 158908 195204 158914
rect 195152 158850 195204 158856
rect 194508 158840 194560 158846
rect 194508 158782 194560 158788
rect 194692 158840 194744 158846
rect 194692 158782 194744 158788
rect 193220 157616 193272 157622
rect 193220 157558 193272 157564
rect 193232 157334 193260 157558
rect 193232 157306 193720 157334
rect 192944 155168 192996 155174
rect 192944 155110 192996 155116
rect 193036 152992 193088 152998
rect 193036 152934 193088 152940
rect 192668 152176 192720 152182
rect 192668 152118 192720 152124
rect 193048 150090 193076 152934
rect 193692 150226 193720 157306
rect 194324 155032 194376 155038
rect 194324 154974 194376 154980
rect 193692 150198 193766 150226
rect 191760 150062 191834 150090
rect 192404 150062 192478 150090
rect 193048 150062 193122 150090
rect 191806 149940 191834 150062
rect 192450 149940 192478 150062
rect 193094 149940 193122 150062
rect 193738 149940 193766 150198
rect 194336 150090 194364 154974
rect 194520 153406 194548 158782
rect 194968 155100 195020 155106
rect 194968 155042 195020 155048
rect 194508 153400 194560 153406
rect 194508 153342 194560 153348
rect 194980 150090 195008 155042
rect 195164 152046 195192 158850
rect 195532 157826 195560 163200
rect 195520 157820 195572 157826
rect 195520 157762 195572 157768
rect 196256 156324 196308 156330
rect 196256 156266 196308 156272
rect 195152 152040 195204 152046
rect 195152 151982 195204 151988
rect 195612 151836 195664 151842
rect 195612 151778 195664 151784
rect 195624 150090 195652 151778
rect 196268 150226 196296 156266
rect 196360 155106 196388 163200
rect 196992 159044 197044 159050
rect 196992 158986 197044 158992
rect 196348 155100 196400 155106
rect 196348 155042 196400 155048
rect 197004 153542 197032 158986
rect 197188 158982 197216 163200
rect 198016 160002 198044 163200
rect 198004 159996 198056 160002
rect 198004 159938 198056 159944
rect 197360 159316 197412 159322
rect 197360 159258 197412 159264
rect 197176 158976 197228 158982
rect 197176 158918 197228 158924
rect 197372 157622 197400 159258
rect 198738 158536 198794 158545
rect 198738 158471 198794 158480
rect 197360 157616 197412 157622
rect 197360 157558 197412 157564
rect 197544 153604 197596 153610
rect 197544 153546 197596 153552
rect 196900 153536 196952 153542
rect 196900 153478 196952 153484
rect 196992 153536 197044 153542
rect 196992 153478 197044 153484
rect 196912 150226 196940 153478
rect 197556 150226 197584 153546
rect 198188 153060 198240 153066
rect 198188 153002 198240 153008
rect 198200 150226 198228 153002
rect 198752 151814 198780 158471
rect 198844 156534 198872 163200
rect 198924 160064 198976 160070
rect 198924 160006 198976 160012
rect 198832 156528 198884 156534
rect 198832 156470 198884 156476
rect 198936 153542 198964 160006
rect 199672 155038 199700 163200
rect 200592 159050 200620 163200
rect 201420 159322 201448 163200
rect 202248 163146 202276 163200
rect 202340 163146 202368 163254
rect 202248 163118 202368 163146
rect 201408 159316 201460 159322
rect 201408 159258 201460 159264
rect 200580 159044 200632 159050
rect 200580 158986 200632 158992
rect 201408 158908 201460 158914
rect 201408 158850 201460 158856
rect 200304 156256 200356 156262
rect 200304 156198 200356 156204
rect 199660 155032 199712 155038
rect 199660 154974 199712 154980
rect 200120 154488 200172 154494
rect 200120 154430 200172 154436
rect 198924 153536 198976 153542
rect 198924 153478 198976 153484
rect 199476 153468 199528 153474
rect 199476 153410 199528 153416
rect 198752 151786 198872 151814
rect 198844 150226 198872 151786
rect 199488 150226 199516 153410
rect 200132 150226 200160 154430
rect 196268 150198 196342 150226
rect 196912 150198 196986 150226
rect 197556 150198 197630 150226
rect 198200 150198 198274 150226
rect 198844 150198 198918 150226
rect 199488 150198 199562 150226
rect 200132 150198 200206 150226
rect 200316 150210 200344 156198
rect 201420 153474 201448 158850
rect 202708 156466 202736 163254
rect 203062 163200 203118 164400
rect 203890 163200 203946 164400
rect 204718 163200 204774 164400
rect 204824 163254 205496 163282
rect 203076 160070 203104 163200
rect 203064 160064 203116 160070
rect 203064 160006 203116 160012
rect 203904 159186 203932 163200
rect 204732 159361 204760 163200
rect 204718 159352 204774 159361
rect 204718 159287 204774 159296
rect 203892 159180 203944 159186
rect 203892 159122 203944 159128
rect 203708 158840 203760 158846
rect 203708 158782 203760 158788
rect 203432 157548 203484 157554
rect 203432 157490 203484 157496
rect 202788 157276 202840 157282
rect 202788 157218 202840 157224
rect 202696 156460 202748 156466
rect 202696 156402 202748 156408
rect 202800 156330 202828 157218
rect 202788 156324 202840 156330
rect 202788 156266 202840 156272
rect 202696 154420 202748 154426
rect 202696 154362 202748 154368
rect 202052 154352 202104 154358
rect 202052 154294 202104 154300
rect 201408 153468 201460 153474
rect 201408 153410 201460 153416
rect 200764 152108 200816 152114
rect 200764 152050 200816 152056
rect 200776 150226 200804 152050
rect 202064 150226 202092 154294
rect 202708 150226 202736 154362
rect 203340 151972 203392 151978
rect 203340 151914 203392 151920
rect 203352 150226 203380 151914
rect 203444 151814 203472 157490
rect 203720 152998 203748 158782
rect 203892 156188 203944 156194
rect 203892 156130 203944 156136
rect 203904 155417 203932 156130
rect 204352 155848 204404 155854
rect 204352 155790 204404 155796
rect 203890 155408 203946 155417
rect 203890 155343 203946 155352
rect 203708 152992 203760 152998
rect 203708 152934 203760 152940
rect 204364 151814 204392 155790
rect 204824 154358 204852 163254
rect 205468 163146 205496 163254
rect 205546 163200 205602 164400
rect 206466 163200 206522 164400
rect 207294 163200 207350 164400
rect 208122 163200 208178 164400
rect 208412 163254 208900 163282
rect 205560 163146 205588 163200
rect 205468 163118 205588 163146
rect 204904 158772 204956 158778
rect 204904 158714 204956 158720
rect 204916 157554 204944 158714
rect 204904 157548 204956 157554
rect 204904 157490 204956 157496
rect 204904 157344 204956 157350
rect 204904 157286 204956 157292
rect 205270 157312 205326 157321
rect 204916 156534 204944 157286
rect 204996 157276 205048 157282
rect 204996 157218 205048 157224
rect 205088 157276 205140 157282
rect 205270 157247 205326 157256
rect 205088 157218 205140 157224
rect 205008 156534 205036 157218
rect 204904 156528 204956 156534
rect 204904 156470 204956 156476
rect 204996 156528 205048 156534
rect 204996 156470 205048 156476
rect 205100 156466 205128 157218
rect 205088 156460 205140 156466
rect 205088 156402 205140 156408
rect 204812 154352 204864 154358
rect 204812 154294 204864 154300
rect 203444 151786 204024 151814
rect 204364 151786 204668 151814
rect 203996 150226 204024 151786
rect 204640 150226 204668 151786
rect 205284 150226 205312 157247
rect 205916 156256 205968 156262
rect 205744 156204 205916 156210
rect 205744 156198 205968 156204
rect 205744 156182 205956 156198
rect 205744 156126 205772 156182
rect 205732 156120 205784 156126
rect 205732 156062 205784 156068
rect 206480 155854 206508 163200
rect 206928 159180 206980 159186
rect 206928 159122 206980 159128
rect 206940 158846 206968 159122
rect 207308 158914 207336 163200
rect 208136 159322 208164 163200
rect 207388 159316 207440 159322
rect 207388 159258 207440 159264
rect 208124 159316 208176 159322
rect 208124 159258 208176 159264
rect 207400 159118 207428 159258
rect 207388 159112 207440 159118
rect 207388 159054 207440 159060
rect 207296 158908 207348 158914
rect 207296 158850 207348 158856
rect 206928 158840 206980 158846
rect 206928 158782 206980 158788
rect 206560 157480 206612 157486
rect 206560 157422 206612 157428
rect 206468 155848 206520 155854
rect 206468 155790 206520 155796
rect 205916 153196 205968 153202
rect 205916 153138 205968 153144
rect 194336 150062 194410 150090
rect 194980 150062 195054 150090
rect 195624 150062 195698 150090
rect 194382 149940 194410 150062
rect 195026 149940 195054 150062
rect 195670 149940 195698 150062
rect 196314 149940 196342 150198
rect 196958 149940 196986 150198
rect 197602 149940 197630 150198
rect 198246 149940 198274 150198
rect 198890 149940 198918 150198
rect 199534 149940 199562 150198
rect 200178 149940 200206 150198
rect 200304 150204 200356 150210
rect 200776 150198 200850 150226
rect 200304 150146 200356 150152
rect 200822 149940 200850 150198
rect 201454 150204 201506 150210
rect 202064 150198 202138 150226
rect 202708 150198 202782 150226
rect 203352 150198 203426 150226
rect 203996 150198 204070 150226
rect 204640 150198 204714 150226
rect 205284 150198 205358 150226
rect 201454 150146 201506 150152
rect 201466 149940 201494 150146
rect 202110 149940 202138 150198
rect 202754 149940 202782 150198
rect 203398 149940 203426 150198
rect 204042 149940 204070 150198
rect 204686 149940 204714 150198
rect 205330 149940 205358 150198
rect 205928 150090 205956 153138
rect 206572 150226 206600 157422
rect 208412 154426 208440 163254
rect 208872 163146 208900 163254
rect 208950 163200 209006 164400
rect 209778 163200 209834 164400
rect 210606 163200 210662 164400
rect 211434 163200 211490 164400
rect 211540 163254 212304 163282
rect 208964 163146 208992 163200
rect 208872 163118 208992 163146
rect 209792 156670 209820 163200
rect 210620 158778 210648 163200
rect 211448 160070 211476 163200
rect 211068 160064 211120 160070
rect 211068 160006 211120 160012
rect 211436 160064 211488 160070
rect 211436 160006 211488 160012
rect 210608 158772 210660 158778
rect 210608 158714 210660 158720
rect 210516 156936 210568 156942
rect 210516 156878 210568 156884
rect 210608 156936 210660 156942
rect 210608 156878 210660 156884
rect 209688 156664 209740 156670
rect 209686 156632 209688 156641
rect 209780 156664 209832 156670
rect 209740 156632 209742 156641
rect 209780 156606 209832 156612
rect 209686 156567 209742 156576
rect 210528 156534 210556 156878
rect 210424 156528 210476 156534
rect 210424 156470 210476 156476
rect 210516 156528 210568 156534
rect 210516 156470 210568 156476
rect 210436 156330 210464 156470
rect 210424 156324 210476 156330
rect 210424 156266 210476 156272
rect 210620 156262 210648 156878
rect 210700 156664 210752 156670
rect 210792 156664 210844 156670
rect 210700 156606 210752 156612
rect 210790 156632 210792 156641
rect 210844 156632 210846 156641
rect 210712 156466 210740 156606
rect 210790 156567 210846 156576
rect 210700 156460 210752 156466
rect 210700 156402 210752 156408
rect 210608 156256 210660 156262
rect 210608 156198 210660 156204
rect 211080 156126 211108 160006
rect 211068 156120 211120 156126
rect 211068 156062 211120 156068
rect 209134 155408 209190 155417
rect 209134 155343 209190 155352
rect 208400 154420 208452 154426
rect 208400 154362 208452 154368
rect 207204 153332 207256 153338
rect 207204 153274 207256 153280
rect 206572 150198 206646 150226
rect 205928 150062 206002 150090
rect 205974 149940 206002 150062
rect 206618 149940 206646 150198
rect 207216 150090 207244 153274
rect 207848 153264 207900 153270
rect 207848 153206 207900 153212
rect 207860 150090 207888 153206
rect 208492 152924 208544 152930
rect 208492 152866 208544 152872
rect 208504 150090 208532 152866
rect 209148 150090 209176 155343
rect 209780 153876 209832 153882
rect 209780 153818 209832 153824
rect 209792 150090 209820 153818
rect 211540 153785 211568 163254
rect 212276 163146 212304 163254
rect 212354 163200 212410 164400
rect 213182 163200 213238 164400
rect 214010 163200 214066 164400
rect 214838 163200 214894 164400
rect 215312 163254 215616 163282
rect 212368 163146 212396 163200
rect 212276 163118 212396 163146
rect 212448 159316 212500 159322
rect 212448 159258 212500 159264
rect 211620 156188 211672 156194
rect 211620 156130 211672 156136
rect 211526 153776 211582 153785
rect 210424 153740 210476 153746
rect 211526 153711 211582 153720
rect 210424 153682 210476 153688
rect 210436 150090 210464 153682
rect 211068 152380 211120 152386
rect 211068 152322 211120 152328
rect 211080 150090 211108 152322
rect 211632 150090 211660 156130
rect 212264 154896 212316 154902
rect 212264 154838 212316 154844
rect 212276 150090 212304 154838
rect 212460 152930 212488 159258
rect 212644 159174 212856 159202
rect 212644 158982 212672 159174
rect 212828 159118 212856 159174
rect 212724 159112 212776 159118
rect 212724 159054 212776 159060
rect 212816 159112 212868 159118
rect 212816 159054 212868 159060
rect 212632 158976 212684 158982
rect 212632 158918 212684 158924
rect 212448 152924 212500 152930
rect 212448 152866 212500 152872
rect 212736 151978 212764 159054
rect 213196 156262 213224 163200
rect 214024 159322 214052 163200
rect 214012 159316 214064 159322
rect 214012 159258 214064 159264
rect 214852 158846 214880 163200
rect 213828 158840 213880 158846
rect 213828 158782 213880 158788
rect 214840 158840 214892 158846
rect 214840 158782 214892 158788
rect 213184 156256 213236 156262
rect 213184 156198 213236 156204
rect 212908 153808 212960 153814
rect 212908 153750 212960 153756
rect 212724 151972 212776 151978
rect 212724 151914 212776 151920
rect 212920 150090 212948 153750
rect 213840 152182 213868 158782
rect 214104 156800 214156 156806
rect 214156 156748 214328 156754
rect 214104 156742 214328 156748
rect 214116 156726 214328 156742
rect 214300 156670 214328 156726
rect 214196 156664 214248 156670
rect 214196 156606 214248 156612
rect 214288 156664 214340 156670
rect 214288 156606 214340 156612
rect 213552 152176 213604 152182
rect 213552 152118 213604 152124
rect 213828 152176 213880 152182
rect 213828 152118 213880 152124
rect 213564 150090 213592 152118
rect 214208 150090 214236 156606
rect 214840 154828 214892 154834
rect 214840 154770 214892 154776
rect 214852 150090 214880 154770
rect 215312 153882 215340 163254
rect 215588 163146 215616 163254
rect 215666 163200 215722 164400
rect 216494 163200 216550 164400
rect 217322 163200 217378 164400
rect 218242 163200 218298 164400
rect 218348 163254 219020 163282
rect 215680 163146 215708 163200
rect 215588 163118 215708 163146
rect 215392 158772 215444 158778
rect 215392 158714 215444 158720
rect 215300 153876 215352 153882
rect 215300 153818 215352 153824
rect 215404 153066 215432 158714
rect 216508 156670 216536 163200
rect 216772 159248 216824 159254
rect 216772 159190 216824 159196
rect 216404 156664 216456 156670
rect 216404 156606 216456 156612
rect 216496 156664 216548 156670
rect 216496 156606 216548 156612
rect 216416 156482 216444 156606
rect 216416 156454 216720 156482
rect 215484 153672 215536 153678
rect 215484 153614 215536 153620
rect 215392 153060 215444 153066
rect 215392 153002 215444 153008
rect 215496 150226 215524 153614
rect 216128 152652 216180 152658
rect 216128 152594 216180 152600
rect 216140 150226 216168 152594
rect 216692 151814 216720 156454
rect 216784 154834 216812 159190
rect 217336 158982 217364 163200
rect 218256 159254 218284 163200
rect 218244 159248 218296 159254
rect 218244 159190 218296 159196
rect 217324 158976 217376 158982
rect 217324 158918 217376 158924
rect 217416 155236 217468 155242
rect 217416 155178 217468 155184
rect 216772 154828 216824 154834
rect 216772 154770 216824 154776
rect 216692 151786 216812 151814
rect 216784 150226 216812 151786
rect 217428 150226 217456 155178
rect 218348 154494 218376 163254
rect 218992 163146 219020 163254
rect 219070 163200 219126 164400
rect 219898 163200 219954 164400
rect 220726 163200 220782 164400
rect 221554 163200 221610 164400
rect 222382 163200 222438 164400
rect 223210 163200 223266 164400
rect 224130 163200 224186 164400
rect 224958 163200 225014 164400
rect 225064 163254 225736 163282
rect 219084 163146 219112 163200
rect 218992 163118 219112 163146
rect 219348 158024 219400 158030
rect 219348 157966 219400 157972
rect 218336 154488 218388 154494
rect 218336 154430 218388 154436
rect 218060 153944 218112 153950
rect 218060 153886 218112 153892
rect 218072 150226 218100 153886
rect 218704 152040 218756 152046
rect 218704 151982 218756 151988
rect 218716 150226 218744 151982
rect 219360 150226 219388 157966
rect 219912 156806 219940 163200
rect 220740 159186 220768 163200
rect 220636 159180 220688 159186
rect 220636 159122 220688 159128
rect 220728 159180 220780 159186
rect 220728 159122 220780 159128
rect 220452 158976 220504 158982
rect 220452 158918 220504 158924
rect 219900 156800 219952 156806
rect 219900 156742 219952 156748
rect 219992 156732 220044 156738
rect 219992 156674 220044 156680
rect 219532 156324 219584 156330
rect 219532 156266 219584 156272
rect 215496 150198 215570 150226
rect 216140 150198 216214 150226
rect 216784 150198 216858 150226
rect 217428 150198 217502 150226
rect 218072 150198 218146 150226
rect 218716 150198 218790 150226
rect 219360 150198 219434 150226
rect 219544 150210 219572 156266
rect 220004 150226 220032 156674
rect 220464 152658 220492 158918
rect 220648 156194 220676 159122
rect 221568 158778 221596 163200
rect 222108 159112 222160 159118
rect 222108 159054 222160 159060
rect 221740 158840 221792 158846
rect 221740 158782 221792 158788
rect 221556 158772 221608 158778
rect 221556 158714 221608 158720
rect 221372 156528 221424 156534
rect 221372 156470 221424 156476
rect 220636 156188 220688 156194
rect 220636 156130 220688 156136
rect 220452 152652 220504 152658
rect 220452 152594 220504 152600
rect 221280 152584 221332 152590
rect 221280 152526 221332 152532
rect 221292 150226 221320 152526
rect 221384 151814 221412 156470
rect 221752 152386 221780 158782
rect 222120 156330 222148 159054
rect 222292 156936 222344 156942
rect 222292 156878 222344 156884
rect 222108 156324 222160 156330
rect 222108 156266 222160 156272
rect 221740 152380 221792 152386
rect 221740 152322 221792 152328
rect 221384 151786 221964 151814
rect 221936 150226 221964 151786
rect 207216 150062 207290 150090
rect 207860 150062 207934 150090
rect 208504 150062 208578 150090
rect 209148 150062 209222 150090
rect 209792 150062 209866 150090
rect 210436 150062 210510 150090
rect 211080 150062 211154 150090
rect 211632 150062 211706 150090
rect 212276 150062 212350 150090
rect 212920 150062 212994 150090
rect 213564 150062 213638 150090
rect 214208 150062 214282 150090
rect 214852 150062 214926 150090
rect 207262 149940 207290 150062
rect 207906 149940 207934 150062
rect 208550 149940 208578 150062
rect 209194 149940 209222 150062
rect 209838 149940 209866 150062
rect 210482 149940 210510 150062
rect 211126 149940 211154 150062
rect 211678 149940 211706 150062
rect 212322 149940 212350 150062
rect 212966 149940 212994 150062
rect 213610 149940 213638 150062
rect 214254 149940 214282 150062
rect 214898 149940 214926 150062
rect 215542 149940 215570 150198
rect 216186 149940 216214 150198
rect 216830 149940 216858 150198
rect 217474 149940 217502 150198
rect 218118 149940 218146 150198
rect 218762 149940 218790 150198
rect 219406 149940 219434 150198
rect 219532 150204 219584 150210
rect 220004 150198 220078 150226
rect 219532 150146 219584 150152
rect 220050 149940 220078 150198
rect 220682 150204 220734 150210
rect 221292 150198 221366 150226
rect 221936 150198 222010 150226
rect 222304 150210 222332 156878
rect 222396 153814 222424 163200
rect 223224 156738 223252 163200
rect 223672 159384 223724 159390
rect 223672 159326 223724 159332
rect 223212 156732 223264 156738
rect 223212 156674 223264 156680
rect 223580 156528 223632 156534
rect 223580 156470 223632 156476
rect 223592 156262 223620 156470
rect 223580 156256 223632 156262
rect 223580 156198 223632 156204
rect 222568 156052 222620 156058
rect 222568 155994 222620 156000
rect 222384 153808 222436 153814
rect 222384 153750 222436 153756
rect 222580 150226 222608 155994
rect 223684 151814 223712 159326
rect 224144 159118 224172 163200
rect 224972 159390 225000 163200
rect 224960 159384 225012 159390
rect 224960 159326 225012 159332
rect 224132 159112 224184 159118
rect 224132 159054 224184 159060
rect 223856 158772 223908 158778
rect 223856 158714 223908 158720
rect 223868 153202 223896 158714
rect 224132 157004 224184 157010
rect 224132 156946 224184 156952
rect 223856 153196 223908 153202
rect 223856 153138 223908 153144
rect 224144 151814 224172 156946
rect 225064 153950 225092 163254
rect 225708 163146 225736 163254
rect 225786 163200 225842 164400
rect 226614 163200 226670 164400
rect 227442 163200 227498 164400
rect 227916 163254 228220 163282
rect 225800 163146 225828 163200
rect 225708 163118 225828 163146
rect 225236 159520 225288 159526
rect 225236 159462 225288 159468
rect 225144 156868 225196 156874
rect 225144 156810 225196 156816
rect 225052 153944 225104 153950
rect 225052 153886 225104 153892
rect 223684 151786 223896 151814
rect 224144 151786 224540 151814
rect 223868 150226 223896 151786
rect 224512 150226 224540 151786
rect 225156 150226 225184 156810
rect 225248 152590 225276 159462
rect 226628 156942 226656 163200
rect 227076 157412 227128 157418
rect 227076 157354 227128 157360
rect 226616 156936 226668 156942
rect 226616 156878 226668 156884
rect 225788 154556 225840 154562
rect 225788 154498 225840 154504
rect 225236 152584 225288 152590
rect 225236 152526 225288 152532
rect 225800 150226 225828 154498
rect 226432 152516 226484 152522
rect 226432 152458 226484 152464
rect 226444 150226 226472 152458
rect 227088 150226 227116 157354
rect 227456 152425 227484 163200
rect 227720 159044 227772 159050
rect 227720 158986 227772 158992
rect 227732 156194 227760 158986
rect 227720 156188 227772 156194
rect 227720 156130 227772 156136
rect 227812 155304 227864 155310
rect 227812 155246 227864 155252
rect 227442 152416 227498 152425
rect 227442 152351 227498 152360
rect 227824 150226 227852 155246
rect 227916 152522 227944 163254
rect 228192 163146 228220 163254
rect 228270 163200 228326 164400
rect 229098 163200 229154 164400
rect 230018 163200 230074 164400
rect 230846 163200 230902 164400
rect 231674 163200 231730 164400
rect 231872 163254 232452 163282
rect 228284 163146 228312 163200
rect 228192 163118 228312 163146
rect 228364 156596 228416 156602
rect 228364 156538 228416 156544
rect 227904 152516 227956 152522
rect 227904 152458 227956 152464
rect 220682 150146 220734 150152
rect 220694 149940 220722 150146
rect 221338 149940 221366 150198
rect 221982 149940 222010 150198
rect 222292 150204 222344 150210
rect 222580 150198 222654 150226
rect 222292 150146 222344 150152
rect 222626 149940 222654 150198
rect 223258 150204 223310 150210
rect 223868 150198 223942 150226
rect 224512 150198 224586 150226
rect 225156 150198 225230 150226
rect 225800 150198 225874 150226
rect 226444 150198 226518 150226
rect 227088 150198 227162 150226
rect 223258 150146 223310 150152
rect 223270 149940 223298 150146
rect 223914 149940 223942 150198
rect 224558 149940 224586 150198
rect 225202 149940 225230 150198
rect 225846 149940 225874 150198
rect 226490 149940 226518 150198
rect 227134 149940 227162 150198
rect 227778 150198 227852 150226
rect 228376 150226 228404 156538
rect 229112 153746 229140 163200
rect 230032 156874 230060 163200
rect 230860 159050 230888 163200
rect 231688 159526 231716 163200
rect 231676 159520 231728 159526
rect 231676 159462 231728 159468
rect 230848 159044 230900 159050
rect 230848 158986 230900 158992
rect 231768 158908 231820 158914
rect 231768 158850 231820 158856
rect 230020 156868 230072 156874
rect 230020 156810 230072 156816
rect 230940 156392 230992 156398
rect 230940 156334 230992 156340
rect 229652 155984 229704 155990
rect 229652 155926 229704 155932
rect 229192 155372 229244 155378
rect 229192 155314 229244 155320
rect 229100 153740 229152 153746
rect 229100 153682 229152 153688
rect 229008 152584 229060 152590
rect 229008 152526 229060 152532
rect 229020 150226 229048 152526
rect 228376 150198 228450 150226
rect 229020 150198 229094 150226
rect 229204 150210 229232 155314
rect 229664 150226 229692 155926
rect 230952 150226 230980 156334
rect 231780 154902 231808 158850
rect 231768 154896 231820 154902
rect 231768 154838 231820 154844
rect 231872 154562 231900 163254
rect 232424 163146 232452 163254
rect 232502 163200 232558 164400
rect 233330 163200 233386 164400
rect 234158 163200 234214 164400
rect 234986 163200 235042 164400
rect 235092 163254 235856 163282
rect 232516 163146 232544 163200
rect 232424 163118 232544 163146
rect 233344 158098 233372 163200
rect 234068 159452 234120 159458
rect 234068 159394 234120 159400
rect 231952 158092 232004 158098
rect 231952 158034 232004 158040
rect 233332 158092 233384 158098
rect 233332 158034 233384 158040
rect 231860 154556 231912 154562
rect 231860 154498 231912 154504
rect 231584 152788 231636 152794
rect 231584 152730 231636 152736
rect 231596 150226 231624 152730
rect 231964 151814 231992 158034
rect 232872 155440 232924 155446
rect 232872 155382 232924 155388
rect 231964 151786 232268 151814
rect 232240 150226 232268 151786
rect 232884 150226 232912 155382
rect 233516 154012 233568 154018
rect 233516 153954 233568 153960
rect 233528 150226 233556 153954
rect 234080 151814 234108 159394
rect 234172 152590 234200 163200
rect 235000 159458 235028 163200
rect 234988 159452 235040 159458
rect 234988 159394 235040 159400
rect 234804 157072 234856 157078
rect 234804 157014 234856 157020
rect 234160 152584 234212 152590
rect 234160 152526 234212 152532
rect 234080 151786 234200 151814
rect 234172 150226 234200 151786
rect 234816 150226 234844 157014
rect 235092 154018 235120 163254
rect 235828 163146 235856 163254
rect 235906 163200 235962 164400
rect 236734 163200 236790 164400
rect 237562 163200 237618 164400
rect 238390 163200 238446 164400
rect 238864 163254 239168 163282
rect 235920 163146 235948 163200
rect 235828 163118 235948 163146
rect 236184 157684 236236 157690
rect 236184 157626 236236 157632
rect 235448 154080 235500 154086
rect 235448 154022 235500 154028
rect 235080 154012 235132 154018
rect 235080 153954 235132 153960
rect 235460 150226 235488 154022
rect 236196 150226 236224 157626
rect 236748 155242 236776 163200
rect 237576 158982 237604 163200
rect 237564 158976 237616 158982
rect 237564 158918 237616 158924
rect 238404 158914 238432 163200
rect 238392 158908 238444 158914
rect 238392 158850 238444 158856
rect 237380 158160 237432 158166
rect 237380 158102 237432 158108
rect 236736 155236 236788 155242
rect 236736 155178 236788 155184
rect 236736 152720 236788 152726
rect 236736 152662 236788 152668
rect 227778 149940 227806 150198
rect 228422 149940 228450 150198
rect 229066 149940 229094 150198
rect 229192 150204 229244 150210
rect 229664 150198 229738 150226
rect 229192 150146 229244 150152
rect 229710 149940 229738 150198
rect 230342 150204 230394 150210
rect 230952 150198 231026 150226
rect 231596 150198 231670 150226
rect 232240 150198 232314 150226
rect 232884 150198 232958 150226
rect 233528 150198 233602 150226
rect 234172 150198 234246 150226
rect 234816 150198 234890 150226
rect 235460 150198 235534 150226
rect 230342 150146 230394 150152
rect 230354 149940 230382 150146
rect 230998 149940 231026 150198
rect 231642 149940 231670 150198
rect 232286 149940 232314 150198
rect 232930 149940 232958 150198
rect 233574 149940 233602 150198
rect 234218 149940 234246 150198
rect 234862 149940 234890 150198
rect 235506 149940 235534 150198
rect 236150 150198 236224 150226
rect 236748 150226 236776 152662
rect 237392 150226 237420 158102
rect 238024 154760 238076 154766
rect 238024 154702 238076 154708
rect 238036 150226 238064 154702
rect 238864 153678 238892 163254
rect 239140 163146 239168 163254
rect 239218 163200 239274 164400
rect 240046 163200 240102 164400
rect 240874 163200 240930 164400
rect 241794 163200 241850 164400
rect 241900 163254 242572 163282
rect 239232 163146 239260 163200
rect 239140 163118 239260 163146
rect 239312 159588 239364 159594
rect 239312 159530 239364 159536
rect 238944 158228 238996 158234
rect 238944 158170 238996 158176
rect 238852 153672 238904 153678
rect 238852 153614 238904 153620
rect 238668 153400 238720 153406
rect 238668 153342 238720 153348
rect 238680 150226 238708 153342
rect 236748 150198 236822 150226
rect 237392 150198 237466 150226
rect 238036 150198 238110 150226
rect 238680 150198 238754 150226
rect 238956 150210 238984 158170
rect 239324 150226 239352 159530
rect 240060 158030 240088 163200
rect 240324 159656 240376 159662
rect 240324 159598 240376 159604
rect 240048 158024 240100 158030
rect 240048 157966 240100 157972
rect 240140 154624 240192 154630
rect 240140 154566 240192 154572
rect 240152 151814 240180 154566
rect 240336 152794 240364 159598
rect 240888 158778 240916 163200
rect 241808 159662 241836 163200
rect 241796 159656 241848 159662
rect 241796 159598 241848 159604
rect 240876 158772 240928 158778
rect 240876 158714 240928 158720
rect 240692 154964 240744 154970
rect 240692 154906 240744 154912
rect 240324 152788 240376 152794
rect 240324 152730 240376 152736
rect 240704 151814 240732 154906
rect 241900 154086 241928 163254
rect 242544 163146 242572 163254
rect 242622 163200 242678 164400
rect 243450 163200 243506 164400
rect 244278 163200 244334 164400
rect 244384 163254 245056 163282
rect 242636 163146 242664 163200
rect 242544 163118 242664 163146
rect 242808 158908 242860 158914
rect 242808 158850 242860 158856
rect 242072 158296 242124 158302
rect 242072 158238 242124 158244
rect 241888 154080 241940 154086
rect 241888 154022 241940 154028
rect 241888 152788 241940 152794
rect 241888 152730 241940 152736
rect 240152 151786 240640 151814
rect 240704 151786 241284 151814
rect 240612 150226 240640 151786
rect 241256 150226 241284 151786
rect 241900 150226 241928 152730
rect 242084 151814 242112 158238
rect 242820 152046 242848 158850
rect 243360 158772 243412 158778
rect 243360 158714 243412 158720
rect 243084 154692 243136 154698
rect 243084 154634 243136 154640
rect 242808 152040 242860 152046
rect 242808 151982 242860 151988
rect 242084 151786 242480 151814
rect 242452 150226 242480 151786
rect 243096 150226 243124 154634
rect 243372 151978 243400 158714
rect 243464 155310 243492 163200
rect 244292 158914 244320 163200
rect 244280 158908 244332 158914
rect 244280 158850 244332 158856
rect 243452 155304 243504 155310
rect 243452 155246 243504 155252
rect 243728 153604 243780 153610
rect 243728 153546 243780 153552
rect 243360 151972 243412 151978
rect 243360 151914 243412 151920
rect 243740 150226 243768 153546
rect 244384 152794 244412 163254
rect 245028 163146 245056 163254
rect 245106 163200 245162 164400
rect 245934 163200 245990 164400
rect 246762 163200 246818 164400
rect 247052 163254 247632 163282
rect 245120 163146 245148 163200
rect 245028 163118 245148 163146
rect 245016 158364 245068 158370
rect 245016 158306 245068 158312
rect 244372 152788 244424 152794
rect 244372 152730 244424 152736
rect 244372 152448 244424 152454
rect 244372 152390 244424 152396
rect 244384 150226 244412 152390
rect 245028 150226 245056 158306
rect 245844 157140 245896 157146
rect 245844 157082 245896 157088
rect 245660 154148 245712 154154
rect 245660 154090 245712 154096
rect 245672 150226 245700 154090
rect 245856 151814 245884 157082
rect 245948 153610 245976 163200
rect 246776 158166 246804 163200
rect 246948 159724 247000 159730
rect 246948 159666 247000 159672
rect 246764 158160 246816 158166
rect 246764 158102 246816 158108
rect 245936 153604 245988 153610
rect 245936 153546 245988 153552
rect 245856 151786 246344 151814
rect 246316 150226 246344 151786
rect 246960 150226 246988 159666
rect 247052 152726 247080 163254
rect 247604 163146 247632 163254
rect 247682 163200 247738 164400
rect 248510 163200 248566 164400
rect 248616 163254 249288 163282
rect 247696 163146 247724 163200
rect 247604 163118 247724 163146
rect 248524 159730 248552 163200
rect 248512 159724 248564 159730
rect 248512 159666 248564 159672
rect 247132 158432 247184 158438
rect 247132 158374 247184 158380
rect 247040 152720 247092 152726
rect 247040 152662 247092 152668
rect 247144 151814 247172 158374
rect 248236 155508 248288 155514
rect 248236 155450 248288 155456
rect 247144 151786 247632 151814
rect 247604 150226 247632 151786
rect 248248 150226 248276 155450
rect 248616 154154 248644 163254
rect 249260 163146 249288 163254
rect 249338 163200 249394 164400
rect 250166 163200 250222 164400
rect 250994 163200 251050 164400
rect 251192 163254 251772 163282
rect 249352 163146 249380 163200
rect 249260 163118 249380 163146
rect 250076 158636 250128 158642
rect 250076 158578 250128 158584
rect 248604 154148 248656 154154
rect 248604 154090 248656 154096
rect 248880 153536 248932 153542
rect 248880 153478 248932 153484
rect 248892 150226 248920 153478
rect 249524 152312 249576 152318
rect 249524 152254 249576 152260
rect 249536 150226 249564 152254
rect 250088 151814 250116 158578
rect 250180 155378 250208 163200
rect 251008 159594 251036 163200
rect 250996 159588 251048 159594
rect 250996 159530 251048 159536
rect 250168 155372 250220 155378
rect 250168 155314 250220 155320
rect 250812 154216 250864 154222
rect 250812 154158 250864 154164
rect 250088 151786 250208 151814
rect 250180 150226 250208 151786
rect 250824 150226 250852 154158
rect 251192 152454 251220 163254
rect 251744 163146 251772 163254
rect 251822 163200 251878 164400
rect 252650 163200 252706 164400
rect 253570 163200 253626 164400
rect 254398 163200 254454 164400
rect 255226 163200 255282 164400
rect 255332 163254 256004 163282
rect 251836 163146 251864 163200
rect 251744 163118 251864 163146
rect 251456 157616 251508 157622
rect 251456 157558 251508 157564
rect 251180 152448 251232 152454
rect 251180 152390 251232 152396
rect 251468 150226 251496 157558
rect 252664 153542 252692 163200
rect 252744 158568 252796 158574
rect 252744 158510 252796 158516
rect 252652 153536 252704 153542
rect 252652 153478 252704 153484
rect 252100 152856 252152 152862
rect 252100 152798 252152 152804
rect 252112 150226 252140 152798
rect 252756 150226 252784 158510
rect 253388 155712 253440 155718
rect 253388 155654 253440 155660
rect 253400 150226 253428 155654
rect 253584 155446 253612 163200
rect 253940 159792 253992 159798
rect 253940 159734 253992 159740
rect 253572 155440 253624 155446
rect 253572 155382 253624 155388
rect 236150 149940 236178 150198
rect 236794 149940 236822 150198
rect 237438 149940 237466 150198
rect 238082 149940 238110 150198
rect 238726 149940 238754 150198
rect 238944 150204 238996 150210
rect 239324 150198 239398 150226
rect 238944 150146 238996 150152
rect 239370 149940 239398 150198
rect 240002 150204 240054 150210
rect 240612 150198 240686 150226
rect 241256 150198 241330 150226
rect 241900 150198 241974 150226
rect 242452 150198 242526 150226
rect 243096 150198 243170 150226
rect 243740 150198 243814 150226
rect 244384 150198 244458 150226
rect 245028 150198 245102 150226
rect 245672 150198 245746 150226
rect 246316 150198 246390 150226
rect 246960 150198 247034 150226
rect 247604 150198 247678 150226
rect 248248 150198 248322 150226
rect 248892 150198 248966 150226
rect 249536 150198 249610 150226
rect 250180 150198 250254 150226
rect 250824 150198 250898 150226
rect 251468 150198 251542 150226
rect 252112 150198 252186 150226
rect 252756 150198 252830 150226
rect 253400 150198 253474 150226
rect 253952 150210 253980 159734
rect 254412 158778 254440 163200
rect 255240 159798 255268 163200
rect 255228 159792 255280 159798
rect 255228 159734 255280 159740
rect 254400 158772 254452 158778
rect 254400 158714 254452 158720
rect 254032 155644 254084 155650
rect 254032 155586 254084 155592
rect 254044 150226 254072 155586
rect 255332 154222 255360 163254
rect 255976 163146 256004 163254
rect 256054 163200 256110 164400
rect 256882 163200 256938 164400
rect 257710 163200 257766 164400
rect 258538 163200 258594 164400
rect 259458 163200 259514 164400
rect 260286 163200 260342 164400
rect 261114 163200 261170 164400
rect 261942 163200 261998 164400
rect 262232 163254 262720 163282
rect 256068 163146 256096 163200
rect 255976 163118 256096 163146
rect 255504 158772 255556 158778
rect 255504 158714 255556 158720
rect 255412 158500 255464 158506
rect 255412 158442 255464 158448
rect 255320 154216 255372 154222
rect 255320 154158 255372 154164
rect 255424 150226 255452 158442
rect 255516 152318 255544 158714
rect 256792 158704 256844 158710
rect 256792 158646 256844 158652
rect 255872 155576 255924 155582
rect 255872 155518 255924 155524
rect 255504 152312 255556 152318
rect 255504 152254 255556 152260
rect 255884 151814 255912 155518
rect 256608 153468 256660 153474
rect 256608 153410 256660 153416
rect 255884 151786 256004 151814
rect 240002 150146 240054 150152
rect 240014 149940 240042 150146
rect 240658 149940 240686 150198
rect 241302 149940 241330 150198
rect 241946 149940 241974 150198
rect 242498 149940 242526 150198
rect 243142 149940 243170 150198
rect 243786 149940 243814 150198
rect 244430 149940 244458 150198
rect 245074 149940 245102 150198
rect 245718 149940 245746 150198
rect 246362 149940 246390 150198
rect 247006 149940 247034 150198
rect 247650 149940 247678 150198
rect 248294 149940 248322 150198
rect 248938 149940 248966 150198
rect 249582 149940 249610 150198
rect 250226 149940 250254 150198
rect 250870 149940 250898 150198
rect 251514 149940 251542 150198
rect 252158 149940 252186 150198
rect 252802 149940 252830 150198
rect 253446 149940 253474 150198
rect 253940 150204 253992 150210
rect 254044 150198 254118 150226
rect 253940 150146 253992 150152
rect 254090 149940 254118 150198
rect 254722 150204 254774 150210
rect 254722 150146 254774 150152
rect 255378 150198 255452 150226
rect 255976 150226 256004 151786
rect 256620 150226 256648 153410
rect 255976 150198 256050 150226
rect 256620 150198 256694 150226
rect 256804 150210 256832 158646
rect 256896 158234 256924 163200
rect 256884 158228 256936 158234
rect 256884 158170 256936 158176
rect 257252 153128 257304 153134
rect 257252 153070 257304 153076
rect 257264 150226 257292 153070
rect 257724 152862 257752 163200
rect 258552 158778 258580 163200
rect 258540 158772 258592 158778
rect 258540 158714 258592 158720
rect 258080 157548 258132 157554
rect 258080 157490 258132 157496
rect 257712 152856 257764 152862
rect 257712 152798 257764 152804
rect 254734 149940 254762 150146
rect 255378 149940 255406 150198
rect 256022 149940 256050 150198
rect 256666 149940 256694 150198
rect 256792 150204 256844 150210
rect 257264 150198 257338 150226
rect 258092 150210 258120 157490
rect 258540 154284 258592 154290
rect 258540 154226 258592 154232
rect 258552 150226 258580 154226
rect 259472 153406 259500 163200
rect 259552 159860 259604 159866
rect 259552 159802 259604 159808
rect 259460 153400 259512 153406
rect 259460 153342 259512 153348
rect 259564 151814 259592 159802
rect 260300 155514 260328 163200
rect 261128 158846 261156 163200
rect 261956 159866 261984 163200
rect 261944 159860 261996 159866
rect 261944 159802 261996 159808
rect 261116 158840 261168 158846
rect 261116 158782 261168 158788
rect 261024 158772 261076 158778
rect 261024 158714 261076 158720
rect 260472 157956 260524 157962
rect 260472 157898 260524 157904
rect 260288 155508 260340 155514
rect 260288 155450 260340 155456
rect 259564 151786 259868 151814
rect 259840 150226 259868 151786
rect 260484 150226 260512 157898
rect 260840 155780 260892 155786
rect 260840 155722 260892 155728
rect 260852 151814 260880 155722
rect 261036 151910 261064 158714
rect 261392 154828 261444 154834
rect 261392 154770 261444 154776
rect 261024 151904 261076 151910
rect 261024 151846 261076 151852
rect 261404 151814 261432 154770
rect 262232 154290 262260 163254
rect 262692 163146 262720 163254
rect 262770 163200 262826 164400
rect 263598 163200 263654 164400
rect 264426 163200 264482 164400
rect 264992 163254 265296 163282
rect 262784 163146 262812 163200
rect 262692 163118 262812 163146
rect 263048 157888 263100 157894
rect 263048 157830 263100 157836
rect 262220 154284 262272 154290
rect 262220 154226 262272 154232
rect 262404 152244 262456 152250
rect 262404 152186 262456 152192
rect 260852 151786 261156 151814
rect 261404 151786 261800 151814
rect 261128 150226 261156 151786
rect 261772 150226 261800 151786
rect 262416 150226 262444 152186
rect 263060 150226 263088 157830
rect 263612 155582 263640 163200
rect 264440 158778 264468 163200
rect 264888 159928 264940 159934
rect 264888 159870 264940 159876
rect 264428 158772 264480 158778
rect 264428 158714 264480 158720
rect 263692 157752 263744 157758
rect 263692 157694 263744 157700
rect 263600 155576 263652 155582
rect 263600 155518 263652 155524
rect 263704 150346 263732 157694
rect 263784 155916 263836 155922
rect 263784 155858 263836 155864
rect 263692 150340 263744 150346
rect 263692 150282 263744 150288
rect 263796 150226 263824 155858
rect 264900 151814 264928 159870
rect 264992 153134 265020 163254
rect 265268 163146 265296 163254
rect 265346 163200 265402 164400
rect 265452 163254 266124 163282
rect 265360 163146 265388 163200
rect 265268 163118 265388 163146
rect 265164 157208 265216 157214
rect 265164 157150 265216 157156
rect 264980 153128 265032 153134
rect 264980 153070 265032 153076
rect 265176 151814 265204 157150
rect 265452 153474 265480 163254
rect 266096 163146 266124 163254
rect 266174 163200 266230 164400
rect 267002 163200 267058 164400
rect 267830 163200 267886 164400
rect 268658 163200 268714 164400
rect 269224 163254 269436 163282
rect 266188 163146 266216 163200
rect 266096 163118 266216 163146
rect 266360 158772 266412 158778
rect 266360 158714 266412 158720
rect 266268 155168 266320 155174
rect 266268 155110 266320 155116
rect 265440 153468 265492 153474
rect 265440 153410 265492 153416
rect 264900 151786 265020 151814
rect 265176 151786 265664 151814
rect 256792 150146 256844 150152
rect 257310 149940 257338 150198
rect 257942 150204 257994 150210
rect 257942 150146 257994 150152
rect 258080 150204 258132 150210
rect 258552 150198 258626 150226
rect 258080 150146 258132 150152
rect 257954 149940 257982 150146
rect 258598 149940 258626 150198
rect 259230 150204 259282 150210
rect 259840 150198 259914 150226
rect 260484 150198 260558 150226
rect 261128 150198 261202 150226
rect 261772 150198 261846 150226
rect 262416 150198 262490 150226
rect 263060 150198 263134 150226
rect 259230 150146 259282 150152
rect 259242 149940 259270 150146
rect 259886 149940 259914 150198
rect 260530 149940 260558 150198
rect 261174 149940 261202 150198
rect 261818 149940 261846 150198
rect 262462 149940 262490 150198
rect 263106 149940 263134 150198
rect 263750 150198 263824 150226
rect 264992 150226 265020 151786
rect 265636 150226 265664 151786
rect 266280 150226 266308 155110
rect 266372 152250 266400 158714
rect 266912 156256 266964 156262
rect 266912 156198 266964 156204
rect 266360 152244 266412 152250
rect 266360 152186 266412 152192
rect 266924 150226 266952 156198
rect 267016 155650 267044 163200
rect 267844 158778 267872 163200
rect 268672 159934 268700 163200
rect 269120 159996 269172 160002
rect 269120 159938 269172 159944
rect 268660 159928 268712 159934
rect 268660 159870 268712 159876
rect 267832 158772 267884 158778
rect 267832 158714 267884 158720
rect 267740 157820 267792 157826
rect 267740 157762 267792 157768
rect 267004 155644 267056 155650
rect 267004 155586 267056 155592
rect 267556 152992 267608 152998
rect 267556 152934 267608 152940
rect 267568 150226 267596 152934
rect 267752 151814 267780 157762
rect 268844 155100 268896 155106
rect 268844 155042 268896 155048
rect 267752 151786 268240 151814
rect 268212 150226 268240 151786
rect 268856 150226 268884 155042
rect 264382 150204 264434 150210
rect 263750 149940 263778 150198
rect 264992 150198 265066 150226
rect 265636 150198 265710 150226
rect 266280 150198 266354 150226
rect 266924 150198 266998 150226
rect 267568 150198 267642 150226
rect 268212 150198 268286 150226
rect 268856 150198 268930 150226
rect 269132 150210 269160 159938
rect 269224 153270 269252 163254
rect 269408 163146 269436 163254
rect 269486 163200 269542 164400
rect 270314 163200 270370 164400
rect 271234 163200 271290 164400
rect 272062 163200 272118 164400
rect 272890 163200 272946 164400
rect 273718 163200 273774 164400
rect 274546 163200 274602 164400
rect 275374 163200 275430 164400
rect 276202 163200 276258 164400
rect 277122 163200 277178 164400
rect 277412 163254 277900 163282
rect 269500 163146 269528 163200
rect 269408 163118 269528 163146
rect 270328 157010 270356 163200
rect 271248 160002 271276 163200
rect 272076 161474 272104 163200
rect 272076 161446 272196 161474
rect 271236 159996 271288 160002
rect 271236 159938 271288 159944
rect 270500 157344 270552 157350
rect 270500 157286 270552 157292
rect 270316 157004 270368 157010
rect 270316 156946 270368 156952
rect 269488 156324 269540 156330
rect 269488 156266 269540 156272
rect 269212 153264 269264 153270
rect 269212 153206 269264 153212
rect 269500 150226 269528 156266
rect 270512 151814 270540 157286
rect 272064 156188 272116 156194
rect 272064 156130 272116 156136
rect 271420 155032 271472 155038
rect 271420 154974 271472 154980
rect 270512 151786 270816 151814
rect 270788 150226 270816 151786
rect 271432 150226 271460 154974
rect 272076 150226 272104 156130
rect 272168 152998 272196 161446
rect 272800 159996 272852 160002
rect 272800 159938 272852 159944
rect 272156 152992 272208 152998
rect 272156 152934 272208 152940
rect 272812 152114 272840 159938
rect 272904 153338 272932 163200
rect 273260 157276 273312 157282
rect 273260 157218 273312 157224
rect 272892 153332 272944 153338
rect 272892 153274 272944 153280
rect 272708 152108 272760 152114
rect 272708 152050 272760 152056
rect 272800 152108 272852 152114
rect 272800 152050 272852 152056
rect 272720 150226 272748 152050
rect 273272 150226 273300 157218
rect 273732 157146 273760 163200
rect 274560 159497 274588 163200
rect 275388 160002 275416 163200
rect 275376 159996 275428 160002
rect 275376 159938 275428 159944
rect 274546 159488 274602 159497
rect 274546 159423 274602 159432
rect 275190 159352 275246 159361
rect 275190 159287 275246 159296
rect 273720 157140 273772 157146
rect 273720 157082 273772 157088
rect 273904 156120 273956 156126
rect 273904 156062 273956 156068
rect 273916 150226 273944 156062
rect 274548 152176 274600 152182
rect 274548 152118 274600 152124
rect 274560 150226 274588 152118
rect 275204 150226 275232 159287
rect 276112 155848 276164 155854
rect 276112 155790 276164 155796
rect 275836 154352 275888 154358
rect 275836 154294 275888 154300
rect 275848 150226 275876 154294
rect 276124 151814 276152 155790
rect 276216 154358 276244 163200
rect 277136 157078 277164 163200
rect 277124 157072 277176 157078
rect 277124 157014 277176 157020
rect 277124 154896 277176 154902
rect 277124 154838 277176 154844
rect 276204 154352 276256 154358
rect 276204 154294 276256 154300
rect 276124 151786 276520 151814
rect 276492 150226 276520 151786
rect 277136 150226 277164 154838
rect 277412 151842 277440 163254
rect 277872 163146 277900 163254
rect 277950 163200 278006 164400
rect 278778 163200 278834 164400
rect 278884 163254 279556 163282
rect 277964 163146 277992 163200
rect 277872 163118 277992 163146
rect 278412 154420 278464 154426
rect 278412 154362 278464 154368
rect 277768 152924 277820 152930
rect 277768 152866 277820 152872
rect 277400 151836 277452 151842
rect 277400 151778 277452 151784
rect 277780 150226 277808 152866
rect 278424 150226 278452 154362
rect 278792 152182 278820 163200
rect 278884 154426 278912 163254
rect 279528 163146 279556 163254
rect 279606 163200 279662 164400
rect 280434 163200 280490 164400
rect 281262 163200 281318 164400
rect 282090 163200 282146 164400
rect 283010 163200 283066 164400
rect 283838 163200 283894 164400
rect 284666 163200 284722 164400
rect 285494 163200 285550 164400
rect 285692 163254 286272 163282
rect 279620 163146 279648 163200
rect 279528 163118 279648 163146
rect 280344 160064 280396 160070
rect 280344 160006 280396 160012
rect 279056 156460 279108 156466
rect 279056 156402 279108 156408
rect 278872 154420 278924 154426
rect 278872 154362 278924 154368
rect 278780 152176 278832 152182
rect 278780 152118 278832 152124
rect 279068 150226 279096 156402
rect 279700 153060 279752 153066
rect 279700 153002 279752 153008
rect 279712 150226 279740 153002
rect 280356 150226 280384 160006
rect 280448 157214 280476 163200
rect 281276 160070 281304 163200
rect 281264 160064 281316 160070
rect 281264 160006 281316 160012
rect 282104 159322 282132 163200
rect 281540 159316 281592 159322
rect 281540 159258 281592 159264
rect 282092 159316 282144 159322
rect 282092 159258 282144 159264
rect 280436 157208 280488 157214
rect 280436 157150 280488 157156
rect 280986 153776 281042 153785
rect 280986 153711 281042 153720
rect 281000 150226 281028 153711
rect 264382 150146 264434 150152
rect 264394 149940 264422 150146
rect 265038 149940 265066 150198
rect 265682 149940 265710 150198
rect 266326 149940 266354 150198
rect 266970 149940 266998 150198
rect 267614 149940 267642 150198
rect 268258 149940 268286 150198
rect 268902 149940 268930 150198
rect 269120 150204 269172 150210
rect 269500 150198 269574 150226
rect 269120 150146 269172 150152
rect 269546 149940 269574 150198
rect 270178 150204 270230 150210
rect 270788 150198 270862 150226
rect 271432 150198 271506 150226
rect 272076 150198 272150 150226
rect 272720 150198 272794 150226
rect 273272 150198 273346 150226
rect 273916 150198 273990 150226
rect 274560 150198 274634 150226
rect 275204 150198 275278 150226
rect 275848 150198 275922 150226
rect 276492 150198 276566 150226
rect 277136 150198 277210 150226
rect 277780 150198 277854 150226
rect 278424 150198 278498 150226
rect 279068 150198 279142 150226
rect 279712 150198 279786 150226
rect 280356 150198 280430 150226
rect 281000 150198 281074 150226
rect 281552 150210 281580 159258
rect 281632 156528 281684 156534
rect 281632 156470 281684 156476
rect 281644 150226 281672 156470
rect 283024 153921 283052 163200
rect 283196 159180 283248 159186
rect 283196 159122 283248 159128
rect 283104 156664 283156 156670
rect 283104 156606 283156 156612
rect 283010 153912 283066 153921
rect 283010 153847 283066 153856
rect 282920 152380 282972 152386
rect 282920 152322 282972 152328
rect 282932 150226 282960 152322
rect 270178 150146 270230 150152
rect 270190 149940 270218 150146
rect 270834 149940 270862 150198
rect 271478 149940 271506 150198
rect 272122 149940 272150 150198
rect 272766 149940 272794 150198
rect 273318 149940 273346 150198
rect 273962 149940 273990 150198
rect 274606 149940 274634 150198
rect 275250 149940 275278 150198
rect 275894 149940 275922 150198
rect 276538 149940 276566 150198
rect 277182 149940 277210 150198
rect 277826 149940 277854 150198
rect 278470 149940 278498 150198
rect 279114 149940 279142 150198
rect 279758 149940 279786 150198
rect 280402 149940 280430 150198
rect 281046 149940 281074 150198
rect 281540 150204 281592 150210
rect 281644 150198 281718 150226
rect 281540 150146 281592 150152
rect 281690 149940 281718 150198
rect 282322 150204 282374 150210
rect 282932 150198 283006 150226
rect 283116 150210 283144 156606
rect 283208 152386 283236 159122
rect 283852 157282 283880 163200
rect 284392 159248 284444 159254
rect 284392 159190 284444 159196
rect 283840 157276 283892 157282
rect 283840 157218 283892 157224
rect 283656 153876 283708 153882
rect 283656 153818 283708 153824
rect 283196 152380 283248 152386
rect 283196 152322 283248 152328
rect 283668 150226 283696 153818
rect 282322 150146 282374 150152
rect 282334 149940 282362 150146
rect 282978 149940 283006 150198
rect 283104 150204 283156 150210
rect 283104 150146 283156 150152
rect 283622 150198 283696 150226
rect 284404 150210 284432 159190
rect 284680 159186 284708 163200
rect 284668 159180 284720 159186
rect 284668 159122 284720 159128
rect 285508 152930 285536 163200
rect 285692 154494 285720 163254
rect 286244 163146 286272 163254
rect 286322 163200 286378 164400
rect 287150 163200 287206 164400
rect 287978 163200 288034 164400
rect 288898 163200 288954 164400
rect 289726 163200 289782 164400
rect 290554 163200 290610 164400
rect 291382 163200 291438 164400
rect 292210 163200 292266 164400
rect 293038 163200 293094 164400
rect 293866 163200 293922 164400
rect 294786 163200 294842 164400
rect 295614 163200 295670 164400
rect 296442 163200 296498 164400
rect 297270 163200 297326 164400
rect 298098 163200 298154 164400
rect 298664 163254 298876 163282
rect 286336 163146 286364 163200
rect 286244 163118 286364 163146
rect 285772 159180 285824 159186
rect 285772 159122 285824 159128
rect 285588 154488 285640 154494
rect 285588 154430 285640 154436
rect 285680 154488 285732 154494
rect 285680 154430 285732 154436
rect 285600 154306 285628 154430
rect 285600 154278 285720 154306
rect 285692 153882 285720 154278
rect 285680 153876 285732 153882
rect 285680 153818 285732 153824
rect 285496 152924 285548 152930
rect 285496 152866 285548 152872
rect 285784 152658 285812 159122
rect 287164 156806 287192 163200
rect 287992 159254 288020 163200
rect 287980 159248 288032 159254
rect 287980 159190 288032 159196
rect 288912 159186 288940 163200
rect 288256 159180 288308 159186
rect 288256 159122 288308 159128
rect 288900 159180 288952 159186
rect 288900 159122 288952 159128
rect 286324 156800 286376 156806
rect 286324 156742 286376 156748
rect 287152 156800 287204 156806
rect 287152 156742 287204 156748
rect 286230 153912 286286 153921
rect 286140 153876 286192 153882
rect 286230 153847 286232 153856
rect 286140 153818 286192 153824
rect 286284 153847 286286 153856
rect 286232 153818 286284 153824
rect 284852 152652 284904 152658
rect 284852 152594 284904 152600
rect 285772 152652 285824 152658
rect 285772 152594 285824 152600
rect 284864 150226 284892 152594
rect 286152 150226 286180 153818
rect 286336 151814 286364 156742
rect 288268 153202 288296 159122
rect 289360 156732 289412 156738
rect 289360 156674 289412 156680
rect 288716 153808 288768 153814
rect 288716 153750 288768 153756
rect 288072 153196 288124 153202
rect 288072 153138 288124 153144
rect 288256 153196 288308 153202
rect 288256 153138 288308 153144
rect 287428 152380 287480 152386
rect 287428 152322 287480 152328
rect 286336 151786 286824 151814
rect 286796 150226 286824 151786
rect 287440 150226 287468 152322
rect 288084 150226 288112 153138
rect 288728 150226 288756 153750
rect 289372 150226 289400 156674
rect 289740 155718 289768 163200
rect 290568 156738 290596 163200
rect 291396 161474 291424 163200
rect 291396 161446 291516 161474
rect 290648 159384 290700 159390
rect 290648 159326 290700 159332
rect 290556 156732 290608 156738
rect 290556 156674 290608 156680
rect 289728 155712 289780 155718
rect 289728 155654 289780 155660
rect 290004 153196 290056 153202
rect 290004 153138 290056 153144
rect 290016 150226 290044 153138
rect 290660 150226 290688 159326
rect 291384 153944 291436 153950
rect 291384 153886 291436 153892
rect 291396 150226 291424 153886
rect 291488 153066 291516 161446
rect 291936 156936 291988 156942
rect 291936 156878 291988 156884
rect 291476 153060 291528 153066
rect 291476 153002 291528 153008
rect 291844 152652 291896 152658
rect 291844 152594 291896 152600
rect 291856 152386 291884 152594
rect 291844 152380 291896 152386
rect 291844 152322 291896 152328
rect 284254 150204 284306 150210
rect 283622 149940 283650 150198
rect 284254 150146 284306 150152
rect 284392 150204 284444 150210
rect 284864 150198 284938 150226
rect 284392 150146 284444 150152
rect 284266 149940 284294 150146
rect 284910 149940 284938 150198
rect 285542 150204 285594 150210
rect 286152 150198 286226 150226
rect 286796 150198 286870 150226
rect 287440 150198 287514 150226
rect 288084 150198 288158 150226
rect 288728 150198 288802 150226
rect 289372 150198 289446 150226
rect 290016 150198 290090 150226
rect 290660 150198 290734 150226
rect 285542 150146 285594 150152
rect 285554 149940 285582 150146
rect 286198 149940 286226 150198
rect 286842 149940 286870 150198
rect 287486 149940 287514 150198
rect 288130 149940 288158 150198
rect 288774 149940 288802 150198
rect 289418 149940 289446 150198
rect 290062 149940 290090 150198
rect 290706 149940 290734 150198
rect 291350 150198 291424 150226
rect 291948 150226 291976 156878
rect 292224 152658 292252 163200
rect 293052 155786 293080 163200
rect 293880 156942 293908 163200
rect 294800 159390 294828 163200
rect 295628 159526 295656 163200
rect 295524 159520 295576 159526
rect 295524 159462 295576 159468
rect 295616 159520 295668 159526
rect 295616 159462 295668 159468
rect 294788 159384 294840 159390
rect 294788 159326 294840 159332
rect 295156 159044 295208 159050
rect 295156 158986 295208 158992
rect 293868 156936 293920 156942
rect 293868 156878 293920 156884
rect 294052 156868 294104 156874
rect 294052 156810 294104 156816
rect 293040 155780 293092 155786
rect 293040 155722 293092 155728
rect 293868 153740 293920 153746
rect 293868 153682 293920 153688
rect 292212 152652 292264 152658
rect 292212 152594 292264 152600
rect 293224 152516 293276 152522
rect 293224 152458 293276 152464
rect 292578 152416 292634 152425
rect 292578 152351 292634 152360
rect 292592 150226 292620 152351
rect 293236 150226 293264 152458
rect 293880 150226 293908 153682
rect 294064 151814 294092 156810
rect 294064 151786 294552 151814
rect 294524 150226 294552 151786
rect 295168 150226 295196 158986
rect 295536 151814 295564 159462
rect 296456 155854 296484 163200
rect 297088 158092 297140 158098
rect 297088 158034 297140 158040
rect 296444 155848 296496 155854
rect 296444 155790 296496 155796
rect 296444 154556 296496 154562
rect 296444 154498 296496 154504
rect 295536 151786 295840 151814
rect 295812 150226 295840 151786
rect 296456 150226 296484 154498
rect 297100 150226 297128 158034
rect 297284 156874 297312 163200
rect 298008 159452 298060 159458
rect 298008 159394 298060 159400
rect 297272 156868 297324 156874
rect 297272 156810 297324 156816
rect 297732 152584 297784 152590
rect 297732 152526 297784 152532
rect 297744 150226 297772 152526
rect 298020 151814 298048 159394
rect 298112 159050 298140 163200
rect 298100 159044 298152 159050
rect 298100 158986 298152 158992
rect 298664 152522 298692 163254
rect 298848 163146 298876 163254
rect 298926 163200 298982 164400
rect 299754 163200 299810 164400
rect 300674 163200 300730 164400
rect 301502 163200 301558 164400
rect 302330 163200 302386 164400
rect 303158 163200 303214 164400
rect 303724 163254 303936 163282
rect 298940 163146 298968 163200
rect 298848 163118 298968 163146
rect 299480 158976 299532 158982
rect 299480 158918 299532 158924
rect 299020 154012 299072 154018
rect 299020 153954 299072 153960
rect 298652 152516 298704 152522
rect 298652 152458 298704 152464
rect 298020 151786 298416 151814
rect 298388 150226 298416 151786
rect 299032 150226 299060 153954
rect 291948 150198 292022 150226
rect 292592 150198 292666 150226
rect 293236 150198 293310 150226
rect 293880 150198 293954 150226
rect 294524 150198 294598 150226
rect 295168 150198 295242 150226
rect 295812 150198 295886 150226
rect 296456 150198 296530 150226
rect 297100 150198 297174 150226
rect 297744 150198 297818 150226
rect 298388 150198 298462 150226
rect 299032 150198 299106 150226
rect 299492 150210 299520 158918
rect 299768 155922 299796 163200
rect 300688 158098 300716 163200
rect 301412 159724 301464 159730
rect 301412 159666 301464 159672
rect 300768 159044 300820 159050
rect 300768 158986 300820 158992
rect 300676 158092 300728 158098
rect 300676 158034 300728 158040
rect 299756 155916 299808 155922
rect 299756 155858 299808 155864
rect 299664 155236 299716 155242
rect 299664 155178 299716 155184
rect 299676 150226 299704 155178
rect 300780 152130 300808 158986
rect 301424 158982 301452 159666
rect 301516 159458 301544 163200
rect 302344 159662 302372 163200
rect 302332 159656 302384 159662
rect 302332 159598 302384 159604
rect 301504 159452 301556 159458
rect 301504 159394 301556 159400
rect 301412 158976 301464 158982
rect 301412 158918 301464 158924
rect 302240 158024 302292 158030
rect 302240 157966 302292 157972
rect 301596 153672 301648 153678
rect 301596 153614 301648 153620
rect 300780 152102 301084 152130
rect 301056 152046 301084 152102
rect 300952 152040 301004 152046
rect 300952 151982 301004 151988
rect 301044 152040 301096 152046
rect 301044 151982 301096 151988
rect 300964 150226 300992 151982
rect 301608 150226 301636 153614
rect 302252 150226 302280 157966
rect 303172 155242 303200 163200
rect 303528 159724 303580 159730
rect 303528 159666 303580 159672
rect 303160 155236 303212 155242
rect 303160 155178 303212 155184
rect 302884 151972 302936 151978
rect 302884 151914 302936 151920
rect 302896 150226 302924 151914
rect 303540 150226 303568 159666
rect 303724 153202 303752 163254
rect 303908 163146 303936 163254
rect 303986 163200 304042 164400
rect 304814 163200 304870 164400
rect 305642 163200 305698 164400
rect 306562 163200 306618 164400
rect 307390 163200 307446 164400
rect 308218 163200 308274 164400
rect 309046 163200 309102 164400
rect 309874 163200 309930 164400
rect 310702 163200 310758 164400
rect 311530 163200 311586 164400
rect 312450 163200 312506 164400
rect 313278 163200 313334 164400
rect 314106 163200 314162 164400
rect 314934 163200 314990 164400
rect 315762 163200 315818 164400
rect 316590 163200 316646 164400
rect 317418 163200 317474 164400
rect 318338 163200 318394 164400
rect 319166 163200 319222 164400
rect 319272 163254 319944 163282
rect 304000 163146 304028 163200
rect 303908 163118 304028 163146
rect 304724 155304 304776 155310
rect 304724 155246 304776 155252
rect 304080 154080 304132 154086
rect 304080 154022 304132 154028
rect 303712 153196 303764 153202
rect 303712 153138 303764 153144
rect 304092 150226 304120 154022
rect 304736 150226 304764 155246
rect 304828 152590 304856 163200
rect 305656 158914 305684 163200
rect 305368 158908 305420 158914
rect 305368 158850 305420 158856
rect 305644 158908 305696 158914
rect 305644 158850 305696 158856
rect 304816 152584 304868 152590
rect 304816 152526 304868 152532
rect 305380 150226 305408 158850
rect 306576 155310 306604 163200
rect 307404 159118 307432 163200
rect 307392 159112 307444 159118
rect 307392 159054 307444 159060
rect 308232 159050 308260 163200
rect 309060 159730 309088 163200
rect 309888 161474 309916 163200
rect 309888 161446 310008 161474
rect 309048 159724 309100 159730
rect 309048 159666 309100 159672
rect 308220 159044 308272 159050
rect 308220 158986 308272 158992
rect 308588 158976 308640 158982
rect 308588 158918 308640 158924
rect 307668 158908 307720 158914
rect 307668 158850 307720 158856
rect 306932 158160 306984 158166
rect 306932 158102 306984 158108
rect 306564 155304 306616 155310
rect 306564 155246 306616 155252
rect 306656 153604 306708 153610
rect 306656 153546 306708 153552
rect 306012 152788 306064 152794
rect 306012 152730 306064 152736
rect 306024 150226 306052 152730
rect 306668 150226 306696 153546
rect 306944 151814 306972 158102
rect 307680 152794 307708 158850
rect 307668 152788 307720 152794
rect 307668 152730 307720 152736
rect 307944 152720 307996 152726
rect 307944 152662 307996 152668
rect 306944 151786 307340 151814
rect 307312 150226 307340 151786
rect 307956 150226 307984 152662
rect 308600 150226 308628 158918
rect 309876 155372 309928 155378
rect 309876 155314 309928 155320
rect 309232 154148 309284 154154
rect 309232 154090 309284 154096
rect 309244 150226 309272 154090
rect 309888 150226 309916 155314
rect 309980 155174 310008 161446
rect 310612 159588 310664 159594
rect 310612 159530 310664 159536
rect 309968 155168 310020 155174
rect 309968 155110 310020 155116
rect 310624 150226 310652 159530
rect 310716 158914 310744 163200
rect 310704 158908 310756 158914
rect 310704 158850 310756 158856
rect 311544 152726 311572 163200
rect 312464 158914 312492 163200
rect 311992 158908 312044 158914
rect 311992 158850 312044 158856
rect 312452 158908 312504 158914
rect 312452 158850 312504 158856
rect 311808 153536 311860 153542
rect 311808 153478 311860 153484
rect 311532 152720 311584 152726
rect 311532 152662 311584 152668
rect 311164 152448 311216 152454
rect 311164 152390 311216 152396
rect 291350 149940 291378 150198
rect 291994 149940 292022 150198
rect 292638 149940 292666 150198
rect 293282 149940 293310 150198
rect 293926 149940 293954 150198
rect 294570 149940 294598 150198
rect 295214 149940 295242 150198
rect 295858 149940 295886 150198
rect 296502 149940 296530 150198
rect 297146 149940 297174 150198
rect 297790 149940 297818 150198
rect 298434 149940 298462 150198
rect 299078 149940 299106 150198
rect 299480 150204 299532 150210
rect 299676 150198 299750 150226
rect 299480 150146 299532 150152
rect 299722 149940 299750 150198
rect 300354 150204 300406 150210
rect 300964 150198 301038 150226
rect 301608 150198 301682 150226
rect 302252 150198 302326 150226
rect 302896 150198 302970 150226
rect 303540 150198 303614 150226
rect 304092 150198 304166 150226
rect 304736 150198 304810 150226
rect 305380 150198 305454 150226
rect 306024 150198 306098 150226
rect 306668 150198 306742 150226
rect 307312 150198 307386 150226
rect 307956 150198 308030 150226
rect 308600 150198 308674 150226
rect 309244 150198 309318 150226
rect 309888 150198 309962 150226
rect 300354 150146 300406 150152
rect 300366 149940 300394 150146
rect 301010 149940 301038 150198
rect 301654 149940 301682 150198
rect 302298 149940 302326 150198
rect 302942 149940 302970 150198
rect 303586 149940 303614 150198
rect 304138 149940 304166 150198
rect 304782 149940 304810 150198
rect 305426 149940 305454 150198
rect 306070 149940 306098 150198
rect 306714 149940 306742 150198
rect 307358 149940 307386 150198
rect 308002 149940 308030 150198
rect 308646 149940 308674 150198
rect 309290 149940 309318 150198
rect 309934 149940 309962 150198
rect 310578 150198 310652 150226
rect 311176 150226 311204 152390
rect 311820 150226 311848 153478
rect 312004 152454 312032 158850
rect 312452 155440 312504 155446
rect 312452 155382 312504 155388
rect 311992 152448 312044 152454
rect 311992 152390 312044 152396
rect 312464 150226 312492 155382
rect 313292 153950 313320 163200
rect 314120 159798 314148 163200
rect 313372 159792 313424 159798
rect 313372 159734 313424 159740
rect 314108 159792 314160 159798
rect 314108 159734 314160 159740
rect 313280 153944 313332 153950
rect 313280 153886 313332 153892
rect 313096 152312 313148 152318
rect 313096 152254 313148 152260
rect 313108 150226 313136 152254
rect 313384 151814 313412 159734
rect 314948 158982 314976 163200
rect 315776 159594 315804 163200
rect 315764 159588 315816 159594
rect 315764 159530 315816 159536
rect 314936 158976 314988 158982
rect 314936 158918 314988 158924
rect 313464 158908 313516 158914
rect 313464 158850 313516 158856
rect 313476 152425 313504 158850
rect 315028 158228 315080 158234
rect 315028 158170 315080 158176
rect 314384 154216 314436 154222
rect 314384 154158 314436 154164
rect 313462 152416 313518 152425
rect 313462 152351 313518 152360
rect 313384 151786 313780 151814
rect 313752 150226 313780 151786
rect 314396 150226 314424 154158
rect 315040 150226 315068 158170
rect 316604 155378 316632 163200
rect 317052 158840 317104 158846
rect 317052 158782 317104 158788
rect 316592 155372 316644 155378
rect 316592 155314 316644 155320
rect 316960 153400 317012 153406
rect 316960 153342 317012 153348
rect 315672 152856 315724 152862
rect 315672 152798 315724 152804
rect 315684 150226 315712 152798
rect 316316 151904 316368 151910
rect 316316 151846 316368 151852
rect 316328 150226 316356 151846
rect 316972 150226 317000 153342
rect 317064 152862 317092 158782
rect 317052 152856 317104 152862
rect 317052 152798 317104 152804
rect 317432 151978 317460 163200
rect 317604 155508 317656 155514
rect 317604 155450 317656 155456
rect 317420 151972 317472 151978
rect 317420 151914 317472 151920
rect 317616 150226 317644 155450
rect 318352 152862 318380 163200
rect 318800 159860 318852 159866
rect 318800 159802 318852 159808
rect 318248 152856 318300 152862
rect 318248 152798 318300 152804
rect 318340 152856 318392 152862
rect 318340 152798 318392 152804
rect 318260 150226 318288 152798
rect 318812 151814 318840 159802
rect 319180 158778 319208 163200
rect 319168 158772 319220 158778
rect 319168 158714 319220 158720
rect 319272 154018 319300 163254
rect 319916 163146 319944 163254
rect 319994 163200 320050 164400
rect 320822 163200 320878 164400
rect 321650 163200 321706 164400
rect 322478 163200 322534 164400
rect 323306 163200 323362 164400
rect 324226 163200 324282 164400
rect 324332 163254 325004 163282
rect 320008 163146 320036 163200
rect 319916 163118 320036 163146
rect 320836 159866 320864 163200
rect 320824 159860 320876 159866
rect 320824 159802 320876 159808
rect 320272 158840 320324 158846
rect 320272 158782 320324 158788
rect 320180 155576 320232 155582
rect 320180 155518 320232 155524
rect 319536 154284 319588 154290
rect 319536 154226 319588 154232
rect 319260 154012 319312 154018
rect 319260 153954 319312 153960
rect 318812 151786 318932 151814
rect 318904 150226 318932 151786
rect 319548 150226 319576 154226
rect 320192 150226 320220 155518
rect 320284 152318 320312 158782
rect 321664 158778 321692 163200
rect 322492 158914 322520 163200
rect 322480 158908 322532 158914
rect 322480 158850 322532 158856
rect 321560 158772 321612 158778
rect 321560 158714 321612 158720
rect 321652 158772 321704 158778
rect 321652 158714 321704 158720
rect 321468 153128 321520 153134
rect 321468 153070 321520 153076
rect 320732 152992 320784 152998
rect 320732 152934 320784 152940
rect 320272 152312 320324 152318
rect 320272 152254 320324 152260
rect 320744 151910 320772 152934
rect 320824 152244 320876 152250
rect 320824 152186 320876 152192
rect 320916 152244 320968 152250
rect 320916 152186 320968 152192
rect 320732 151904 320784 151910
rect 320732 151846 320784 151852
rect 320836 150226 320864 152186
rect 320928 151978 320956 152186
rect 320916 151972 320968 151978
rect 320916 151914 320968 151920
rect 321480 150226 321508 153070
rect 321572 151978 321600 158714
rect 321744 155644 321796 155650
rect 321744 155586 321796 155592
rect 321560 151972 321612 151978
rect 321560 151914 321612 151920
rect 311176 150198 311250 150226
rect 311820 150198 311894 150226
rect 312464 150198 312538 150226
rect 313108 150198 313182 150226
rect 313752 150198 313826 150226
rect 314396 150198 314470 150226
rect 315040 150198 315114 150226
rect 315684 150198 315758 150226
rect 316328 150198 316402 150226
rect 316972 150198 317046 150226
rect 317616 150198 317690 150226
rect 318260 150198 318334 150226
rect 318904 150198 318978 150226
rect 319548 150198 319622 150226
rect 320192 150198 320266 150226
rect 320836 150198 320910 150226
rect 321480 150198 321554 150226
rect 321756 150210 321784 155586
rect 323320 154086 323348 163200
rect 324044 159928 324096 159934
rect 324044 159870 324096 159876
rect 323308 154080 323360 154086
rect 323308 154022 323360 154028
rect 322204 153468 322256 153474
rect 322204 153410 322256 153416
rect 322216 150226 322244 153410
rect 323124 152312 323176 152318
rect 323124 152254 323176 152260
rect 323136 151814 323164 152254
rect 323136 151786 323440 151814
rect 310578 149940 310606 150198
rect 311222 149940 311250 150198
rect 311866 149940 311894 150198
rect 312510 149940 312538 150198
rect 313154 149940 313182 150198
rect 313798 149940 313826 150198
rect 314442 149940 314470 150198
rect 315086 149940 315114 150198
rect 315730 149940 315758 150198
rect 316374 149940 316402 150198
rect 317018 149940 317046 150198
rect 317662 149940 317690 150198
rect 318306 149940 318334 150198
rect 318950 149940 318978 150198
rect 319594 149940 319622 150198
rect 320238 149940 320266 150198
rect 320882 149940 320910 150198
rect 321526 149940 321554 150198
rect 321744 150204 321796 150210
rect 321744 150146 321796 150152
rect 322170 150198 322244 150226
rect 323412 150226 323440 151786
rect 324056 150226 324084 159870
rect 324240 153134 324268 163200
rect 324228 153128 324280 153134
rect 324228 153070 324280 153076
rect 324332 152250 324360 163254
rect 324976 163146 325004 163254
rect 325054 163200 325110 164400
rect 325882 163200 325938 164400
rect 326710 163200 326766 164400
rect 327538 163200 327594 164400
rect 328366 163200 328422 164400
rect 329194 163200 329250 164400
rect 330114 163200 330170 164400
rect 330942 163200 330998 164400
rect 331232 163254 331720 163282
rect 325068 163146 325096 163200
rect 324976 163118 325096 163146
rect 325332 157004 325384 157010
rect 325332 156946 325384 156952
rect 324688 153264 324740 153270
rect 324688 153206 324740 153212
rect 324320 152244 324372 152250
rect 324320 152186 324372 152192
rect 324700 150226 324728 153206
rect 325344 150226 325372 156946
rect 325896 151978 325924 163200
rect 326724 154154 326752 163200
rect 327552 158846 327580 163200
rect 328380 159934 328408 163200
rect 329208 160002 329236 163200
rect 329104 159996 329156 160002
rect 329104 159938 329156 159944
rect 329196 159996 329248 160002
rect 329196 159938 329248 159944
rect 328368 159928 328420 159934
rect 328368 159870 328420 159876
rect 328550 159488 328606 159497
rect 328550 159423 328606 159432
rect 327540 158840 327592 158846
rect 327540 158782 327592 158788
rect 327908 157140 327960 157146
rect 327908 157082 327960 157088
rect 326712 154148 326764 154154
rect 326712 154090 326764 154096
rect 327264 153332 327316 153338
rect 327264 153274 327316 153280
rect 325976 152108 326028 152114
rect 325976 152050 326028 152056
rect 325608 151972 325660 151978
rect 325608 151914 325660 151920
rect 325884 151972 325936 151978
rect 325884 151914 325936 151920
rect 325620 151774 325648 151914
rect 325608 151768 325660 151774
rect 325608 151710 325660 151716
rect 325988 150226 326016 152050
rect 326620 151904 326672 151910
rect 326620 151846 326672 151852
rect 326632 150226 326660 151846
rect 327276 150226 327304 153274
rect 327920 150226 327948 157082
rect 328564 150226 328592 159423
rect 329116 151814 329144 159938
rect 330128 155446 330156 163200
rect 330484 158840 330536 158846
rect 330536 158788 330708 158794
rect 330484 158782 330708 158788
rect 330496 158778 330708 158782
rect 330496 158772 330720 158778
rect 330496 158766 330668 158772
rect 330668 158714 330720 158720
rect 330484 157072 330536 157078
rect 330484 157014 330536 157020
rect 330116 155440 330168 155446
rect 330116 155382 330168 155388
rect 329932 154352 329984 154358
rect 329932 154294 329984 154300
rect 329116 151786 329236 151814
rect 329208 150226 329236 151786
rect 329944 150226 329972 154294
rect 322802 150204 322854 150210
rect 322170 149940 322198 150198
rect 323412 150198 323486 150226
rect 324056 150198 324130 150226
rect 324700 150198 324774 150226
rect 325344 150198 325418 150226
rect 325988 150198 326062 150226
rect 326632 150198 326706 150226
rect 327276 150198 327350 150226
rect 327920 150198 327994 150226
rect 328564 150198 328638 150226
rect 329208 150198 329282 150226
rect 322802 150146 322854 150152
rect 322814 149940 322842 150146
rect 323458 149940 323486 150198
rect 324102 149940 324130 150198
rect 324746 149940 324774 150198
rect 325390 149940 325418 150198
rect 326034 149940 326062 150198
rect 326678 149940 326706 150198
rect 327322 149940 327350 150198
rect 327966 149940 327994 150198
rect 328610 149940 328638 150198
rect 329254 149940 329282 150198
rect 329898 150198 329972 150226
rect 330496 150226 330524 157014
rect 330956 152998 330984 163200
rect 331232 153542 331260 163254
rect 331692 163146 331720 163254
rect 331770 163200 331826 164400
rect 332598 163200 332654 164400
rect 333426 163200 333482 164400
rect 334254 163200 334310 164400
rect 335082 163200 335138 164400
rect 335372 163254 335952 163282
rect 331784 163146 331812 163200
rect 331692 163118 331812 163146
rect 332416 154420 332468 154426
rect 332416 154362 332468 154368
rect 331220 153536 331272 153542
rect 331220 153478 331272 153484
rect 330944 152992 330996 152998
rect 330944 152934 330996 152940
rect 331772 152176 331824 152182
rect 331772 152118 331824 152124
rect 331128 151904 331180 151910
rect 331128 151846 331180 151852
rect 331140 150226 331168 151846
rect 330496 150198 330570 150226
rect 331140 150198 331214 150226
rect 329898 149940 329926 150198
rect 330542 149940 330570 150198
rect 331186 149940 331214 150198
rect 331784 150090 331812 152118
rect 332428 150090 332456 154362
rect 332612 151910 332640 163200
rect 332692 160064 332744 160070
rect 332692 160006 332744 160012
rect 332704 157334 332732 160006
rect 332704 157306 333376 157334
rect 333060 157208 333112 157214
rect 333060 157150 333112 157156
rect 332600 151904 332652 151910
rect 332600 151846 332652 151852
rect 333072 150090 333100 157150
rect 333348 150226 333376 157306
rect 333440 155514 333468 163200
rect 334268 159322 334296 163200
rect 335096 160070 335124 163200
rect 335084 160064 335136 160070
rect 335084 160006 335136 160012
rect 334164 159316 334216 159322
rect 334164 159258 334216 159264
rect 334256 159316 334308 159322
rect 334256 159258 334308 159264
rect 334176 157334 334204 159258
rect 334176 157306 334388 157334
rect 333428 155508 333480 155514
rect 333428 155450 333480 155456
rect 334360 150226 334388 157306
rect 334900 153876 334952 153882
rect 334900 153818 334952 153824
rect 333348 150198 333790 150226
rect 334360 150198 334434 150226
rect 331784 150062 331858 150090
rect 332428 150062 332502 150090
rect 333072 150062 333146 150090
rect 331830 149940 331858 150062
rect 332474 149940 332502 150062
rect 333118 149940 333146 150062
rect 333762 149940 333790 150198
rect 334406 149940 334434 150198
rect 334912 150090 334940 153818
rect 335372 152114 335400 163254
rect 335924 163146 335952 163254
rect 336002 163200 336058 164400
rect 336830 163200 336886 164400
rect 337658 163200 337714 164400
rect 338486 163200 338542 164400
rect 339314 163200 339370 164400
rect 339512 163254 340092 163282
rect 336016 163146 336044 163200
rect 335924 163118 336044 163146
rect 335544 157276 335596 157282
rect 335544 157218 335596 157224
rect 335360 152108 335412 152114
rect 335360 152050 335412 152056
rect 335556 150090 335584 157218
rect 336844 154290 336872 163200
rect 337672 156670 337700 163200
rect 338500 159186 338528 163200
rect 339328 159254 339356 163200
rect 338764 159248 338816 159254
rect 338764 159190 338816 159196
rect 339316 159248 339368 159254
rect 339316 159190 339368 159196
rect 338396 159180 338448 159186
rect 338396 159122 338448 159128
rect 338488 159180 338540 159186
rect 338488 159122 338540 159128
rect 338120 156800 338172 156806
rect 338120 156742 338172 156748
rect 337660 156664 337712 156670
rect 337660 156606 337712 156612
rect 337476 154488 337528 154494
rect 337476 154430 337528 154436
rect 336832 154284 336884 154290
rect 336832 154226 336884 154232
rect 337016 153536 337068 153542
rect 337016 153478 337068 153484
rect 335740 153066 335952 153082
rect 335728 153060 335952 153066
rect 335780 153054 335952 153060
rect 335728 153002 335780 153008
rect 335924 152930 335952 153054
rect 336096 153060 336148 153066
rect 336096 153002 336148 153008
rect 335820 152924 335872 152930
rect 335820 152866 335872 152872
rect 335912 152924 335964 152930
rect 335912 152866 335964 152872
rect 335832 152182 335860 152866
rect 336108 152674 336136 153002
rect 335924 152646 336136 152674
rect 335924 152522 335952 152646
rect 335912 152516 335964 152522
rect 335912 152458 335964 152464
rect 336004 152516 336056 152522
rect 336004 152458 336056 152464
rect 335820 152176 335872 152182
rect 335820 152118 335872 152124
rect 336016 152046 336044 152458
rect 336188 152380 336240 152386
rect 336188 152322 336240 152328
rect 336004 152040 336056 152046
rect 336004 151982 336056 151988
rect 336200 150090 336228 152322
rect 336832 152176 336884 152182
rect 336832 152118 336884 152124
rect 336924 152176 336976 152182
rect 336924 152118 336976 152124
rect 336844 150090 336872 152118
rect 336936 151910 336964 152118
rect 337028 151910 337056 153478
rect 336924 151904 336976 151910
rect 336924 151846 336976 151852
rect 337016 151904 337068 151910
rect 337016 151846 337068 151852
rect 337488 150090 337516 154430
rect 338132 150090 338160 156742
rect 338408 150210 338436 159122
rect 338776 150226 338804 159190
rect 339512 153882 339540 163254
rect 340064 163146 340092 163254
rect 340142 163200 340198 164400
rect 340970 163200 341026 164400
rect 341890 163200 341946 164400
rect 342718 163200 342774 164400
rect 342824 163254 343496 163282
rect 340156 163146 340184 163200
rect 340064 163118 340184 163146
rect 340788 159180 340840 159186
rect 340788 159122 340840 159128
rect 340696 156732 340748 156738
rect 340696 156674 340748 156680
rect 340052 155712 340104 155718
rect 340052 155654 340104 155660
rect 339500 153876 339552 153882
rect 339500 153818 339552 153824
rect 338396 150204 338448 150210
rect 338776 150198 338850 150226
rect 338396 150146 338448 150152
rect 334912 150062 334986 150090
rect 335556 150062 335630 150090
rect 336200 150062 336274 150090
rect 336844 150062 336918 150090
rect 337488 150062 337562 150090
rect 338132 150062 338206 150090
rect 334958 149940 334986 150062
rect 335602 149940 335630 150062
rect 336246 149940 336274 150062
rect 336890 149940 336918 150062
rect 337534 149940 337562 150062
rect 338178 149940 338206 150062
rect 338822 149940 338850 150198
rect 339454 150204 339506 150210
rect 339454 150146 339506 150152
rect 339466 149940 339494 150146
rect 340064 150090 340092 155654
rect 340708 150090 340736 156674
rect 340800 153082 340828 159122
rect 340984 155582 341012 163200
rect 341904 159186 341932 163200
rect 342444 159520 342496 159526
rect 342444 159462 342496 159468
rect 342260 159384 342312 159390
rect 342260 159326 342312 159332
rect 341892 159180 341944 159186
rect 341892 159122 341944 159128
rect 340972 155576 341024 155582
rect 340972 155518 341024 155524
rect 340800 153054 341472 153082
rect 341444 152930 341472 153054
rect 341340 152924 341392 152930
rect 341340 152866 341392 152872
rect 341432 152924 341484 152930
rect 341432 152866 341484 152872
rect 341352 150226 341380 152866
rect 342272 152658 342300 159326
rect 342352 155780 342404 155786
rect 342352 155722 342404 155728
rect 341984 152652 342036 152658
rect 341984 152594 342036 152600
rect 342260 152652 342312 152658
rect 342260 152594 342312 152600
rect 341996 150226 342024 152594
rect 342364 151814 342392 155722
rect 342456 152046 342484 159462
rect 342732 159390 342760 163200
rect 342720 159384 342772 159390
rect 342720 159326 342772 159332
rect 342720 156936 342772 156942
rect 342720 156878 342772 156884
rect 342444 152040 342496 152046
rect 342444 151982 342496 151988
rect 342732 151814 342760 156878
rect 342824 154222 342852 163254
rect 343468 163146 343496 163254
rect 343546 163200 343602 164400
rect 344374 163200 344430 164400
rect 345202 163200 345258 164400
rect 346030 163200 346086 164400
rect 346412 163254 346808 163282
rect 343560 163146 343588 163200
rect 343468 163118 343588 163146
rect 343640 159384 343692 159390
rect 343640 159326 343692 159332
rect 342812 154216 342864 154222
rect 342812 154158 342864 154164
rect 343652 152386 343680 159326
rect 344388 156738 344416 163200
rect 345216 161474 345244 163200
rect 345216 161446 345336 161474
rect 345112 156868 345164 156874
rect 345112 156810 345164 156816
rect 344376 156732 344428 156738
rect 344376 156674 344428 156680
rect 343916 152652 343968 152658
rect 343916 152594 343968 152600
rect 343640 152380 343692 152386
rect 343640 152322 343692 152328
rect 342364 151786 342668 151814
rect 342732 151786 343312 151814
rect 342640 150226 342668 151786
rect 343284 150226 343312 151786
rect 343928 150226 343956 152594
rect 344560 152040 344612 152046
rect 344560 151982 344612 151988
rect 344572 150226 344600 151982
rect 341352 150198 341426 150226
rect 341996 150198 342070 150226
rect 342640 150198 342714 150226
rect 343284 150198 343358 150226
rect 343928 150198 344002 150226
rect 344572 150198 344646 150226
rect 345124 150210 345152 156810
rect 345204 155848 345256 155854
rect 345204 155790 345256 155796
rect 345216 150226 345244 155790
rect 345308 152658 345336 161446
rect 346044 159390 346072 163200
rect 346032 159384 346084 159390
rect 346032 159326 346084 159332
rect 346412 154358 346440 163254
rect 346780 163146 346808 163254
rect 346858 163200 346914 164400
rect 347778 163200 347834 164400
rect 347976 163254 348556 163282
rect 346872 163146 346900 163200
rect 346780 163118 346900 163146
rect 347688 159520 347740 159526
rect 347688 159462 347740 159468
rect 347700 159050 347728 159462
rect 347792 159050 347820 163200
rect 347688 159044 347740 159050
rect 347688 158986 347740 158992
rect 347780 159044 347832 159050
rect 347780 158986 347832 158992
rect 347872 155916 347924 155922
rect 347872 155858 347924 155864
rect 346400 154352 346452 154358
rect 346400 154294 346452 154300
rect 347136 153060 347188 153066
rect 347136 153002 347188 153008
rect 345296 152652 345348 152658
rect 345296 152594 345348 152600
rect 346492 152516 346544 152522
rect 346492 152458 346544 152464
rect 346504 150226 346532 152458
rect 347148 150226 347176 153002
rect 347884 150226 347912 155858
rect 347976 152522 348004 163254
rect 348528 163146 348556 163254
rect 348606 163200 348662 164400
rect 349172 163254 349384 163282
rect 348620 163146 348648 163200
rect 348528 163118 348648 163146
rect 349068 159452 349120 159458
rect 349068 159394 349120 159400
rect 348056 158092 348108 158098
rect 348056 158034 348108 158040
rect 347964 152516 348016 152522
rect 347964 152458 348016 152464
rect 348068 151814 348096 158034
rect 348068 151786 348464 151814
rect 340064 150062 340138 150090
rect 340708 150062 340782 150090
rect 340110 149940 340138 150062
rect 340754 149940 340782 150062
rect 341398 149940 341426 150198
rect 342042 149940 342070 150198
rect 342686 149940 342714 150198
rect 343330 149940 343358 150198
rect 343974 149940 344002 150198
rect 344618 149940 344646 150198
rect 345112 150204 345164 150210
rect 345216 150198 345290 150226
rect 345112 150146 345164 150152
rect 345262 149940 345290 150198
rect 345894 150204 345946 150210
rect 346504 150198 346578 150226
rect 347148 150198 347222 150226
rect 345894 150146 345946 150152
rect 345906 149940 345934 150146
rect 346550 149940 346578 150198
rect 347194 149940 347222 150198
rect 347838 150198 347912 150226
rect 348436 150226 348464 151786
rect 349080 150226 349108 159394
rect 349172 153066 349200 163254
rect 349356 163146 349384 163254
rect 349434 163200 349490 164400
rect 349540 163254 350212 163282
rect 349448 163146 349476 163200
rect 349356 163118 349476 163146
rect 349252 159656 349304 159662
rect 349252 159598 349304 159604
rect 349160 153060 349212 153066
rect 349160 153002 349212 153008
rect 349264 151814 349292 159598
rect 349344 159452 349396 159458
rect 349344 159394 349396 159400
rect 349356 159118 349384 159394
rect 349344 159112 349396 159118
rect 349344 159054 349396 159060
rect 349540 154426 349568 163254
rect 350184 163146 350212 163254
rect 350262 163200 350318 164400
rect 351090 163200 351146 164400
rect 351918 163200 351974 164400
rect 352024 163254 352696 163282
rect 350276 163146 350304 163200
rect 350184 163118 350304 163146
rect 351104 159118 351132 163200
rect 351932 159662 351960 163200
rect 351920 159656 351972 159662
rect 351920 159598 351972 159604
rect 351092 159112 351144 159118
rect 351092 159054 351144 159060
rect 350356 155236 350408 155242
rect 350356 155178 350408 155184
rect 349528 154420 349580 154426
rect 349528 154362 349580 154368
rect 349264 151786 349752 151814
rect 349724 150226 349752 151786
rect 350368 150226 350396 155178
rect 352024 153202 352052 163254
rect 352668 163146 352696 163254
rect 352746 163200 352802 164400
rect 353666 163200 353722 164400
rect 354494 163200 354550 164400
rect 354692 163254 355272 163282
rect 352760 163146 352788 163200
rect 352668 163118 352788 163146
rect 353208 159452 353260 159458
rect 353208 159394 353260 159400
rect 352472 155304 352524 155310
rect 352472 155246 352524 155252
rect 351000 153196 351052 153202
rect 351000 153138 351052 153144
rect 352012 153196 352064 153202
rect 352012 153138 352064 153144
rect 351012 150226 351040 153138
rect 352288 152788 352340 152794
rect 352288 152730 352340 152736
rect 351644 152584 351696 152590
rect 351644 152526 351696 152532
rect 351656 150226 351684 152526
rect 352300 150226 352328 152730
rect 352484 151814 352512 155246
rect 353220 151814 353248 159394
rect 353680 154562 353708 163200
rect 354220 159520 354272 159526
rect 354220 159462 354272 159468
rect 353668 154556 353720 154562
rect 353668 154498 353720 154504
rect 352484 151786 352972 151814
rect 353220 151786 353616 151814
rect 352944 150226 352972 151786
rect 353588 150226 353616 151786
rect 354232 150226 354260 159462
rect 354508 152590 354536 163200
rect 354496 152584 354548 152590
rect 354496 152526 354548 152532
rect 354692 152046 354720 163254
rect 355244 163146 355272 163254
rect 355322 163200 355378 164400
rect 356150 163200 356206 164400
rect 356256 163254 356928 163282
rect 355336 163146 355364 163200
rect 355244 163118 355364 163146
rect 354864 159724 354916 159730
rect 354864 159666 354916 159672
rect 354680 152040 354732 152046
rect 354680 151982 354732 151988
rect 354876 150226 354904 159666
rect 356164 159526 356192 163200
rect 356152 159520 356204 159526
rect 356152 159462 356204 159468
rect 355508 155168 355560 155174
rect 355508 155110 355560 155116
rect 355520 150226 355548 155110
rect 356256 154494 356284 163254
rect 356900 163146 356928 163254
rect 356978 163200 357034 164400
rect 357806 163200 357862 164400
rect 358634 163200 358690 164400
rect 358832 163254 359504 163282
rect 356992 163146 357020 163200
rect 356900 163118 357020 163146
rect 357820 159730 357848 163200
rect 357992 159792 358044 159798
rect 357992 159734 358044 159740
rect 357808 159724 357860 159730
rect 357808 159666 357860 159672
rect 357440 158976 357492 158982
rect 357440 158918 357492 158924
rect 356244 154488 356296 154494
rect 356244 154430 356296 154436
rect 357452 152794 357480 158918
rect 357808 153944 357860 153950
rect 357808 153886 357860 153892
rect 357440 152788 357492 152794
rect 357440 152730 357492 152736
rect 356796 152720 356848 152726
rect 356796 152662 356848 152668
rect 356152 152448 356204 152454
rect 356152 152390 356204 152396
rect 356164 150226 356192 152390
rect 356808 150226 356836 152662
rect 357438 152416 357494 152425
rect 357438 152351 357494 152360
rect 357452 150226 357480 152351
rect 357820 151814 357848 153886
rect 358004 151814 358032 159734
rect 358648 159458 358676 163200
rect 358636 159452 358688 159458
rect 358636 159394 358688 159400
rect 358832 152726 358860 163254
rect 359476 163146 359504 163254
rect 359554 163200 359610 164400
rect 360382 163200 360438 164400
rect 361210 163200 361266 164400
rect 361592 163254 361988 163282
rect 359568 163146 359596 163200
rect 359476 163118 359596 163146
rect 358912 159588 358964 159594
rect 358912 159530 358964 159536
rect 358820 152720 358872 152726
rect 358820 152662 358872 152668
rect 357820 151786 357940 151814
rect 358004 151786 358768 151814
rect 357912 150226 357940 151786
rect 358740 150226 358768 151786
rect 348436 150198 348510 150226
rect 349080 150198 349154 150226
rect 349724 150198 349798 150226
rect 350368 150198 350442 150226
rect 351012 150198 351086 150226
rect 351656 150198 351730 150226
rect 352300 150198 352374 150226
rect 352944 150198 353018 150226
rect 353588 150198 353662 150226
rect 354232 150198 354306 150226
rect 354876 150198 354950 150226
rect 355520 150198 355594 150226
rect 356164 150198 356238 150226
rect 356808 150198 356882 150226
rect 357452 150198 357526 150226
rect 357912 150198 358170 150226
rect 358740 150198 358814 150226
rect 358924 150210 358952 159530
rect 360396 153950 360424 163200
rect 361224 158982 361252 163200
rect 361212 158976 361264 158982
rect 361212 158918 361264 158924
rect 360660 155372 360712 155378
rect 360660 155314 360712 155320
rect 360384 153944 360436 153950
rect 360384 153886 360436 153892
rect 359372 152788 359424 152794
rect 359372 152730 359424 152736
rect 359464 152788 359516 152794
rect 359464 152730 359516 152736
rect 359384 150226 359412 152730
rect 359476 152046 359504 152730
rect 359464 152040 359516 152046
rect 359464 151982 359516 151988
rect 360672 150226 360700 155314
rect 361592 152454 361620 163254
rect 361960 163146 361988 163254
rect 362038 163200 362094 164400
rect 362866 163200 362922 164400
rect 363064 163254 363644 163282
rect 362052 163146 362080 163200
rect 361960 163118 362080 163146
rect 362880 159594 362908 163200
rect 362960 159860 363012 159866
rect 362960 159802 363012 159808
rect 362868 159588 362920 159594
rect 362868 159530 362920 159536
rect 361948 152856 362000 152862
rect 361948 152798 362000 152804
rect 361580 152448 361632 152454
rect 361580 152390 361632 152396
rect 361304 152312 361356 152318
rect 361304 152254 361356 152260
rect 361316 150226 361344 152254
rect 361960 150226 361988 152798
rect 362592 151836 362644 151842
rect 362592 151778 362644 151784
rect 362604 150226 362632 151778
rect 347838 149940 347866 150198
rect 348482 149940 348510 150198
rect 349126 149940 349154 150198
rect 349770 149940 349798 150198
rect 350414 149940 350442 150198
rect 351058 149940 351086 150198
rect 351702 149940 351730 150198
rect 352346 149940 352374 150198
rect 352990 149940 353018 150198
rect 353634 149940 353662 150198
rect 354278 149940 354306 150198
rect 354922 149940 354950 150198
rect 355566 149940 355594 150198
rect 356210 149940 356238 150198
rect 356854 149940 356882 150198
rect 357498 149940 357526 150198
rect 358142 149940 358170 150198
rect 358786 149940 358814 150198
rect 358912 150204 358964 150210
rect 359384 150198 359458 150226
rect 358912 150146 358964 150152
rect 359430 149940 359458 150198
rect 360062 150204 360114 150210
rect 360672 150198 360746 150226
rect 361316 150198 361390 150226
rect 361960 150198 362034 150226
rect 362604 150198 362678 150226
rect 362972 150210 363000 159802
rect 363064 153814 363092 163254
rect 363616 163146 363644 163254
rect 363694 163200 363750 164400
rect 364522 163200 364578 164400
rect 365442 163200 365498 164400
rect 365732 163254 366220 163282
rect 363708 163146 363736 163200
rect 363616 163118 363736 163146
rect 363144 158840 363196 158846
rect 363144 158782 363196 158788
rect 363052 153808 363104 153814
rect 363052 153750 363104 153756
rect 363156 151842 363184 158782
rect 363236 154012 363288 154018
rect 363236 153954 363288 153960
rect 363144 151836 363196 151842
rect 363144 151778 363196 151784
rect 363248 150226 363276 153954
rect 364536 152318 364564 163200
rect 365456 159798 365484 163200
rect 365444 159792 365496 159798
rect 365444 159734 365496 159740
rect 365168 158908 365220 158914
rect 365168 158850 365220 158856
rect 364524 152312 364576 152318
rect 364524 152254 364576 152260
rect 364524 151836 364576 151842
rect 364524 151778 364576 151784
rect 364536 150226 364564 151778
rect 365180 150226 365208 158850
rect 365732 152862 365760 163254
rect 366192 163146 366220 163254
rect 366270 163200 366326 164400
rect 367098 163200 367154 164400
rect 367926 163200 367982 164400
rect 368492 163254 368704 163282
rect 366284 163146 366312 163200
rect 366192 163118 366312 163146
rect 367112 155242 367140 163200
rect 367940 158914 367968 163200
rect 367928 158908 367980 158914
rect 367928 158850 367980 158856
rect 367192 158772 367244 158778
rect 367192 158714 367244 158720
rect 367100 155236 367152 155242
rect 367100 155178 367152 155184
rect 365812 154080 365864 154086
rect 365812 154022 365864 154028
rect 365720 152856 365772 152862
rect 365720 152798 365772 152804
rect 365824 150226 365852 154022
rect 366364 153128 366416 153134
rect 366364 153070 366416 153076
rect 360062 150146 360114 150152
rect 360074 149940 360102 150146
rect 360718 149940 360746 150198
rect 361362 149940 361390 150198
rect 362006 149940 362034 150198
rect 362650 149940 362678 150198
rect 362960 150204 363012 150210
rect 363248 150198 363322 150226
rect 362960 150146 363012 150152
rect 363294 149940 363322 150198
rect 363926 150204 363978 150210
rect 364536 150198 364610 150226
rect 365180 150198 365254 150226
rect 363926 150146 363978 150152
rect 363938 149940 363966 150146
rect 364582 149940 364610 150198
rect 365226 149940 365254 150198
rect 365778 150198 365852 150226
rect 366376 150226 366404 153070
rect 367204 152862 367232 158714
rect 368296 154148 368348 154154
rect 368296 154090 368348 154096
rect 367008 152856 367060 152862
rect 367008 152798 367060 152804
rect 367192 152856 367244 152862
rect 367192 152798 367244 152804
rect 367020 152402 367048 152798
rect 367020 152374 367140 152402
rect 367112 152250 367140 152374
rect 367008 152244 367060 152250
rect 367008 152186 367060 152192
rect 367100 152244 367152 152250
rect 367100 152186 367152 152192
rect 367020 150226 367048 152186
rect 367652 151972 367704 151978
rect 367652 151914 367704 151920
rect 367664 150226 367692 151914
rect 368308 150226 368336 154090
rect 368492 153134 368520 163254
rect 368676 163146 368704 163254
rect 368754 163200 368810 164400
rect 369582 163200 369638 164400
rect 369964 163254 370360 163282
rect 368768 163146 368796 163200
rect 368676 163118 368796 163146
rect 369492 159928 369544 159934
rect 369492 159870 369544 159876
rect 369216 159724 369268 159730
rect 369216 159666 369268 159672
rect 369228 158982 369256 159666
rect 369216 158976 369268 158982
rect 369216 158918 369268 158924
rect 368480 153128 368532 153134
rect 368480 153070 368532 153076
rect 368940 152856 368992 152862
rect 368940 152798 368992 152804
rect 369032 152856 369084 152862
rect 369032 152798 369084 152804
rect 368952 150226 368980 152798
rect 369044 152318 369072 152798
rect 369032 152312 369084 152318
rect 369032 152254 369084 152260
rect 369504 151814 369532 159870
rect 369596 159730 369624 163200
rect 369860 159996 369912 160002
rect 369860 159938 369912 159944
rect 369584 159724 369636 159730
rect 369584 159666 369636 159672
rect 369872 151814 369900 159938
rect 369964 154018 369992 163254
rect 370332 163146 370360 163254
rect 370410 163200 370466 164400
rect 371330 163200 371386 164400
rect 372158 163200 372214 164400
rect 372632 163254 372936 163282
rect 370424 163146 370452 163200
rect 370332 163118 370452 163146
rect 370872 155440 370924 155446
rect 370872 155382 370924 155388
rect 369952 154012 370004 154018
rect 369952 153954 370004 153960
rect 369504 151786 369624 151814
rect 369872 151786 370268 151814
rect 369596 150226 369624 151786
rect 370240 150226 370268 151786
rect 370884 150226 370912 155382
rect 371344 152250 371372 163200
rect 372172 160002 372200 163200
rect 372160 159996 372212 160002
rect 372160 159938 372212 159944
rect 372632 152998 372660 163254
rect 372908 163146 372936 163254
rect 372986 163200 373042 164400
rect 373814 163200 373870 164400
rect 374642 163200 374698 164400
rect 375470 163200 375526 164400
rect 376298 163200 376354 164400
rect 376864 163254 377168 163282
rect 373000 163146 373028 163200
rect 372908 163118 373028 163146
rect 373448 155508 373500 155514
rect 373448 155450 373500 155456
rect 371516 152992 371568 152998
rect 371516 152934 371568 152940
rect 372620 152992 372672 152998
rect 372620 152934 372672 152940
rect 371332 152244 371384 152250
rect 371332 152186 371384 152192
rect 371528 150226 371556 152934
rect 372804 152176 372856 152182
rect 372804 152118 372856 152124
rect 372160 151904 372212 151910
rect 372160 151846 372212 151852
rect 372172 150226 372200 151846
rect 372816 150226 372844 152118
rect 373460 150226 373488 155450
rect 373828 155310 373856 163200
rect 374000 160064 374052 160070
rect 374000 160006 374052 160012
rect 373816 155304 373868 155310
rect 373816 155246 373868 155252
rect 366376 150198 366450 150226
rect 367020 150198 367094 150226
rect 367664 150198 367738 150226
rect 368308 150198 368382 150226
rect 368952 150198 369026 150226
rect 369596 150198 369670 150226
rect 370240 150198 370314 150226
rect 370884 150198 370958 150226
rect 371528 150198 371602 150226
rect 372172 150198 372246 150226
rect 372816 150198 372890 150226
rect 373460 150198 373534 150226
rect 374012 150210 374040 160006
rect 374092 159316 374144 159322
rect 374092 159258 374144 159264
rect 374104 150226 374132 159258
rect 374656 158778 374684 163200
rect 374644 158772 374696 158778
rect 374644 158714 374696 158720
rect 375380 152108 375432 152114
rect 375380 152050 375432 152056
rect 375392 150226 375420 152050
rect 375484 151978 375512 163200
rect 376312 159866 376340 163200
rect 376300 159860 376352 159866
rect 376300 159802 376352 159808
rect 376668 156664 376720 156670
rect 376668 156606 376720 156612
rect 376024 154284 376076 154290
rect 376024 154226 376076 154232
rect 375472 151972 375524 151978
rect 375472 151914 375524 151920
rect 376036 150226 376064 154226
rect 376680 150226 376708 156606
rect 376864 154086 376892 163254
rect 377140 163146 377168 163254
rect 377218 163200 377274 164400
rect 378046 163200 378102 164400
rect 378874 163200 378930 164400
rect 379702 163200 379758 164400
rect 380176 163254 380480 163282
rect 377232 163146 377260 163200
rect 377140 163118 377260 163146
rect 378060 159322 378088 163200
rect 378888 160070 378916 163200
rect 378876 160064 378928 160070
rect 378876 160006 378928 160012
rect 379716 159934 379744 163200
rect 379704 159928 379756 159934
rect 379704 159870 379756 159876
rect 378048 159316 378100 159322
rect 378048 159258 378100 159264
rect 377956 159248 378008 159254
rect 377956 159190 378008 159196
rect 376852 154080 376904 154086
rect 376852 154022 376904 154028
rect 377312 152924 377364 152930
rect 377312 152866 377364 152872
rect 377324 150226 377352 152866
rect 377968 150226 377996 159190
rect 378232 159180 378284 159186
rect 378232 159122 378284 159128
rect 378140 155576 378192 155582
rect 378140 155518 378192 155524
rect 365778 149940 365806 150198
rect 366422 149940 366450 150198
rect 367066 149940 367094 150198
rect 367710 149940 367738 150198
rect 368354 149940 368382 150198
rect 368998 149940 369026 150198
rect 369642 149940 369670 150198
rect 370286 149940 370314 150198
rect 370930 149940 370958 150198
rect 371574 149940 371602 150198
rect 372218 149940 372246 150198
rect 372862 149940 372890 150198
rect 373506 149940 373534 150198
rect 374000 150204 374052 150210
rect 374104 150198 374178 150226
rect 374000 150146 374052 150152
rect 374150 149940 374178 150198
rect 374782 150204 374834 150210
rect 375392 150198 375466 150226
rect 376036 150198 376110 150226
rect 376680 150198 376754 150226
rect 377324 150198 377398 150226
rect 377968 150198 378042 150226
rect 378152 150210 378180 155518
rect 378244 152930 378272 159122
rect 378784 159044 378836 159050
rect 378784 158986 378836 158992
rect 378600 153876 378652 153882
rect 378600 153818 378652 153824
rect 378232 152924 378284 152930
rect 378232 152866 378284 152872
rect 378612 150226 378640 153818
rect 378796 152046 378824 158986
rect 380176 153882 380204 163254
rect 380452 163146 380480 163254
rect 380530 163200 380586 164400
rect 380912 163254 381308 163282
rect 380544 163146 380572 163200
rect 380452 163118 380572 163146
rect 380164 153876 380216 153882
rect 380164 153818 380216 153824
rect 380912 152930 380940 163254
rect 381280 163146 381308 163254
rect 381358 163200 381414 164400
rect 381464 163254 382136 163282
rect 381372 163146 381400 163200
rect 381280 163118 381400 163146
rect 381176 154216 381228 154222
rect 381176 154158 381228 154164
rect 379888 152924 379940 152930
rect 379888 152866 379940 152872
rect 380900 152924 380952 152930
rect 380900 152866 380952 152872
rect 378784 152040 378836 152046
rect 378784 151982 378836 151988
rect 379900 150226 379928 152866
rect 380532 152380 380584 152386
rect 380532 152322 380584 152328
rect 380544 150226 380572 152322
rect 381188 150226 381216 154158
rect 381464 152386 381492 163254
rect 382108 163146 382136 163254
rect 382186 163200 382242 164400
rect 383106 163200 383162 164400
rect 383672 163254 383884 163282
rect 382200 163146 382228 163200
rect 382108 163118 382228 163146
rect 383120 159390 383148 163200
rect 382832 159384 382884 159390
rect 382832 159326 382884 159332
rect 383108 159384 383160 159390
rect 383108 159326 383160 159332
rect 382280 159112 382332 159118
rect 382280 159054 382332 159060
rect 381820 156732 381872 156738
rect 381820 156674 381872 156680
rect 381452 152380 381504 152386
rect 381452 152322 381504 152328
rect 381832 150226 381860 156674
rect 382292 152114 382320 159054
rect 382464 152652 382516 152658
rect 382464 152594 382516 152600
rect 382280 152108 382332 152114
rect 382280 152050 382332 152056
rect 382476 150226 382504 152594
rect 382844 151814 382872 159326
rect 383672 154154 383700 163254
rect 383856 163146 383884 163254
rect 383934 163200 383990 164400
rect 384762 163200 384818 164400
rect 385590 163200 385646 164400
rect 386418 163200 386474 164400
rect 386524 163254 387196 163282
rect 383948 163146 383976 163200
rect 383856 163118 383976 163146
rect 384672 159044 384724 159050
rect 384672 158986 384724 158992
rect 384684 158778 384712 158986
rect 384776 158778 384804 163200
rect 385316 159656 385368 159662
rect 385316 159598 385368 159604
rect 384948 158976 385000 158982
rect 384948 158918 385000 158924
rect 384672 158772 384724 158778
rect 384672 158714 384724 158720
rect 384764 158772 384816 158778
rect 384764 158714 384816 158720
rect 383752 154352 383804 154358
rect 383752 154294 383804 154300
rect 383660 154148 383712 154154
rect 383660 154090 383712 154096
rect 382844 151786 383148 151814
rect 383120 150226 383148 151786
rect 383764 150226 383792 154294
rect 384960 152182 384988 158918
rect 385328 152522 385356 159598
rect 385604 159254 385632 163200
rect 385592 159248 385644 159254
rect 385592 159190 385644 159196
rect 386236 158908 386288 158914
rect 386236 158850 386288 158856
rect 385776 158840 385828 158846
rect 385776 158782 385828 158788
rect 385592 153060 385644 153066
rect 385592 153002 385644 153008
rect 385040 152516 385092 152522
rect 385040 152458 385092 152464
rect 385316 152516 385368 152522
rect 385316 152458 385368 152464
rect 384948 152176 385000 152182
rect 384948 152118 385000 152124
rect 384396 152040 384448 152046
rect 384396 151982 384448 151988
rect 384408 150226 384436 151982
rect 385052 150226 385080 152458
rect 385604 151814 385632 153002
rect 385788 152046 385816 158782
rect 386248 153066 386276 158850
rect 386328 154420 386380 154426
rect 386328 154362 386380 154368
rect 386236 153060 386288 153066
rect 386236 153002 386288 153008
rect 385776 152040 385828 152046
rect 385776 151982 385828 151988
rect 385604 151786 385724 151814
rect 385696 150226 385724 151786
rect 386340 150226 386368 154362
rect 386432 152658 386460 163200
rect 386524 154222 386552 163254
rect 387168 163146 387196 163254
rect 387246 163200 387302 164400
rect 388074 163200 388130 164400
rect 388994 163200 389050 164400
rect 389822 163200 389878 164400
rect 390650 163200 390706 164400
rect 391478 163200 391534 164400
rect 392306 163200 392362 164400
rect 393134 163200 393190 164400
rect 393332 163254 393912 163282
rect 387260 163146 387288 163200
rect 387168 163118 387288 163146
rect 388088 158846 388116 163200
rect 388352 159316 388404 159322
rect 388352 159258 388404 159264
rect 388076 158840 388128 158846
rect 388076 158782 388128 158788
rect 386512 154216 386564 154222
rect 386512 154158 386564 154164
rect 388260 153196 388312 153202
rect 388260 153138 388312 153144
rect 386420 152652 386472 152658
rect 386420 152594 386472 152600
rect 387616 152516 387668 152522
rect 387616 152458 387668 152464
rect 386972 152108 387024 152114
rect 386972 152050 387024 152056
rect 386984 150226 387012 152050
rect 387628 150226 387656 152458
rect 388272 150226 388300 153138
rect 388364 152114 388392 159258
rect 389008 159050 389036 163200
rect 389836 159662 389864 163200
rect 389824 159656 389876 159662
rect 389824 159598 389876 159604
rect 390560 159520 390612 159526
rect 390560 159462 390612 159468
rect 388444 159044 388496 159050
rect 388444 158986 388496 158992
rect 388996 159044 389048 159050
rect 388996 158986 389048 158992
rect 388352 152108 388404 152114
rect 388352 152050 388404 152056
rect 388456 151842 388484 158986
rect 390376 158840 390428 158846
rect 390376 158782 390428 158788
rect 389180 158772 389232 158778
rect 389180 158714 389232 158720
rect 388904 154556 388956 154562
rect 388904 154498 388956 154504
rect 388444 151836 388496 151842
rect 388444 151778 388496 151784
rect 388916 150226 388944 154498
rect 389192 153202 389220 158714
rect 389180 153196 389232 153202
rect 389180 153138 389232 153144
rect 390192 152788 390244 152794
rect 390192 152730 390244 152736
rect 389548 152584 389600 152590
rect 389548 152526 389600 152532
rect 389560 150226 389588 152526
rect 390204 150226 390232 152730
rect 390388 152658 390416 158782
rect 390376 152652 390428 152658
rect 390376 152594 390428 152600
rect 390572 151814 390600 159462
rect 390664 154358 390692 163200
rect 391492 158914 391520 163200
rect 392320 159526 392348 163200
rect 392308 159520 392360 159526
rect 392308 159462 392360 159468
rect 392768 159452 392820 159458
rect 392768 159394 392820 159400
rect 391480 158908 391532 158914
rect 391480 158850 391532 158856
rect 391480 154488 391532 154494
rect 391480 154430 391532 154436
rect 390652 154352 390704 154358
rect 390652 154294 390704 154300
rect 390572 151786 390876 151814
rect 390848 150226 390876 151786
rect 391492 150226 391520 154430
rect 392124 152176 392176 152182
rect 392124 152118 392176 152124
rect 392136 150226 392164 152118
rect 392780 150226 392808 159394
rect 393148 152522 393176 163200
rect 393332 154290 393360 163254
rect 393884 163146 393912 163254
rect 393962 163200 394018 164400
rect 394882 163200 394938 164400
rect 395710 163200 395766 164400
rect 396538 163200 396594 164400
rect 397366 163200 397422 164400
rect 397472 163254 398144 163282
rect 393976 163146 394004 163200
rect 393884 163118 394004 163146
rect 394332 158908 394384 158914
rect 394332 158850 394384 158856
rect 393320 154284 393372 154290
rect 393320 154226 393372 154232
rect 394056 153944 394108 153950
rect 394056 153886 394108 153892
rect 393412 152720 393464 152726
rect 393412 152662 393464 152668
rect 393136 152516 393188 152522
rect 393136 152458 393188 152464
rect 393424 150226 393452 152662
rect 394068 150226 394096 153886
rect 394344 152182 394372 158850
rect 394896 152590 394924 163200
rect 395528 159792 395580 159798
rect 395528 159734 395580 159740
rect 395540 152726 395568 159734
rect 395724 159322 395752 163200
rect 396172 159996 396224 160002
rect 396172 159938 396224 159944
rect 395988 159588 396040 159594
rect 395988 159530 396040 159536
rect 395712 159316 395764 159322
rect 395712 159258 395764 159264
rect 395528 152720 395580 152726
rect 395528 152662 395580 152668
rect 394884 152584 394936 152590
rect 394884 152526 394936 152532
rect 395344 152448 395396 152454
rect 395344 152390 395396 152396
rect 394332 152176 394384 152182
rect 394332 152118 394384 152124
rect 394700 152040 394752 152046
rect 394700 151982 394752 151988
rect 394712 150226 394740 151982
rect 395356 150226 395384 152390
rect 396000 150226 396028 159530
rect 396184 151910 396212 159938
rect 396552 159798 396580 163200
rect 396540 159792 396592 159798
rect 396540 159734 396592 159740
rect 397380 153950 397408 163200
rect 397472 154426 397500 163254
rect 398116 163146 398144 163254
rect 398194 163200 398250 164400
rect 399022 163200 399078 164400
rect 399128 163254 399800 163282
rect 398208 163146 398236 163200
rect 398116 163118 398236 163146
rect 398564 160064 398616 160070
rect 398564 160006 398616 160012
rect 397460 154420 397512 154426
rect 397460 154362 397512 154368
rect 397368 153944 397420 153950
rect 397368 153886 397420 153892
rect 396540 153808 396592 153814
rect 396540 153750 396592 153756
rect 396172 151904 396224 151910
rect 396172 151846 396224 151852
rect 396552 150226 396580 153750
rect 397184 152856 397236 152862
rect 397184 152798 397236 152804
rect 397196 150226 397224 152798
rect 397828 152720 397880 152726
rect 397828 152662 397880 152668
rect 397840 150226 397868 152662
rect 398576 152318 398604 160006
rect 399036 160002 399064 163200
rect 399024 159996 399076 160002
rect 399024 159938 399076 159944
rect 398840 159248 398892 159254
rect 398840 159190 398892 159196
rect 398852 152454 398880 159190
rect 399024 155236 399076 155242
rect 399024 155178 399076 155184
rect 398840 152448 398892 152454
rect 398840 152390 398892 152396
rect 398472 152312 398524 152318
rect 398472 152254 398524 152260
rect 398564 152312 398616 152318
rect 398564 152254 398616 152260
rect 398484 150226 398512 152254
rect 399036 151814 399064 155178
rect 399128 152726 399156 163254
rect 399772 163146 399800 163254
rect 399850 163200 399906 164400
rect 400324 163254 400720 163282
rect 399864 163146 399892 163200
rect 399772 163118 399892 163146
rect 400324 154494 400352 163254
rect 400692 163146 400720 163254
rect 400770 163200 400826 164400
rect 401598 163200 401654 164400
rect 401704 163254 402376 163282
rect 400784 163146 400812 163200
rect 400692 163118 400812 163146
rect 401048 159724 401100 159730
rect 401048 159666 401100 159672
rect 400312 154488 400364 154494
rect 400312 154430 400364 154436
rect 400404 153128 400456 153134
rect 400404 153070 400456 153076
rect 399760 153060 399812 153066
rect 399760 153002 399812 153008
rect 399116 152720 399168 152726
rect 399116 152662 399168 152668
rect 399036 151786 399156 151814
rect 399128 150226 399156 151786
rect 399772 150226 399800 153002
rect 400416 150226 400444 153070
rect 401060 150226 401088 159666
rect 401612 155242 401640 163200
rect 401600 155236 401652 155242
rect 401600 155178 401652 155184
rect 401600 154012 401652 154018
rect 401600 153954 401652 153960
rect 401612 151814 401640 153954
rect 401704 152862 401732 163254
rect 402348 163146 402376 163254
rect 402426 163200 402482 164400
rect 403254 163200 403310 164400
rect 404082 163200 404138 164400
rect 404372 163254 404860 163282
rect 402440 163146 402468 163200
rect 402348 163118 402468 163146
rect 403268 159730 403296 163200
rect 403256 159724 403308 159730
rect 403256 159666 403308 159672
rect 404096 159458 404124 163200
rect 404268 159520 404320 159526
rect 404268 159462 404320 159468
rect 404084 159452 404136 159458
rect 404084 159394 404136 159400
rect 403256 159044 403308 159050
rect 403256 158986 403308 158992
rect 403164 155304 403216 155310
rect 403164 155246 403216 155252
rect 401692 152856 401744 152862
rect 401692 152798 401744 152804
rect 402336 152244 402388 152250
rect 402336 152186 402388 152192
rect 401612 151786 401732 151814
rect 401704 150226 401732 151786
rect 402348 150226 402376 152186
rect 402980 151904 403032 151910
rect 402980 151846 403032 151852
rect 402992 150226 403020 151846
rect 374782 150146 374834 150152
rect 374794 149940 374822 150146
rect 375438 149940 375466 150198
rect 376082 149940 376110 150198
rect 376726 149940 376754 150198
rect 377370 149940 377398 150198
rect 378014 149940 378042 150198
rect 378140 150204 378192 150210
rect 378612 150198 378686 150226
rect 378140 150146 378192 150152
rect 378658 149940 378686 150198
rect 379290 150204 379342 150210
rect 379900 150198 379974 150226
rect 380544 150198 380618 150226
rect 381188 150198 381262 150226
rect 381832 150198 381906 150226
rect 382476 150198 382550 150226
rect 383120 150198 383194 150226
rect 383764 150198 383838 150226
rect 384408 150198 384482 150226
rect 385052 150198 385126 150226
rect 385696 150198 385770 150226
rect 386340 150198 386414 150226
rect 386984 150198 387058 150226
rect 387628 150198 387702 150226
rect 388272 150198 388346 150226
rect 388916 150198 388990 150226
rect 389560 150198 389634 150226
rect 390204 150198 390278 150226
rect 390848 150198 390922 150226
rect 391492 150198 391566 150226
rect 392136 150198 392210 150226
rect 392780 150198 392854 150226
rect 393424 150198 393498 150226
rect 394068 150198 394142 150226
rect 394712 150198 394786 150226
rect 395356 150198 395430 150226
rect 396000 150198 396074 150226
rect 396552 150198 396626 150226
rect 397196 150198 397270 150226
rect 397840 150198 397914 150226
rect 398484 150198 398558 150226
rect 399128 150198 399202 150226
rect 399772 150198 399846 150226
rect 400416 150198 400490 150226
rect 401060 150198 401134 150226
rect 401704 150198 401778 150226
rect 402348 150198 402422 150226
rect 402992 150198 403066 150226
rect 403176 150210 403204 155246
rect 403268 153134 403296 158986
rect 403256 153128 403308 153134
rect 403256 153070 403308 153076
rect 403624 152992 403676 152998
rect 403624 152934 403676 152940
rect 403636 150226 403664 152934
rect 404280 151910 404308 159462
rect 404372 152998 404400 163254
rect 404832 163146 404860 163254
rect 404910 163200 404966 164400
rect 405738 163200 405794 164400
rect 406658 163200 406714 164400
rect 407486 163200 407542 164400
rect 407684 163254 408264 163282
rect 404924 163146 404952 163200
rect 404832 163118 404952 163146
rect 404728 159316 404780 159322
rect 404728 159258 404780 159264
rect 404360 152992 404412 152998
rect 404360 152934 404412 152940
rect 404740 152046 404768 159258
rect 405752 158846 405780 163200
rect 405832 159928 405884 159934
rect 405832 159870 405884 159876
rect 405740 158840 405792 158846
rect 405740 158782 405792 158788
rect 405844 152250 405872 159870
rect 406200 159860 406252 159866
rect 406200 159802 406252 159808
rect 405832 152244 405884 152250
rect 405832 152186 405884 152192
rect 404728 152040 404780 152046
rect 404728 151982 404780 151988
rect 405556 151972 405608 151978
rect 405556 151914 405608 151920
rect 404268 151904 404320 151910
rect 404268 151846 404320 151852
rect 404912 151836 404964 151842
rect 404912 151778 404964 151784
rect 404924 150226 404952 151778
rect 405568 150226 405596 151914
rect 406212 150226 406240 159802
rect 406672 153066 406700 163200
rect 407500 159594 407528 163200
rect 407488 159588 407540 159594
rect 407488 159530 407540 159536
rect 406844 154080 406896 154086
rect 406844 154022 406896 154028
rect 406660 153060 406712 153066
rect 406660 153002 406712 153008
rect 406856 150226 406884 154022
rect 407684 152425 407712 163254
rect 408236 163146 408264 163254
rect 408314 163200 408370 164400
rect 409142 163200 409198 164400
rect 409970 163200 410026 164400
rect 410798 163200 410854 164400
rect 411272 163254 411576 163282
rect 408328 163146 408356 163200
rect 408236 163118 408356 163146
rect 408500 159996 408552 160002
rect 408500 159938 408552 159944
rect 407670 152416 407726 152425
rect 407670 152351 407726 152360
rect 408132 152312 408184 152318
rect 408132 152254 408184 152260
rect 407488 152108 407540 152114
rect 407488 152050 407540 152056
rect 407500 150226 407528 152050
rect 408144 150226 408172 152254
rect 408512 152114 408540 159938
rect 409156 159118 409184 163200
rect 409984 159866 410012 163200
rect 409972 159860 410024 159866
rect 409972 159802 410024 159808
rect 410812 159526 410840 163200
rect 410800 159520 410852 159526
rect 410800 159462 410852 159468
rect 409144 159112 409196 159118
rect 409144 159054 409196 159060
rect 410892 159112 410944 159118
rect 410892 159054 410944 159060
rect 409236 158840 409288 158846
rect 409236 158782 409288 158788
rect 409248 152250 409276 158782
rect 409420 153876 409472 153882
rect 409420 153818 409472 153824
rect 408776 152244 408828 152250
rect 408776 152186 408828 152192
rect 409236 152244 409288 152250
rect 409236 152186 409288 152192
rect 408500 152108 408552 152114
rect 408500 152050 408552 152056
rect 408788 150226 408816 152186
rect 409432 150226 409460 153818
rect 410064 152924 410116 152930
rect 410064 152866 410116 152872
rect 410076 150226 410104 152866
rect 410708 152380 410760 152386
rect 410708 152322 410760 152328
rect 410720 150226 410748 152322
rect 410904 152318 410932 159054
rect 411272 152930 411300 163254
rect 411548 163146 411576 163254
rect 411626 163200 411682 164400
rect 412546 163200 412602 164400
rect 413374 163200 413430 164400
rect 414202 163200 414258 164400
rect 414400 163254 414980 163282
rect 411640 163146 411668 163200
rect 411548 163118 411668 163146
rect 411352 159384 411404 159390
rect 411352 159326 411404 159332
rect 411260 152924 411312 152930
rect 411260 152866 411312 152872
rect 410892 152312 410944 152318
rect 410892 152254 410944 152260
rect 411364 150226 411392 159326
rect 412560 158914 412588 163200
rect 413192 159792 413244 159798
rect 413192 159734 413244 159740
rect 412548 158908 412600 158914
rect 412548 158850 412600 158856
rect 413100 158908 413152 158914
rect 413100 158850 413152 158856
rect 411996 154148 412048 154154
rect 411996 154090 412048 154096
rect 412008 150226 412036 154090
rect 413112 153202 413140 158850
rect 412640 153196 412692 153202
rect 412640 153138 412692 153144
rect 413100 153196 413152 153202
rect 413100 153138 413152 153144
rect 412652 150226 412680 153138
rect 413204 152386 413232 159734
rect 413388 158846 413416 163200
rect 413836 159656 413888 159662
rect 413836 159598 413888 159604
rect 413376 158840 413428 158846
rect 413376 158782 413428 158788
rect 413848 152454 413876 159598
rect 414216 159390 414244 163200
rect 414204 159384 414256 159390
rect 414204 159326 414256 159332
rect 414400 152658 414428 163254
rect 414952 163146 414980 163254
rect 415030 163200 415086 164400
rect 415412 163254 415808 163282
rect 415044 163146 415072 163200
rect 414952 163118 415072 163146
rect 414572 154216 414624 154222
rect 414572 154158 414624 154164
rect 413928 152652 413980 152658
rect 413928 152594 413980 152600
rect 414388 152652 414440 152658
rect 414388 152594 414440 152600
rect 413284 152448 413336 152454
rect 413284 152390 413336 152396
rect 413836 152448 413888 152454
rect 413836 152390 413888 152396
rect 413192 152380 413244 152386
rect 413192 152322 413244 152328
rect 413296 150226 413324 152390
rect 413940 150226 413968 152594
rect 414584 150226 414612 154158
rect 415412 152794 415440 163254
rect 415780 163146 415808 163254
rect 415858 163200 415914 164400
rect 416686 163200 416742 164400
rect 417514 163200 417570 164400
rect 418434 163200 418490 164400
rect 419262 163200 419318 164400
rect 420090 163200 420146 164400
rect 420918 163200 420974 164400
rect 421208 163254 421696 163282
rect 415872 163146 415900 163200
rect 415780 163118 415900 163146
rect 416596 159724 416648 159730
rect 416596 159666 416648 159672
rect 415860 153128 415912 153134
rect 415860 153070 415912 153076
rect 415216 152788 415268 152794
rect 415216 152730 415268 152736
rect 415400 152788 415452 152794
rect 415400 152730 415452 152736
rect 415228 150226 415256 152730
rect 415872 150226 415900 153070
rect 416504 152448 416556 152454
rect 416504 152390 416556 152396
rect 416516 150226 416544 152390
rect 416608 151978 416636 159666
rect 416700 158778 416728 163200
rect 417424 159860 417476 159866
rect 417424 159802 417476 159808
rect 416688 158772 416740 158778
rect 416688 158714 416740 158720
rect 417148 154352 417200 154358
rect 417148 154294 417200 154300
rect 416596 151972 416648 151978
rect 416596 151914 416648 151920
rect 417160 150226 417188 154294
rect 417436 151842 417464 159802
rect 417528 159662 417556 163200
rect 417516 159656 417568 159662
rect 417516 159598 417568 159604
rect 418448 152454 418476 163200
rect 419276 153134 419304 163200
rect 420104 158982 420132 163200
rect 420932 159730 420960 163200
rect 420920 159724 420972 159730
rect 420920 159666 420972 159672
rect 420092 158976 420144 158982
rect 420092 158918 420144 158924
rect 419632 158840 419684 158846
rect 419632 158782 419684 158788
rect 419540 158772 419592 158778
rect 419540 158714 419592 158720
rect 419264 153128 419316 153134
rect 419264 153070 419316 153076
rect 419080 152516 419132 152522
rect 419080 152458 419132 152464
rect 418436 152448 418488 152454
rect 418436 152390 418488 152396
rect 417792 152176 417844 152182
rect 417792 152118 417844 152124
rect 417424 151836 417476 151842
rect 417424 151778 417476 151784
rect 417804 150226 417832 152118
rect 418436 151904 418488 151910
rect 418436 151846 418488 151852
rect 418448 150226 418476 151846
rect 419092 150226 419120 152458
rect 419552 151910 419580 158714
rect 419644 152182 419672 158782
rect 419724 154284 419776 154290
rect 419724 154226 419776 154232
rect 419632 152176 419684 152182
rect 419632 152118 419684 152124
rect 419540 151904 419592 151910
rect 419540 151846 419592 151852
rect 419736 150226 419764 154226
rect 420368 152584 420420 152590
rect 420368 152526 420420 152532
rect 420380 150226 420408 152526
rect 421208 152522 421236 163254
rect 421668 163146 421696 163254
rect 421746 163200 421802 164400
rect 422574 163200 422630 164400
rect 423402 163200 423458 164400
rect 424322 163200 424378 164400
rect 425150 163200 425206 164400
rect 425978 163200 426034 164400
rect 426452 163254 426756 163282
rect 421760 163146 421788 163200
rect 421668 163118 421788 163146
rect 422484 153944 422536 153950
rect 422484 153886 422536 153892
rect 421196 152516 421248 152522
rect 421196 152458 421248 152464
rect 421656 152380 421708 152386
rect 421656 152322 421708 152328
rect 421012 152040 421064 152046
rect 421012 151982 421064 151988
rect 421024 150226 421052 151982
rect 421668 150226 421696 152322
rect 422496 151814 422524 153886
rect 422588 151978 422616 163200
rect 423036 154420 423088 154426
rect 423036 154362 423088 154368
rect 422576 151972 422628 151978
rect 422576 151914 422628 151920
rect 422404 151786 422524 151814
rect 422404 150226 422432 151786
rect 423048 150226 423076 154362
rect 423416 152590 423444 163200
rect 424336 159798 424364 163200
rect 424324 159792 424376 159798
rect 424324 159734 424376 159740
rect 423588 158976 423640 158982
rect 423588 158918 423640 158924
rect 423404 152584 423456 152590
rect 423404 152526 423456 152532
rect 423600 152266 423628 158918
rect 424876 154488 424928 154494
rect 424876 154430 424928 154436
rect 424232 152720 424284 152726
rect 424232 152662 424284 152668
rect 423600 152238 423720 152266
rect 423692 152114 423720 152238
rect 423588 152108 423640 152114
rect 423588 152050 423640 152056
rect 423680 152108 423732 152114
rect 423680 152050 423732 152056
rect 379290 150146 379342 150152
rect 379302 149940 379330 150146
rect 379946 149940 379974 150198
rect 380590 149940 380618 150198
rect 381234 149940 381262 150198
rect 381878 149940 381906 150198
rect 382522 149940 382550 150198
rect 383166 149940 383194 150198
rect 383810 149940 383838 150198
rect 384454 149940 384482 150198
rect 385098 149940 385126 150198
rect 385742 149940 385770 150198
rect 386386 149940 386414 150198
rect 387030 149940 387058 150198
rect 387674 149940 387702 150198
rect 388318 149940 388346 150198
rect 388962 149940 388990 150198
rect 389606 149940 389634 150198
rect 390250 149940 390278 150198
rect 390894 149940 390922 150198
rect 391538 149940 391566 150198
rect 392182 149940 392210 150198
rect 392826 149940 392854 150198
rect 393470 149940 393498 150198
rect 394114 149940 394142 150198
rect 394758 149940 394786 150198
rect 395402 149940 395430 150198
rect 396046 149940 396074 150198
rect 396598 149940 396626 150198
rect 397242 149940 397270 150198
rect 397886 149940 397914 150198
rect 398530 149940 398558 150198
rect 399174 149940 399202 150198
rect 399818 149940 399846 150198
rect 400462 149940 400490 150198
rect 401106 149940 401134 150198
rect 401750 149940 401778 150198
rect 402394 149940 402422 150198
rect 403038 149940 403066 150198
rect 403164 150204 403216 150210
rect 403636 150198 403710 150226
rect 403164 150146 403216 150152
rect 403682 149940 403710 150198
rect 404314 150204 404366 150210
rect 404924 150198 404998 150226
rect 405568 150198 405642 150226
rect 406212 150198 406286 150226
rect 406856 150198 406930 150226
rect 407500 150198 407574 150226
rect 408144 150198 408218 150226
rect 408788 150198 408862 150226
rect 409432 150198 409506 150226
rect 410076 150198 410150 150226
rect 410720 150198 410794 150226
rect 411364 150198 411438 150226
rect 412008 150198 412082 150226
rect 412652 150198 412726 150226
rect 413296 150198 413370 150226
rect 413940 150198 414014 150226
rect 414584 150198 414658 150226
rect 415228 150198 415302 150226
rect 415872 150198 415946 150226
rect 416516 150198 416590 150226
rect 417160 150198 417234 150226
rect 417804 150198 417878 150226
rect 418448 150198 418522 150226
rect 419092 150198 419166 150226
rect 419736 150198 419810 150226
rect 420380 150198 420454 150226
rect 421024 150198 421098 150226
rect 421668 150198 421742 150226
rect 404314 150146 404366 150152
rect 404326 149940 404354 150146
rect 404970 149940 404998 150198
rect 405614 149940 405642 150198
rect 406258 149940 406286 150198
rect 406902 149940 406930 150198
rect 407546 149940 407574 150198
rect 408190 149940 408218 150198
rect 408834 149940 408862 150198
rect 409478 149940 409506 150198
rect 410122 149940 410150 150198
rect 410766 149940 410794 150198
rect 411410 149940 411438 150198
rect 412054 149940 412082 150198
rect 412698 149940 412726 150198
rect 413342 149940 413370 150198
rect 413986 149940 414014 150198
rect 414630 149940 414658 150198
rect 415274 149940 415302 150198
rect 415918 149940 415946 150198
rect 416562 149940 416590 150198
rect 417206 149940 417234 150198
rect 417850 149940 417878 150198
rect 418494 149940 418522 150198
rect 419138 149940 419166 150198
rect 419782 149940 419810 150198
rect 420426 149940 420454 150198
rect 421070 149940 421098 150198
rect 421714 149940 421742 150198
rect 422358 150198 422432 150226
rect 423002 150198 423076 150226
rect 423600 150226 423628 152050
rect 424244 150226 424272 152662
rect 424888 150226 424916 154430
rect 425164 152386 425192 163200
rect 425520 155236 425572 155242
rect 425520 155178 425572 155184
rect 425152 152380 425204 152386
rect 425152 152322 425204 152328
rect 425532 150226 425560 155178
rect 425992 153338 426020 163200
rect 426452 153814 426480 163254
rect 426728 163146 426756 163254
rect 426806 163200 426862 164400
rect 427634 163200 427690 164400
rect 427832 163254 428412 163282
rect 426820 163146 426848 163200
rect 426728 163118 426848 163146
rect 427648 159458 427676 163200
rect 427360 159452 427412 159458
rect 427360 159394 427412 159400
rect 427636 159452 427688 159458
rect 427636 159394 427688 159400
rect 426440 153808 426492 153814
rect 426440 153750 426492 153756
rect 425980 153332 426032 153338
rect 425980 153274 426032 153280
rect 426164 152856 426216 152862
rect 426164 152798 426216 152804
rect 426348 152856 426400 152862
rect 426348 152798 426400 152804
rect 426176 150226 426204 152798
rect 426360 152114 426388 152798
rect 426716 152244 426768 152250
rect 426716 152186 426768 152192
rect 426348 152108 426400 152114
rect 426348 152050 426400 152056
rect 423600 150198 423674 150226
rect 424244 150198 424318 150226
rect 424888 150198 424962 150226
rect 425532 150198 425606 150226
rect 426176 150198 426250 150226
rect 426728 150210 426756 152186
rect 426808 152040 426860 152046
rect 426808 151982 426860 151988
rect 426820 150226 426848 151982
rect 427372 150226 427400 159394
rect 427832 157334 427860 163254
rect 428384 163146 428412 163254
rect 428462 163200 428518 164400
rect 429290 163200 429346 164400
rect 430210 163200 430266 164400
rect 430592 163254 430988 163282
rect 428476 163146 428504 163200
rect 428384 163118 428504 163146
rect 429304 157334 429332 163200
rect 429936 159588 429988 159594
rect 429936 159530 429988 159536
rect 427832 157306 428228 157334
rect 429304 157306 429424 157334
rect 428096 153264 428148 153270
rect 428096 153206 428148 153212
rect 427912 153196 427964 153202
rect 427832 153156 427912 153184
rect 427636 152992 427688 152998
rect 427636 152934 427688 152940
rect 427648 150249 427676 152934
rect 427832 152794 427860 153156
rect 427912 153138 427964 153144
rect 428108 152998 428136 153206
rect 428096 152992 428148 152998
rect 428096 152934 428148 152940
rect 427820 152788 427872 152794
rect 427820 152730 427872 152736
rect 428200 152726 428228 157306
rect 429292 153060 429344 153066
rect 429292 153002 429344 153008
rect 428188 152720 428240 152726
rect 428188 152662 428240 152668
rect 427728 152176 427780 152182
rect 427728 152118 427780 152124
rect 427634 150240 427690 150249
rect 422358 149940 422386 150198
rect 423002 149940 423030 150198
rect 423646 149940 423674 150198
rect 424290 149940 424318 150198
rect 424934 149940 424962 150198
rect 425578 149940 425606 150198
rect 426222 149940 426250 150198
rect 426716 150204 426768 150210
rect 426820 150198 426894 150226
rect 427372 150198 427446 150226
rect 426716 150146 426768 150152
rect 426866 149940 426894 150198
rect 427418 149940 427446 150198
rect 427634 150175 427690 150184
rect 427740 150142 427768 152118
rect 428048 150240 428104 150249
rect 428048 150175 428104 150184
rect 428694 150204 428746 150210
rect 427728 150136 427780 150142
rect 427728 150078 427780 150084
rect 428062 149940 428090 150175
rect 428694 150146 428746 150152
rect 428706 149940 428734 150146
rect 429304 150090 429332 153002
rect 429396 152250 429424 157306
rect 429844 152584 429896 152590
rect 429844 152526 429896 152532
rect 429384 152244 429436 152250
rect 429384 152186 429436 152192
rect 429856 151978 429884 152526
rect 429844 151972 429896 151978
rect 429844 151914 429896 151920
rect 429948 150226 429976 159530
rect 430224 152862 430252 163200
rect 430592 152998 430620 163254
rect 430960 163146 430988 163254
rect 431038 163200 431094 164400
rect 431236 163254 431816 163282
rect 431052 163146 431080 163200
rect 430960 163118 431080 163146
rect 430580 152992 430632 152998
rect 430580 152934 430632 152940
rect 430212 152856 430264 152862
rect 430212 152798 430264 152804
rect 430028 152788 430080 152794
rect 430028 152730 430080 152736
rect 430040 152454 430068 152730
rect 431236 152561 431264 163254
rect 431788 163146 431816 163254
rect 431866 163200 431922 164400
rect 431972 163254 432644 163282
rect 431880 163146 431908 163200
rect 431788 163118 431908 163146
rect 431316 153332 431368 153338
rect 431316 153274 431368 153280
rect 431222 152552 431278 152561
rect 431222 152487 431278 152496
rect 430028 152448 430080 152454
rect 430028 152390 430080 152396
rect 430578 152416 430634 152425
rect 430578 152351 430634 152360
rect 429948 150198 430022 150226
rect 429304 150062 429378 150090
rect 429350 149940 429378 150062
rect 429994 149940 430022 150198
rect 430592 150090 430620 152351
rect 431328 152182 431356 153274
rect 431868 153264 431920 153270
rect 431868 153206 431920 153212
rect 431880 153066 431908 153206
rect 431972 153066 432000 163254
rect 432616 163146 432644 163254
rect 432694 163200 432750 164400
rect 433522 163200 433578 164400
rect 434350 163200 434406 164400
rect 434732 163254 435128 163282
rect 432708 163146 432736 163200
rect 432616 163118 432736 163146
rect 432512 159520 432564 159526
rect 432512 159462 432564 159468
rect 432420 153808 432472 153814
rect 432420 153750 432472 153756
rect 431868 153060 431920 153066
rect 431868 153002 431920 153008
rect 431960 153060 432012 153066
rect 431960 153002 432012 153008
rect 431224 152176 431276 152182
rect 431224 152118 431276 152124
rect 431316 152176 431368 152182
rect 431316 152118 431368 152124
rect 431236 150090 431264 152118
rect 432432 152114 432460 153750
rect 432420 152108 432472 152114
rect 432420 152050 432472 152056
rect 431868 151836 431920 151842
rect 431868 151778 431920 151784
rect 431880 150090 431908 151778
rect 432524 150226 432552 159462
rect 432696 153196 432748 153202
rect 432696 153138 432748 153144
rect 432708 152522 432736 153138
rect 432788 153128 432840 153134
rect 432788 153070 432840 153076
rect 432604 152516 432656 152522
rect 432604 152458 432656 152464
rect 432696 152516 432748 152522
rect 432696 152458 432748 152464
rect 432616 151842 432644 152458
rect 432800 152318 432828 153070
rect 433536 152930 433564 163200
rect 434364 153202 434392 163200
rect 433800 153196 433852 153202
rect 433800 153138 433852 153144
rect 434352 153196 434404 153202
rect 434352 153138 434404 153144
rect 433156 152924 433208 152930
rect 433156 152866 433208 152872
rect 433524 152924 433576 152930
rect 433524 152866 433576 152872
rect 432696 152312 432748 152318
rect 432696 152254 432748 152260
rect 432788 152312 432840 152318
rect 432788 152254 432840 152260
rect 432708 152046 432736 152254
rect 432696 152040 432748 152046
rect 432696 151982 432748 151988
rect 432604 151836 432656 151842
rect 432604 151778 432656 151784
rect 432524 150198 432598 150226
rect 430592 150062 430666 150090
rect 431236 150062 431310 150090
rect 431880 150062 431954 150090
rect 430638 149940 430666 150062
rect 431282 149940 431310 150062
rect 431926 149940 431954 150062
rect 432570 149940 432598 150198
rect 433168 150090 433196 152866
rect 433812 150090 433840 153138
rect 434732 152794 434760 163254
rect 435100 163146 435128 163254
rect 435178 163200 435234 164400
rect 436098 163200 436154 164400
rect 436204 163254 436876 163282
rect 435192 163146 435220 163200
rect 435100 163118 435220 163146
rect 435088 159384 435140 159390
rect 435088 159326 435140 159332
rect 434536 152788 434588 152794
rect 434536 152730 434588 152736
rect 434720 152788 434772 152794
rect 434720 152730 434772 152736
rect 434548 151978 434576 152730
rect 434536 151972 434588 151978
rect 434536 151914 434588 151920
rect 435100 150226 435128 159326
rect 436112 153134 436140 163200
rect 436100 153128 436152 153134
rect 436100 153070 436152 153076
rect 436204 152522 436232 163254
rect 436848 163146 436876 163254
rect 436926 163200 436982 164400
rect 437492 163254 437704 163282
rect 436940 163146 436968 163200
rect 436848 163118 436968 163146
rect 437112 152652 437164 152658
rect 437112 152594 437164 152600
rect 436192 152516 436244 152522
rect 436192 152458 436244 152464
rect 435732 152448 435784 152454
rect 435732 152390 435784 152396
rect 436376 152448 436428 152454
rect 436376 152390 436428 152396
rect 435100 150198 435174 150226
rect 434490 150136 434542 150142
rect 433168 150062 433242 150090
rect 433812 150062 433886 150090
rect 434490 150078 434542 150084
rect 433214 149940 433242 150062
rect 433858 149940 433886 150062
rect 434502 149940 434530 150078
rect 435146 149940 435174 150198
rect 435744 150090 435772 152390
rect 436388 150090 436416 152390
rect 437124 151910 437152 152594
rect 437492 152454 437520 163254
rect 437676 163146 437704 163254
rect 437754 163200 437810 164400
rect 437860 163254 438532 163282
rect 437768 163146 437796 163200
rect 437676 163118 437796 163146
rect 437664 159656 437716 159662
rect 437664 159598 437716 159604
rect 437572 153400 437624 153406
rect 437572 153342 437624 153348
rect 437584 153134 437612 153342
rect 437572 153128 437624 153134
rect 437572 153070 437624 153076
rect 437480 152448 437532 152454
rect 437480 152390 437532 152396
rect 437020 151904 437072 151910
rect 437020 151846 437072 151852
rect 437112 151904 437164 151910
rect 437112 151846 437164 151852
rect 437032 150090 437060 151846
rect 437676 150226 437704 159598
rect 437860 153202 437888 163254
rect 438504 163146 438532 163254
rect 438582 163200 438638 164400
rect 438872 163254 439360 163282
rect 438596 163146 438624 163200
rect 438504 163118 438624 163146
rect 437848 153196 437900 153202
rect 437848 153138 437900 153144
rect 438400 153196 438452 153202
rect 438400 153138 438452 153144
rect 438412 152386 438440 153138
rect 438872 152794 438900 163254
rect 439332 163146 439360 163254
rect 439410 163200 439466 164400
rect 440238 163200 440294 164400
rect 440344 163254 441016 163282
rect 439424 163146 439452 163200
rect 439332 163118 439452 163146
rect 440252 153202 440280 163200
rect 440240 153196 440292 153202
rect 440240 153138 440292 153144
rect 438860 152788 438912 152794
rect 438860 152730 438912 152736
rect 440344 152726 440372 163254
rect 440988 163146 441016 163254
rect 441066 163200 441122 164400
rect 441632 163254 441936 163282
rect 441080 163146 441108 163200
rect 440988 163118 441108 163146
rect 440424 159724 440476 159730
rect 440424 159666 440476 159672
rect 440240 152720 440292 152726
rect 440240 152662 440292 152668
rect 440332 152720 440384 152726
rect 440332 152662 440384 152668
rect 438308 152380 438360 152386
rect 438308 152322 438360 152328
rect 438400 152380 438452 152386
rect 438400 152322 438452 152328
rect 437676 150198 437750 150226
rect 435744 150062 435818 150090
rect 436388 150062 436462 150090
rect 437032 150062 437106 150090
rect 435790 149940 435818 150062
rect 436434 149940 436462 150062
rect 437078 149940 437106 150062
rect 437722 149940 437750 150198
rect 438320 150090 438348 152322
rect 438952 152312 439004 152318
rect 438952 152254 439004 152260
rect 438964 150090 438992 152254
rect 440252 151978 440280 152662
rect 439596 151972 439648 151978
rect 439596 151914 439648 151920
rect 440240 151972 440292 151978
rect 440240 151914 440292 151920
rect 439608 150090 439636 151914
rect 440436 150226 440464 159666
rect 440516 153196 440568 153202
rect 440516 153138 440568 153144
rect 440528 152318 440556 153138
rect 441632 152658 441660 163254
rect 441908 163146 441936 163254
rect 441986 163200 442042 164400
rect 442092 163254 442764 163282
rect 442000 163146 442028 163200
rect 441908 163118 442028 163146
rect 441988 153264 442040 153270
rect 441988 153206 442040 153212
rect 442000 153066 442028 153206
rect 441988 153060 442040 153066
rect 441988 153002 442040 153008
rect 441436 152652 441488 152658
rect 441436 152594 441488 152600
rect 441620 152652 441672 152658
rect 441620 152594 441672 152600
rect 440516 152312 440568 152318
rect 440516 152254 440568 152260
rect 441448 151842 441476 152594
rect 442092 152590 442120 163254
rect 442736 163146 442764 163254
rect 442814 163200 442870 164400
rect 443196 163254 443592 163282
rect 442828 163146 442856 163200
rect 442736 163118 442856 163146
rect 442816 159792 442868 159798
rect 442816 159734 442868 159740
rect 442172 153196 442224 153202
rect 442172 153138 442224 153144
rect 442184 152946 442212 153138
rect 442540 153128 442592 153134
rect 442276 153076 442540 153082
rect 442276 153070 442592 153076
rect 442276 153066 442580 153070
rect 442264 153060 442580 153066
rect 442316 153054 442580 153060
rect 442264 153002 442316 153008
rect 442356 152992 442408 152998
rect 442184 152918 442304 152946
rect 442540 152992 442592 152998
rect 442408 152940 442540 152946
rect 442356 152934 442592 152940
rect 442368 152918 442580 152934
rect 441528 152584 441580 152590
rect 441528 152526 441580 152532
rect 442080 152584 442132 152590
rect 442080 152526 442132 152532
rect 440884 151836 440936 151842
rect 440884 151778 440936 151784
rect 441436 151836 441488 151842
rect 441436 151778 441488 151784
rect 440298 150198 440464 150226
rect 440896 150226 440924 151778
rect 440896 150198 440970 150226
rect 438320 150062 438394 150090
rect 438964 150062 439038 150090
rect 439608 150062 439682 150090
rect 438366 149940 438394 150062
rect 439010 149940 439038 150062
rect 439654 149940 439682 150062
rect 440298 149940 440326 150198
rect 440942 149940 440970 150198
rect 441540 150090 441568 152526
rect 442276 151910 442304 152918
rect 442172 151904 442224 151910
rect 442172 151846 442224 151852
rect 442264 151904 442316 151910
rect 442264 151846 442316 151852
rect 442184 150226 442212 151846
rect 442828 150226 442856 159734
rect 443196 152930 443224 163254
rect 443564 163146 443592 163254
rect 443642 163200 443698 164400
rect 444470 163200 444526 164400
rect 445298 163200 445354 164400
rect 446126 163200 446182 164400
rect 446324 163254 446904 163282
rect 443656 163146 443684 163200
rect 443564 163118 443684 163146
rect 444484 153134 444512 163200
rect 443552 153128 443604 153134
rect 443552 153070 443604 153076
rect 444472 153128 444524 153134
rect 444472 153070 444524 153076
rect 443184 152924 443236 152930
rect 443184 152866 443236 152872
rect 443564 152046 443592 153070
rect 444654 152688 444710 152697
rect 444654 152623 444710 152632
rect 444748 152652 444800 152658
rect 444668 152590 444696 152623
rect 444748 152594 444800 152600
rect 444656 152584 444708 152590
rect 444656 152526 444708 152532
rect 444760 152538 444788 152594
rect 444564 152516 444616 152522
rect 444760 152510 445156 152538
rect 444564 152458 444616 152464
rect 444472 152448 444524 152454
rect 444472 152390 444524 152396
rect 444576 152402 444604 152458
rect 444104 152176 444156 152182
rect 444104 152118 444156 152124
rect 443460 152040 443512 152046
rect 443460 151982 443512 151988
rect 443552 152040 443604 152046
rect 443552 151982 443604 151988
rect 442184 150198 442258 150226
rect 442828 150198 442902 150226
rect 441540 150062 441614 150090
rect 441586 149940 441614 150062
rect 442230 149940 442258 150198
rect 442874 149940 442902 150198
rect 443472 150090 443500 151982
rect 444116 150090 444144 152118
rect 444484 150210 444512 152390
rect 444576 152374 444880 152402
rect 445128 152386 445156 152510
rect 444748 152108 444800 152114
rect 444748 152050 444800 152056
rect 444472 150204 444524 150210
rect 444472 150146 444524 150152
rect 444760 150090 444788 152050
rect 444852 151910 444880 152374
rect 445116 152380 445168 152386
rect 445116 152322 445168 152328
rect 445312 152046 445340 163200
rect 445392 159452 445444 159458
rect 445392 159394 445444 159400
rect 445300 152040 445352 152046
rect 445300 151982 445352 151988
rect 444840 151904 444892 151910
rect 444840 151846 444892 151852
rect 445404 150226 445432 159394
rect 446140 158982 446168 163200
rect 446128 158976 446180 158982
rect 446128 158918 446180 158924
rect 445484 152720 445536 152726
rect 445484 152662 445536 152668
rect 445574 152688 445630 152697
rect 445496 152522 445524 152662
rect 445574 152623 445630 152632
rect 445588 152590 445616 152623
rect 445576 152584 445628 152590
rect 445576 152526 445628 152532
rect 445484 152516 445536 152522
rect 445484 152458 445536 152464
rect 446324 152114 446352 163254
rect 446876 163146 446904 163254
rect 446954 163200 447010 164400
rect 447874 163200 447930 164400
rect 448702 163200 448758 164400
rect 449530 163200 449586 164400
rect 450358 163200 450414 164400
rect 451186 163200 451242 164400
rect 452014 163200 452070 164400
rect 452842 163200 452898 164400
rect 453762 163200 453818 164400
rect 454590 163200 454646 164400
rect 455418 163200 455474 164400
rect 456246 163200 456302 164400
rect 457074 163200 457130 164400
rect 457902 163200 457958 164400
rect 458730 163200 458786 164400
rect 459650 163200 459706 164400
rect 460478 163200 460534 164400
rect 461306 163200 461362 164400
rect 462134 163200 462190 164400
rect 462962 163200 463018 164400
rect 463790 163200 463846 164400
rect 464618 163200 464674 164400
rect 465538 163200 465594 164400
rect 466366 163200 466422 164400
rect 467194 163200 467250 164400
rect 468022 163200 468078 164400
rect 468850 163200 468906 164400
rect 469678 163200 469734 164400
rect 470506 163200 470562 164400
rect 471426 163200 471482 164400
rect 472254 163200 472310 164400
rect 473082 163200 473138 164400
rect 473910 163200 473966 164400
rect 474738 163200 474794 164400
rect 475566 163200 475622 164400
rect 476394 163200 476450 164400
rect 477314 163200 477370 164400
rect 478142 163200 478198 164400
rect 478970 163200 479026 164400
rect 479798 163200 479854 164400
rect 480626 163200 480682 164400
rect 481454 163200 481510 164400
rect 482282 163200 482338 164400
rect 483202 163200 483258 164400
rect 484030 163200 484086 164400
rect 484504 163254 484808 163282
rect 446968 163146 446996 163200
rect 446876 163118 446996 163146
rect 447888 159390 447916 163200
rect 448716 159662 448744 163200
rect 448704 159656 448756 159662
rect 448704 159598 448756 159604
rect 449544 159526 449572 163200
rect 450372 159594 450400 163200
rect 450360 159588 450412 159594
rect 450360 159530 450412 159536
rect 449532 159520 449584 159526
rect 449532 159462 449584 159468
rect 451200 159458 451228 163200
rect 451188 159452 451240 159458
rect 451188 159394 451240 159400
rect 447876 159384 447928 159390
rect 447876 159326 447928 159332
rect 452028 158778 452056 163200
rect 452856 159118 452884 163200
rect 453776 159254 453804 163200
rect 453764 159248 453816 159254
rect 453764 159190 453816 159196
rect 452844 159112 452896 159118
rect 452844 159054 452896 159060
rect 454604 158982 454632 163200
rect 455432 159050 455460 163200
rect 455880 159656 455932 159662
rect 455880 159598 455932 159604
rect 455512 159520 455564 159526
rect 455512 159462 455564 159468
rect 455420 159044 455472 159050
rect 455420 158986 455472 158992
rect 453856 158976 453908 158982
rect 453856 158918 453908 158924
rect 454592 158976 454644 158982
rect 454592 158918 454644 158924
rect 452016 158772 452068 158778
rect 452016 158714 452068 158720
rect 453868 153202 453896 158918
rect 449256 153196 449308 153202
rect 449256 153138 449308 153144
rect 453856 153196 453908 153202
rect 453856 153138 453908 153144
rect 447968 152992 448020 152998
rect 447968 152934 448020 152940
rect 447324 152856 447376 152862
rect 447324 152798 447376 152804
rect 446680 152244 446732 152250
rect 446680 152186 446732 152192
rect 446312 152108 446364 152114
rect 446312 152050 446364 152056
rect 446036 151700 446088 151706
rect 446036 151642 446088 151648
rect 445404 150198 445478 150226
rect 443472 150062 443546 150090
rect 444116 150062 444190 150090
rect 444760 150062 444834 150090
rect 443518 149940 443546 150062
rect 444162 149940 444190 150062
rect 444806 149940 444834 150062
rect 445450 149940 445478 150198
rect 446048 150090 446076 151642
rect 446692 150090 446720 152186
rect 447336 150226 447364 152798
rect 447980 150226 448008 152934
rect 448610 152552 448666 152561
rect 448610 152487 448666 152496
rect 448624 150226 448652 152487
rect 449268 150226 449296 153138
rect 449900 153060 449952 153066
rect 449900 153002 449952 153008
rect 449912 150226 449940 153002
rect 451188 152924 451240 152930
rect 451188 152866 451240 152872
rect 450544 152176 450596 152182
rect 450544 152118 450596 152124
rect 450556 150226 450584 152118
rect 451200 151978 451228 152866
rect 454408 152788 454460 152794
rect 454408 152730 454460 152736
rect 453764 152448 453816 152454
rect 453764 152390 453816 152396
rect 451096 151972 451148 151978
rect 451096 151914 451148 151920
rect 451188 151972 451240 151978
rect 451188 151914 451240 151920
rect 451108 151814 451136 151914
rect 452476 151904 452528 151910
rect 452476 151846 452528 151852
rect 451832 151836 451884 151842
rect 451108 151786 451228 151814
rect 451200 150226 451228 151786
rect 451832 151778 451884 151784
rect 451844 150226 451872 151778
rect 452488 150226 452516 151846
rect 453776 150226 453804 152390
rect 454420 150226 454448 152730
rect 455524 152318 455552 159462
rect 455696 152516 455748 152522
rect 455696 152458 455748 152464
rect 455052 152312 455104 152318
rect 455052 152254 455104 152260
rect 455512 152312 455564 152318
rect 455512 152254 455564 152260
rect 455064 150226 455092 152254
rect 455708 150226 455736 152458
rect 455892 152182 455920 159598
rect 456260 158914 456288 163200
rect 457088 159526 457116 163200
rect 457168 159588 457220 159594
rect 457168 159530 457220 159536
rect 457076 159520 457128 159526
rect 457076 159462 457128 159468
rect 456800 159452 456852 159458
rect 456800 159394 456852 159400
rect 456248 158908 456300 158914
rect 456248 158850 456300 158856
rect 456340 152380 456392 152386
rect 456340 152322 456392 152328
rect 455880 152176 455932 152182
rect 455880 152118 455932 152124
rect 456352 150226 456380 152322
rect 456812 152250 456840 159394
rect 456892 159384 456944 159390
rect 456892 159326 456944 159332
rect 456904 153066 456932 159326
rect 456892 153060 456944 153066
rect 456892 153002 456944 153008
rect 456984 152584 457036 152590
rect 456984 152526 457036 152532
rect 456800 152244 456852 152250
rect 456800 152186 456852 152192
rect 456996 150226 457024 152526
rect 457180 151842 457208 159530
rect 457916 159186 457944 163200
rect 458744 159594 458772 163200
rect 458732 159588 458784 159594
rect 458732 159530 458784 159536
rect 459664 159458 459692 163200
rect 459652 159452 459704 159458
rect 459652 159394 459704 159400
rect 460492 159322 460520 163200
rect 460480 159316 460532 159322
rect 460480 159258 460532 159264
rect 459560 159248 459612 159254
rect 459560 159190 459612 159196
rect 457904 159180 457956 159186
rect 457904 159122 457956 159128
rect 458180 158772 458232 158778
rect 458180 158714 458232 158720
rect 458192 152590 458220 158714
rect 459468 153196 459520 153202
rect 459468 153138 459520 153144
rect 458272 153128 458324 153134
rect 458272 153070 458324 153076
rect 458180 152584 458232 152590
rect 458180 152526 458232 152532
rect 457628 151972 457680 151978
rect 457628 151914 457680 151920
rect 457168 151836 457220 151842
rect 457168 151778 457220 151784
rect 457640 150226 457668 151914
rect 458284 150226 458312 153070
rect 458824 152040 458876 152046
rect 458824 151982 458876 151988
rect 447336 150198 447410 150226
rect 447980 150198 448054 150226
rect 448624 150198 448698 150226
rect 449268 150198 449342 150226
rect 449912 150198 449986 150226
rect 450556 150198 450630 150226
rect 451200 150198 451274 150226
rect 451844 150198 451918 150226
rect 452488 150198 452562 150226
rect 446048 150062 446122 150090
rect 446692 150062 446766 150090
rect 446094 149940 446122 150062
rect 446738 149940 446766 150062
rect 447382 149940 447410 150198
rect 448026 149940 448054 150198
rect 448670 149940 448698 150198
rect 449314 149940 449342 150198
rect 449958 149940 449986 150198
rect 450602 149940 450630 150198
rect 451246 149940 451274 150198
rect 451890 149940 451918 150198
rect 452534 149940 452562 150198
rect 453166 150204 453218 150210
rect 453776 150198 453850 150226
rect 454420 150198 454494 150226
rect 455064 150198 455138 150226
rect 455708 150198 455782 150226
rect 456352 150198 456426 150226
rect 456996 150198 457070 150226
rect 457640 150198 457714 150226
rect 453166 150146 453218 150152
rect 453178 149940 453206 150146
rect 453822 149940 453850 150198
rect 454466 149940 454494 150198
rect 455110 149940 455138 150198
rect 455754 149940 455782 150198
rect 456398 149940 456426 150198
rect 457042 149940 457070 150198
rect 457686 149940 457714 150198
rect 458238 150198 458312 150226
rect 458836 150226 458864 151982
rect 459480 150226 459508 153138
rect 459572 152658 459600 159190
rect 461320 159118 461348 163200
rect 459652 159112 459704 159118
rect 459652 159054 459704 159060
rect 461308 159112 461360 159118
rect 461308 159054 461360 159060
rect 459664 152930 459692 159054
rect 461860 158976 461912 158982
rect 461860 158918 461912 158924
rect 461872 153202 461900 158918
rect 462148 158778 462176 163200
rect 462976 159254 463004 163200
rect 462964 159248 463016 159254
rect 462964 159190 463016 159196
rect 463516 159044 463568 159050
rect 463516 158986 463568 158992
rect 462964 158908 463016 158914
rect 462964 158850 463016 158856
rect 462136 158772 462188 158778
rect 462136 158714 462188 158720
rect 461860 153196 461912 153202
rect 461860 153138 461912 153144
rect 462976 153134 463004 158850
rect 462964 153128 463016 153134
rect 462964 153070 463016 153076
rect 463528 153066 463556 158986
rect 463804 158846 463832 163200
rect 464344 159520 464396 159526
rect 464344 159462 464396 159468
rect 463884 159180 463936 159186
rect 463884 159122 463936 159128
rect 463792 158840 463844 158846
rect 463792 158782 463844 158788
rect 460756 153060 460808 153066
rect 460756 153002 460808 153008
rect 463516 153060 463568 153066
rect 463516 153002 463568 153008
rect 459652 152924 459704 152930
rect 459652 152866 459704 152872
rect 459560 152652 459612 152658
rect 459560 152594 459612 152600
rect 460112 152108 460164 152114
rect 460112 152050 460164 152056
rect 460124 150226 460152 152050
rect 460768 150226 460796 153002
rect 463896 152998 463924 159122
rect 463884 152992 463936 152998
rect 463884 152934 463936 152940
rect 463976 152584 464028 152590
rect 463976 152526 464028 152532
rect 462044 152312 462096 152318
rect 462044 152254 462096 152260
rect 461400 152176 461452 152182
rect 461400 152118 461452 152124
rect 461412 150226 461440 152118
rect 462056 150226 462084 152254
rect 463332 152244 463384 152250
rect 463332 152186 463384 152192
rect 462688 151836 462740 151842
rect 462688 151778 462740 151784
rect 462700 150226 462728 151778
rect 463344 150226 463372 152186
rect 463988 150226 464016 152526
rect 464356 151842 464384 159462
rect 464632 158982 464660 163200
rect 465080 159588 465132 159594
rect 465080 159530 465132 159536
rect 464620 158976 464672 158982
rect 464620 158918 464672 158924
rect 465092 152930 465120 159530
rect 465552 159050 465580 163200
rect 465540 159044 465592 159050
rect 465540 158986 465592 158992
rect 466380 158914 466408 163200
rect 467208 159866 467236 163200
rect 467196 159860 467248 159866
rect 467196 159802 467248 159808
rect 468036 159594 468064 163200
rect 468024 159588 468076 159594
rect 468024 159530 468076 159536
rect 468864 159458 468892 163200
rect 466460 159452 466512 159458
rect 466460 159394 466512 159400
rect 468852 159452 468904 159458
rect 468852 159394 468904 159400
rect 466368 158908 466420 158914
rect 466368 158850 466420 158856
rect 466472 153202 466500 159394
rect 469692 159390 469720 163200
rect 470520 159934 470548 163200
rect 471440 159934 471468 163200
rect 470508 159928 470560 159934
rect 470508 159870 470560 159876
rect 471428 159928 471480 159934
rect 471428 159870 471480 159876
rect 472268 159798 472296 163200
rect 472256 159792 472308 159798
rect 472256 159734 472308 159740
rect 469680 159384 469732 159390
rect 469680 159326 469732 159332
rect 466644 159316 466696 159322
rect 466644 159258 466696 159264
rect 465908 153196 465960 153202
rect 465908 153138 465960 153144
rect 466460 153196 466512 153202
rect 466460 153138 466512 153144
rect 464620 152924 464672 152930
rect 464620 152866 464672 152872
rect 465080 152924 465132 152930
rect 465080 152866 465132 152872
rect 464344 151836 464396 151842
rect 464344 151778 464396 151784
rect 464632 150226 464660 152866
rect 465264 152652 465316 152658
rect 465264 152594 465316 152600
rect 465276 150226 465304 152594
rect 465920 150226 465948 153138
rect 466656 153066 466684 159258
rect 469220 159248 469272 159254
rect 469220 159190 469272 159196
rect 467840 159112 467892 159118
rect 467840 159054 467892 159060
rect 467288 153128 467340 153134
rect 467288 153070 467340 153076
rect 466552 153060 466604 153066
rect 466552 153002 466604 153008
rect 466644 153060 466696 153066
rect 466644 153002 466696 153008
rect 466564 150226 466592 153002
rect 467300 150226 467328 153070
rect 467852 151910 467880 159054
rect 467932 158772 467984 158778
rect 467932 158714 467984 158720
rect 467840 151904 467892 151910
rect 467840 151846 467892 151852
rect 467944 151842 467972 158714
rect 468392 152992 468444 152998
rect 468392 152934 468444 152940
rect 467748 151836 467800 151842
rect 467932 151836 467984 151842
rect 467800 151786 467880 151814
rect 467748 151778 467800 151784
rect 458836 150198 458910 150226
rect 459480 150198 459554 150226
rect 460124 150198 460198 150226
rect 460768 150198 460842 150226
rect 461412 150198 461486 150226
rect 462056 150198 462130 150226
rect 462700 150198 462774 150226
rect 463344 150198 463418 150226
rect 463988 150198 464062 150226
rect 464632 150198 464706 150226
rect 465276 150198 465350 150226
rect 465920 150198 465994 150226
rect 466564 150198 466638 150226
rect 458238 149940 458266 150198
rect 458882 149940 458910 150198
rect 459526 149940 459554 150198
rect 460170 149940 460198 150198
rect 460814 149940 460842 150198
rect 461458 149940 461486 150198
rect 462102 149940 462130 150198
rect 462746 149940 462774 150198
rect 463390 149940 463418 150198
rect 464034 149940 464062 150198
rect 464678 149940 464706 150198
rect 465322 149940 465350 150198
rect 465966 149940 465994 150198
rect 466610 149940 466638 150198
rect 467254 150198 467328 150226
rect 467852 150226 467880 151786
rect 468404 151814 468432 152934
rect 469128 152924 469180 152930
rect 469128 152866 469180 152872
rect 468404 151786 468524 151814
rect 467932 151778 467984 151784
rect 468496 150226 468524 151786
rect 469140 150226 469168 152866
rect 469232 151978 469260 159190
rect 472440 159044 472492 159050
rect 472440 158986 472492 158992
rect 471244 158976 471296 158982
rect 471244 158918 471296 158924
rect 469772 153196 469824 153202
rect 469772 153138 469824 153144
rect 469220 151972 469272 151978
rect 469220 151914 469272 151920
rect 469784 150226 469812 153138
rect 471256 153134 471284 158918
rect 472348 158908 472400 158914
rect 472348 158850 472400 158856
rect 471428 158840 471480 158846
rect 471428 158782 471480 158788
rect 471440 153202 471468 158782
rect 471428 153196 471480 153202
rect 471428 153138 471480 153144
rect 471244 153128 471296 153134
rect 471244 153070 471296 153076
rect 472360 153066 472388 158850
rect 470416 153060 470468 153066
rect 470416 153002 470468 153008
rect 472348 153060 472400 153066
rect 472348 153002 472400 153008
rect 470428 150226 470456 153002
rect 472452 152998 472480 158986
rect 473096 158778 473124 163200
rect 473360 159860 473412 159866
rect 473360 159802 473412 159808
rect 473084 158772 473136 158778
rect 473084 158714 473136 158720
rect 473372 153202 473400 159802
rect 473924 159050 473952 163200
rect 473912 159044 473964 159050
rect 473912 158986 473964 158992
rect 474752 158914 474780 163200
rect 474832 159452 474884 159458
rect 474832 159394 474884 159400
rect 474740 158908 474792 158914
rect 474740 158850 474792 158856
rect 472992 153196 473044 153202
rect 472992 153138 473044 153144
rect 473360 153196 473412 153202
rect 473360 153138 473412 153144
rect 472440 152992 472492 152998
rect 472440 152934 472492 152940
rect 472348 151972 472400 151978
rect 472348 151914 472400 151920
rect 471060 151904 471112 151910
rect 471060 151846 471112 151852
rect 471072 150226 471100 151846
rect 471704 151836 471756 151842
rect 471704 151778 471756 151784
rect 471716 150226 471744 151778
rect 472360 150226 472388 151914
rect 473004 150226 473032 153138
rect 474844 153134 474872 159394
rect 475580 158982 475608 163200
rect 476120 159996 476172 160002
rect 476120 159938 476172 159944
rect 476028 159588 476080 159594
rect 476028 159530 476080 159536
rect 475568 158976 475620 158982
rect 475568 158918 475620 158924
rect 475568 153196 475620 153202
rect 475568 153138 475620 153144
rect 473636 153128 473688 153134
rect 473636 153070 473688 153076
rect 474832 153128 474884 153134
rect 474832 153070 474884 153076
rect 473648 150226 473676 153070
rect 474924 153060 474976 153066
rect 474924 153002 474976 153008
rect 474280 152992 474332 152998
rect 474280 152934 474332 152940
rect 474292 150226 474320 152934
rect 474936 150226 474964 153002
rect 475580 150226 475608 153138
rect 476040 151814 476068 159530
rect 476132 153202 476160 159938
rect 476408 158846 476436 163200
rect 477328 159458 477356 163200
rect 477684 159928 477736 159934
rect 477684 159870 477736 159876
rect 477316 159452 477368 159458
rect 477316 159394 477368 159400
rect 477408 159384 477460 159390
rect 477408 159326 477460 159332
rect 476396 158840 476448 158846
rect 476396 158782 476448 158788
rect 476120 153196 476172 153202
rect 476120 153138 476172 153144
rect 476948 153128 477000 153134
rect 476948 153070 477000 153076
rect 476040 151786 476252 151814
rect 476224 150226 476252 151786
rect 476960 150226 476988 153070
rect 477420 151814 477448 159326
rect 477420 151786 477540 151814
rect 467852 150198 467926 150226
rect 468496 150198 468570 150226
rect 469140 150198 469214 150226
rect 469784 150198 469858 150226
rect 470428 150198 470502 150226
rect 471072 150198 471146 150226
rect 471716 150198 471790 150226
rect 472360 150198 472434 150226
rect 473004 150198 473078 150226
rect 473648 150198 473722 150226
rect 474292 150198 474366 150226
rect 474936 150198 475010 150226
rect 475580 150198 475654 150226
rect 476224 150198 476298 150226
rect 467254 149940 467282 150198
rect 467898 149940 467926 150198
rect 468542 149940 468570 150198
rect 469186 149940 469214 150198
rect 469830 149940 469858 150198
rect 470474 149940 470502 150198
rect 471118 149940 471146 150198
rect 471762 149940 471790 150198
rect 472406 149940 472434 150198
rect 473050 149940 473078 150198
rect 473694 149940 473722 150198
rect 474338 149940 474366 150198
rect 474982 149940 475010 150198
rect 475626 149940 475654 150198
rect 476270 149940 476298 150198
rect 476914 150198 476988 150226
rect 477512 150226 477540 151786
rect 477512 150198 477586 150226
rect 477696 150210 477724 159870
rect 478156 159390 478184 163200
rect 478984 159594 479012 163200
rect 479812 159798 479840 163200
rect 480640 159934 480668 163200
rect 480628 159928 480680 159934
rect 480628 159870 480680 159876
rect 479432 159792 479484 159798
rect 479432 159734 479484 159740
rect 479800 159792 479852 159798
rect 479800 159734 479852 159740
rect 478972 159588 479024 159594
rect 478972 159530 479024 159536
rect 478144 159384 478196 159390
rect 478144 159326 478196 159332
rect 478972 158772 479024 158778
rect 478972 158714 479024 158720
rect 478144 153196 478196 153202
rect 478144 153138 478196 153144
rect 478156 150226 478184 153138
rect 476914 149940 476942 150198
rect 477558 149940 477586 150198
rect 477684 150204 477736 150210
rect 478156 150198 478230 150226
rect 478984 150210 479012 158714
rect 479444 150226 479472 159734
rect 480260 159044 480312 159050
rect 480260 158986 480312 158992
rect 480272 151814 480300 158986
rect 481468 158914 481496 163200
rect 482008 158976 482060 158982
rect 482008 158918 482060 158924
rect 481364 158908 481416 158914
rect 481364 158850 481416 158856
rect 481456 158908 481508 158914
rect 481456 158850 481508 158856
rect 480272 151786 480760 151814
rect 480732 150226 480760 151786
rect 481376 150226 481404 158850
rect 481640 158840 481692 158846
rect 481640 158782 481692 158788
rect 477684 150146 477736 150152
rect 478202 149940 478230 150198
rect 478834 150204 478886 150210
rect 478834 150146 478886 150152
rect 478972 150204 479024 150210
rect 479444 150198 479518 150226
rect 478972 150146 479024 150152
rect 478846 149940 478874 150146
rect 479490 149940 479518 150198
rect 480122 150204 480174 150210
rect 480732 150198 480806 150226
rect 481376 150198 481450 150226
rect 481652 150210 481680 158782
rect 482020 150226 482048 158918
rect 482296 158778 482324 163200
rect 483216 161474 483244 163200
rect 483124 161446 483244 161474
rect 482284 158772 482336 158778
rect 482284 158714 482336 158720
rect 483124 152998 483152 161446
rect 483296 159452 483348 159458
rect 483296 159394 483348 159400
rect 483204 159384 483256 159390
rect 483204 159326 483256 159332
rect 483112 152992 483164 152998
rect 483112 152934 483164 152940
rect 480122 150146 480174 150152
rect 480134 149940 480162 150146
rect 480778 149940 480806 150198
rect 481422 149940 481450 150198
rect 481640 150204 481692 150210
rect 482020 150198 482094 150226
rect 483216 150210 483244 159326
rect 483308 150226 483336 159394
rect 484044 153134 484072 163200
rect 484032 153128 484084 153134
rect 484032 153070 484084 153076
rect 484504 153066 484532 163254
rect 484780 163146 484808 163254
rect 484858 163200 484914 164400
rect 485686 163200 485742 164400
rect 485792 163254 486464 163282
rect 484872 163146 484900 163200
rect 484780 163118 484900 163146
rect 485228 159792 485280 159798
rect 485228 159734 485280 159740
rect 484584 159588 484636 159594
rect 484584 159530 484636 159536
rect 484492 153060 484544 153066
rect 484492 153002 484544 153008
rect 484596 150226 484624 159530
rect 485240 150226 485268 159734
rect 485700 153202 485728 163200
rect 485688 153196 485740 153202
rect 485688 153138 485740 153144
rect 485792 152046 485820 163254
rect 486436 163146 486464 163254
rect 486514 163200 486570 164400
rect 487342 163200 487398 164400
rect 488170 163200 488226 164400
rect 488552 163254 489040 163282
rect 486528 163146 486556 163200
rect 486436 163118 486556 163146
rect 485964 159928 486016 159934
rect 485964 159870 486016 159876
rect 485780 152040 485832 152046
rect 485780 151982 485832 151988
rect 485976 150226 486004 159870
rect 486516 158908 486568 158914
rect 486516 158850 486568 158856
rect 481640 150146 481692 150152
rect 482066 149940 482094 150198
rect 482698 150204 482750 150210
rect 482698 150146 482750 150152
rect 483204 150204 483256 150210
rect 483308 150198 483382 150226
rect 483204 150146 483256 150152
rect 482710 149940 482738 150146
rect 483354 149940 483382 150198
rect 483986 150204 484038 150210
rect 484596 150198 484670 150226
rect 485240 150198 485314 150226
rect 483986 150146 484038 150152
rect 483998 149940 484026 150146
rect 484642 149940 484670 150198
rect 485286 149940 485314 150198
rect 485930 150198 486004 150226
rect 486528 150226 486556 158850
rect 487252 158772 487304 158778
rect 487252 158714 487304 158720
rect 487264 150226 487292 158714
rect 487356 151978 487384 163200
rect 487804 152992 487856 152998
rect 487804 152934 487856 152940
rect 487344 151972 487396 151978
rect 487344 151914 487396 151920
rect 486528 150198 486602 150226
rect 485930 149940 485958 150198
rect 486574 149940 486602 150198
rect 487218 150198 487292 150226
rect 487816 150226 487844 152934
rect 488184 151842 488212 163200
rect 488448 153128 488500 153134
rect 488448 153070 488500 153076
rect 488172 151836 488224 151842
rect 488172 151778 488224 151784
rect 488460 150226 488488 153070
rect 488552 151910 488580 163254
rect 489012 163146 489040 163254
rect 489090 163200 489146 164400
rect 489918 163200 489974 164400
rect 490746 163200 490802 164400
rect 491312 163254 491524 163282
rect 489104 163146 489132 163200
rect 489012 163118 489132 163146
rect 489644 153196 489696 153202
rect 489644 153138 489696 153144
rect 489000 153060 489052 153066
rect 489000 153002 489052 153008
rect 488540 151904 488592 151910
rect 488540 151846 488592 151852
rect 489012 150226 489040 153002
rect 489656 150226 489684 153138
rect 489932 153134 489960 163200
rect 490760 153202 490788 163200
rect 490748 153196 490800 153202
rect 490748 153138 490800 153144
rect 489920 153128 489972 153134
rect 489920 153070 489972 153076
rect 491312 152930 491340 163254
rect 491496 163146 491524 163254
rect 491574 163200 491630 164400
rect 491680 163254 492352 163282
rect 491588 163146 491616 163200
rect 491496 163118 491616 163146
rect 491680 152998 491708 163254
rect 492324 163146 492352 163254
rect 492402 163200 492458 164400
rect 492692 163254 493180 163282
rect 492416 163146 492444 163200
rect 492324 163118 492444 163146
rect 492692 153066 492720 163254
rect 493152 163146 493180 163254
rect 493230 163200 493286 164400
rect 494058 163200 494114 164400
rect 494164 163254 494928 163282
rect 493244 163146 493272 163200
rect 493152 163118 493272 163146
rect 494072 153202 494100 163200
rect 493508 153196 493560 153202
rect 493508 153138 493560 153144
rect 494060 153196 494112 153202
rect 494060 153138 494112 153144
rect 492864 153128 492916 153134
rect 492864 153070 492916 153076
rect 492680 153060 492732 153066
rect 492680 153002 492732 153008
rect 491668 152992 491720 152998
rect 491668 152934 491720 152940
rect 491300 152924 491352 152930
rect 491300 152866 491352 152872
rect 490288 152040 490340 152046
rect 490288 151982 490340 151988
rect 490300 150226 490328 151982
rect 490932 151972 490984 151978
rect 490932 151914 490984 151920
rect 490944 150226 490972 151914
rect 492220 151904 492272 151910
rect 492220 151846 492272 151852
rect 491576 151836 491628 151842
rect 491576 151778 491628 151784
rect 491588 150226 491616 151778
rect 492232 150226 492260 151846
rect 492876 150226 492904 153070
rect 493520 150226 493548 153138
rect 494164 153134 494192 163254
rect 494900 163146 494928 163254
rect 494978 163200 495034 164400
rect 495544 163254 495756 163282
rect 494992 163146 495020 163200
rect 494900 163118 495020 163146
rect 494152 153128 494204 153134
rect 494152 153070 494204 153076
rect 495544 153066 495572 163254
rect 495728 163146 495756 163254
rect 495806 163200 495862 164400
rect 496634 163200 496690 164400
rect 496832 163254 497412 163282
rect 495820 163146 495848 163200
rect 495728 163118 495848 163146
rect 496648 153202 496676 163200
rect 496084 153196 496136 153202
rect 496084 153138 496136 153144
rect 496636 153196 496688 153202
rect 496636 153138 496688 153144
rect 495440 153060 495492 153066
rect 495440 153002 495492 153008
rect 495532 153060 495584 153066
rect 495532 153002 495584 153008
rect 494796 152992 494848 152998
rect 494796 152934 494848 152940
rect 494152 152924 494204 152930
rect 494152 152866 494204 152872
rect 494164 150226 494192 152866
rect 494808 150226 494836 152934
rect 495452 150226 495480 153002
rect 496096 150226 496124 153138
rect 496832 153134 496860 163254
rect 497384 163146 497412 163254
rect 497462 163200 497518 164400
rect 498290 163200 498346 164400
rect 499118 163200 499174 164400
rect 499946 163200 500002 164400
rect 500052 163254 500632 163282
rect 497476 163146 497504 163200
rect 497384 163118 497504 163146
rect 498304 156670 498332 163200
rect 498292 156664 498344 156670
rect 498292 156606 498344 156612
rect 498016 153196 498068 153202
rect 498016 153138 498068 153144
rect 496728 153128 496780 153134
rect 496728 153070 496780 153076
rect 496820 153128 496872 153134
rect 496820 153070 496872 153076
rect 496740 150226 496768 153070
rect 497372 153060 497424 153066
rect 497372 153002 497424 153008
rect 497384 150226 497412 153002
rect 498028 150226 498056 153138
rect 498660 153128 498712 153134
rect 498660 153070 498712 153076
rect 498672 150226 498700 153070
rect 499132 151842 499160 163200
rect 499960 163146 499988 163200
rect 500052 163146 500080 163254
rect 499960 163118 500080 163146
rect 499304 156664 499356 156670
rect 499304 156606 499356 156612
rect 499120 151836 499172 151842
rect 499120 151778 499172 151784
rect 499316 150226 499344 156606
rect 499948 151836 500000 151842
rect 499948 151778 500000 151784
rect 499960 150226 499988 151778
rect 500604 150226 500632 163254
rect 500866 163200 500922 164400
rect 501694 163200 501750 164400
rect 502522 163200 502578 164400
rect 503350 163200 503406 164400
rect 503824 163254 504128 163282
rect 500880 151814 500908 163200
rect 501708 161474 501736 163200
rect 501708 161446 501920 161474
rect 500880 151786 501276 151814
rect 501248 150226 501276 151786
rect 501892 150226 501920 161446
rect 502536 150226 502564 163200
rect 503364 151814 503392 163200
rect 503272 151786 503392 151814
rect 503272 150226 503300 151786
rect 487816 150198 487890 150226
rect 488460 150198 488534 150226
rect 489012 150198 489086 150226
rect 489656 150198 489730 150226
rect 490300 150198 490374 150226
rect 490944 150198 491018 150226
rect 491588 150198 491662 150226
rect 492232 150198 492306 150226
rect 492876 150198 492950 150226
rect 493520 150198 493594 150226
rect 494164 150198 494238 150226
rect 494808 150198 494882 150226
rect 495452 150198 495526 150226
rect 496096 150198 496170 150226
rect 496740 150198 496814 150226
rect 497384 150198 497458 150226
rect 498028 150198 498102 150226
rect 498672 150198 498746 150226
rect 499316 150198 499390 150226
rect 499960 150198 500034 150226
rect 500604 150198 500678 150226
rect 501248 150198 501322 150226
rect 501892 150198 501966 150226
rect 502536 150198 502610 150226
rect 487218 149940 487246 150198
rect 487862 149940 487890 150198
rect 488506 149940 488534 150198
rect 489058 149940 489086 150198
rect 489702 149940 489730 150198
rect 490346 149940 490374 150198
rect 490990 149940 491018 150198
rect 491634 149940 491662 150198
rect 492278 149940 492306 150198
rect 492922 149940 492950 150198
rect 493566 149940 493594 150198
rect 494210 149940 494238 150198
rect 494854 149940 494882 150198
rect 495498 149940 495526 150198
rect 496142 149940 496170 150198
rect 496786 149940 496814 150198
rect 497430 149940 497458 150198
rect 498074 149940 498102 150198
rect 498718 149940 498746 150198
rect 499362 149940 499390 150198
rect 500006 149940 500034 150198
rect 500650 149940 500678 150198
rect 501294 149940 501322 150198
rect 501938 149940 501966 150198
rect 502582 149940 502610 150198
rect 503226 150198 503300 150226
rect 503824 150226 503852 163254
rect 504100 163146 504128 163254
rect 504178 163200 504234 164400
rect 504468 163254 504956 163282
rect 504192 163146 504220 163200
rect 504100 163118 504220 163146
rect 504468 150226 504496 163254
rect 504928 163146 504956 163254
rect 505006 163200 505062 164400
rect 505112 163254 505784 163282
rect 505020 163146 505048 163200
rect 504928 163118 505048 163146
rect 505112 150226 505140 163254
rect 505756 163146 505784 163254
rect 505834 163200 505890 164400
rect 506754 163200 506810 164400
rect 507582 163200 507638 164400
rect 508410 163200 508466 164400
rect 509238 163200 509294 164400
rect 509344 163254 509556 163282
rect 505848 163146 505876 163200
rect 505756 163118 505876 163146
rect 505284 158840 505336 158846
rect 505284 158782 505336 158788
rect 503824 150198 503898 150226
rect 504468 150198 504542 150226
rect 505112 150198 505186 150226
rect 505296 150210 505324 158782
rect 506768 158778 506796 163200
rect 507596 158846 507624 163200
rect 508320 158908 508372 158914
rect 508320 158850 508372 158856
rect 507584 158840 507636 158846
rect 507584 158782 507636 158788
rect 505744 158772 505796 158778
rect 505744 158714 505796 158720
rect 506756 158772 506808 158778
rect 506756 158714 506808 158720
rect 507032 158772 507084 158778
rect 507032 158714 507084 158720
rect 505756 150226 505784 158714
rect 507044 150226 507072 158714
rect 507768 151904 507820 151910
rect 507768 151846 507820 151852
rect 507780 150226 507808 151846
rect 503226 149940 503254 150198
rect 503870 149940 503898 150198
rect 504514 149940 504542 150198
rect 505158 149940 505186 150198
rect 505284 150204 505336 150210
rect 505756 150198 505830 150226
rect 505284 150146 505336 150152
rect 505802 149940 505830 150198
rect 506434 150204 506486 150210
rect 507044 150198 507118 150226
rect 506434 150146 506486 150152
rect 506446 149940 506474 150146
rect 507090 149940 507118 150198
rect 507734 150198 507808 150226
rect 508332 150226 508360 158850
rect 508424 158778 508452 163200
rect 509252 163146 509280 163200
rect 509344 163146 509372 163254
rect 509252 163118 509372 163146
rect 508412 158772 508464 158778
rect 508412 158714 508464 158720
rect 509424 158772 509476 158778
rect 509424 158714 509476 158720
rect 509056 151972 509108 151978
rect 509056 151914 509108 151920
rect 509068 150226 509096 151914
rect 509436 151814 509464 158714
rect 509528 151910 509556 163254
rect 510066 163200 510122 164400
rect 510894 163200 510950 164400
rect 511722 163200 511778 164400
rect 512012 163254 512592 163282
rect 510080 158914 510108 163200
rect 510068 158908 510120 158914
rect 510068 158850 510120 158856
rect 510344 152856 510396 152862
rect 510344 152798 510396 152804
rect 509516 151904 509568 151910
rect 509516 151846 509568 151852
rect 509436 151786 509648 151814
rect 508332 150198 508406 150226
rect 507734 149940 507762 150198
rect 508378 149940 508406 150198
rect 509022 150198 509096 150226
rect 509620 150226 509648 151786
rect 510356 150226 510384 152798
rect 510908 151978 510936 163200
rect 511736 158778 511764 163200
rect 511724 158772 511776 158778
rect 511724 158714 511776 158720
rect 510988 153128 511040 153134
rect 510988 153070 511040 153076
rect 510896 151972 510948 151978
rect 510896 151914 510948 151920
rect 511000 150226 511028 153070
rect 512012 152862 512040 163254
rect 512564 163146 512592 163254
rect 512642 163200 512698 164400
rect 513470 163200 513526 164400
rect 513760 163254 514248 163282
rect 512656 163146 512684 163200
rect 512564 163118 512684 163146
rect 512920 153196 512972 153202
rect 512920 153138 512972 153144
rect 512276 152992 512328 152998
rect 512276 152934 512328 152940
rect 512000 152856 512052 152862
rect 512000 152798 512052 152804
rect 511632 152788 511684 152794
rect 511632 152730 511684 152736
rect 511644 150226 511672 152730
rect 512288 150226 512316 152934
rect 512932 150226 512960 153138
rect 513484 153134 513512 163200
rect 513472 153128 513524 153134
rect 513472 153070 513524 153076
rect 513564 152924 513616 152930
rect 513564 152866 513616 152872
rect 513576 150226 513604 152866
rect 513760 152794 513788 163254
rect 514220 163146 514248 163254
rect 514298 163200 514354 164400
rect 514772 163254 515076 163282
rect 514312 163146 514340 163200
rect 514220 163118 514340 163146
rect 514208 153128 514260 153134
rect 514208 153070 514260 153076
rect 513748 152788 513800 152794
rect 513748 152730 513800 152736
rect 514220 150226 514248 153070
rect 514772 152998 514800 163254
rect 515048 163146 515076 163254
rect 515126 163200 515182 164400
rect 515232 163254 515904 163282
rect 515140 163146 515168 163200
rect 515048 163118 515168 163146
rect 514944 158772 514996 158778
rect 514944 158714 514996 158720
rect 514760 152992 514812 152998
rect 514760 152934 514812 152940
rect 514956 151814 514984 158714
rect 515232 153202 515260 163254
rect 515876 163146 515904 163254
rect 515954 163200 516010 164400
rect 516152 163254 516732 163282
rect 515968 163146 515996 163200
rect 515876 163118 515996 163146
rect 515220 153196 515272 153202
rect 515220 153138 515272 153144
rect 516152 152930 516180 163254
rect 516704 163146 516732 163254
rect 516782 163200 516838 164400
rect 517610 163200 517666 164400
rect 518530 163200 518586 164400
rect 519004 163254 519308 163282
rect 516796 163146 516824 163200
rect 516704 163118 516824 163146
rect 517624 161474 517652 163200
rect 517532 161446 517652 161474
rect 517532 158794 517560 161446
rect 517440 158766 517560 158794
rect 518544 158778 518572 163200
rect 518808 159452 518860 159458
rect 518808 159394 518860 159400
rect 518716 159384 518768 159390
rect 518716 159326 518768 159332
rect 518532 158772 518584 158778
rect 517440 153134 517468 158766
rect 518532 158714 518584 158720
rect 517428 153128 517480 153134
rect 517428 153070 517480 153076
rect 516140 152924 516192 152930
rect 516140 152866 516192 152872
rect 516692 152040 516744 152046
rect 516692 151982 516744 151988
rect 515496 151972 515548 151978
rect 515496 151914 515548 151920
rect 514864 151786 514984 151814
rect 514864 150226 514892 151786
rect 515508 150226 515536 151914
rect 516048 151904 516100 151910
rect 516048 151846 516100 151852
rect 509620 150198 509694 150226
rect 509022 149940 509050 150198
rect 509666 149940 509694 150198
rect 510310 150198 510384 150226
rect 510954 150198 511028 150226
rect 511598 150198 511672 150226
rect 512242 150198 512316 150226
rect 512886 150198 512960 150226
rect 513530 150198 513604 150226
rect 514174 150198 514248 150226
rect 514818 150198 514892 150226
rect 515462 150198 515536 150226
rect 516060 150226 516088 151846
rect 516704 150226 516732 151982
rect 517428 151836 517480 151842
rect 517428 151778 517480 151784
rect 517440 150226 517468 151778
rect 518728 150226 518756 159326
rect 516060 150198 516134 150226
rect 516704 150198 516778 150226
rect 510310 149940 510338 150198
rect 510954 149940 510982 150198
rect 511598 149940 511626 150198
rect 512242 149940 512270 150198
rect 512886 149940 512914 150198
rect 513530 149940 513558 150198
rect 514174 149940 514202 150198
rect 514818 149940 514846 150198
rect 515462 149940 515490 150198
rect 516106 149940 516134 150198
rect 516750 149940 516778 150198
rect 517394 150198 517468 150226
rect 518026 150204 518078 150210
rect 517394 149940 517422 150198
rect 518026 150146 518078 150152
rect 518682 150198 518756 150226
rect 518820 150210 518848 159394
rect 519004 151978 519032 163254
rect 519280 163146 519308 163254
rect 519358 163200 519414 164400
rect 519924 163254 520136 163282
rect 519372 163146 519400 163200
rect 519280 163118 519400 163146
rect 519726 163160 519782 163169
rect 519726 163095 519782 163104
rect 519542 161664 519598 161673
rect 519542 161599 519598 161608
rect 519358 158672 519414 158681
rect 519358 158607 519414 158616
rect 518992 151972 519044 151978
rect 518992 151914 519044 151920
rect 518808 150204 518860 150210
rect 518038 149940 518066 150146
rect 518682 149940 518710 150198
rect 518808 150146 518860 150152
rect 519372 145761 519400 158607
rect 519556 148481 519584 161599
rect 519634 160168 519690 160177
rect 519634 160103 519690 160112
rect 519542 148472 519598 148481
rect 519542 148407 519598 148416
rect 519648 147121 519676 160103
rect 519740 149841 519768 163095
rect 519924 151910 519952 163254
rect 520108 163146 520136 163254
rect 520186 163200 520242 164400
rect 520292 163254 520964 163282
rect 520200 163146 520228 163200
rect 520108 163118 520228 163146
rect 520002 157176 520058 157185
rect 520002 157111 520058 157120
rect 519912 151904 519964 151910
rect 519912 151846 519964 151852
rect 519818 151192 519874 151201
rect 519818 151127 519874 151136
rect 519726 149832 519782 149841
rect 519726 149767 519782 149776
rect 519726 148200 519782 148209
rect 519726 148135 519782 148144
rect 519634 147112 519690 147121
rect 519634 147047 519690 147056
rect 519358 145752 519414 145761
rect 519358 145687 519414 145696
rect 519542 145208 519598 145217
rect 519542 145143 519598 145152
rect 519266 140584 519322 140593
rect 519266 140519 519322 140528
rect 519280 129441 519308 140519
rect 519358 139088 519414 139097
rect 519358 139023 519414 139032
rect 519266 129432 519322 129441
rect 519266 129367 519322 129376
rect 519372 128081 519400 139023
rect 519450 137456 519506 137465
rect 519450 137391 519506 137400
rect 519358 128072 519414 128081
rect 519358 128007 519414 128016
rect 519464 126721 519492 137391
rect 519556 133521 519584 145143
rect 519634 142216 519690 142225
rect 519634 142151 519690 142160
rect 519542 133512 519598 133521
rect 519542 133447 519598 133456
rect 519542 131608 519598 131617
rect 519542 131543 519598 131552
rect 519450 126712 519506 126721
rect 519450 126647 519506 126656
rect 519266 122496 519322 122505
rect 519266 122431 519322 122440
rect 117240 113206 117360 113234
rect 117332 113174 117360 113206
rect 117240 113146 117360 113174
rect 117240 107409 117268 113146
rect 519280 113121 519308 122431
rect 519556 121281 519584 131543
rect 519648 130801 519676 142151
rect 519740 136241 519768 148135
rect 519832 138961 519860 151127
rect 519910 149696 519966 149705
rect 519910 149631 519966 149640
rect 519818 138952 519874 138961
rect 519818 138887 519874 138896
rect 519924 137601 519952 149631
rect 520016 144401 520044 157111
rect 520094 155680 520150 155689
rect 520094 155615 520150 155624
rect 520002 144392 520058 144401
rect 520002 144327 520058 144336
rect 520108 143041 520136 155615
rect 520186 154184 520242 154193
rect 520186 154119 520242 154128
rect 520094 143032 520150 143041
rect 520094 142967 520150 142976
rect 520200 141681 520228 154119
rect 520292 152046 520320 163254
rect 520936 163146 520964 163254
rect 521014 163200 521070 164400
rect 521842 163200 521898 164400
rect 522670 163200 522726 164400
rect 523498 163200 523554 164400
rect 521028 163146 521056 163200
rect 520936 163118 521056 163146
rect 521856 161474 521884 163200
rect 521672 161446 521884 161474
rect 521672 158794 521700 161446
rect 522684 159458 522712 163200
rect 522672 159452 522724 159458
rect 522672 159394 522724 159400
rect 523512 159390 523540 163200
rect 523500 159384 523552 159390
rect 523500 159326 523552 159332
rect 521580 158766 521700 158794
rect 521106 152688 521162 152697
rect 521106 152623 521162 152632
rect 520280 152040 520332 152046
rect 520280 151982 520332 151988
rect 521014 146704 521070 146713
rect 521014 146639 521070 146648
rect 520922 143712 520978 143721
rect 520922 143647 520978 143656
rect 520186 141672 520242 141681
rect 520186 141607 520242 141616
rect 519910 137592 519966 137601
rect 519910 137527 519966 137536
rect 519726 136232 519782 136241
rect 519726 136167 519782 136176
rect 520186 136096 520242 136105
rect 520186 136031 520242 136040
rect 520002 134600 520058 134609
rect 520002 134535 520058 134544
rect 519634 130792 519690 130801
rect 519634 130727 519690 130736
rect 519818 130112 519874 130121
rect 519818 130047 519874 130056
rect 519634 128616 519690 128625
rect 519634 128551 519690 128560
rect 519542 121272 519598 121281
rect 519542 121207 519598 121216
rect 519358 121136 519414 121145
rect 519358 121071 519414 121080
rect 519266 113112 519322 113121
rect 519266 113047 519322 113056
rect 519372 111761 519400 121071
rect 519450 119640 519506 119649
rect 519450 119575 519506 119584
rect 519358 111752 519414 111761
rect 519358 111687 519414 111696
rect 519464 110401 519492 119575
rect 519648 118561 519676 128551
rect 519726 127120 519782 127129
rect 519726 127055 519782 127064
rect 519634 118552 519690 118561
rect 519634 118487 519690 118496
rect 519740 117201 519768 127055
rect 519832 119921 519860 130047
rect 519910 125624 519966 125633
rect 519910 125559 519966 125568
rect 519818 119912 519874 119921
rect 519818 119847 519874 119856
rect 519818 118144 519874 118153
rect 519818 118079 519874 118088
rect 519726 117192 519782 117201
rect 519726 117127 519782 117136
rect 519726 113520 519782 113529
rect 519726 113455 519782 113464
rect 519634 112024 519690 112033
rect 519634 111959 519690 111968
rect 519542 110528 519598 110537
rect 519542 110463 519598 110472
rect 519450 110392 519506 110401
rect 519450 110327 519506 110336
rect 117226 107400 117282 107409
rect 117226 107335 117282 107344
rect 117134 104544 117190 104553
rect 117134 104479 117190 104488
rect 117042 103184 117098 103193
rect 117042 103119 117098 103128
rect 519556 102105 519584 110463
rect 519648 103465 519676 111959
rect 519740 104825 519768 113455
rect 519832 109041 519860 118079
rect 519924 115569 519952 125559
rect 520016 124001 520044 134535
rect 520094 133104 520150 133113
rect 520094 133039 520150 133048
rect 520002 123992 520058 124001
rect 520002 123927 520058 123936
rect 520108 122641 520136 133039
rect 520200 125225 520228 136031
rect 520936 132161 520964 143647
rect 521028 134745 521056 146639
rect 521120 140321 521148 152623
rect 521580 151842 521608 158766
rect 521568 151836 521620 151842
rect 521568 151778 521620 151784
rect 521106 140312 521162 140321
rect 521106 140247 521162 140256
rect 521014 134736 521070 134745
rect 521014 134671 521070 134680
rect 520922 132152 520978 132161
rect 520922 132087 520978 132096
rect 520186 125216 520242 125225
rect 520186 125151 520242 125160
rect 520186 124128 520242 124137
rect 520186 124063 520242 124072
rect 520094 122632 520150 122641
rect 520094 122567 520150 122576
rect 520002 116512 520058 116521
rect 520002 116447 520058 116456
rect 519910 115560 519966 115569
rect 519910 115495 519966 115504
rect 519818 109032 519874 109041
rect 519818 108967 519874 108976
rect 520016 107545 520044 116447
rect 520094 115016 520150 115025
rect 520094 114951 520150 114960
rect 520002 107536 520058 107545
rect 520002 107471 520058 107480
rect 520108 106049 520136 114951
rect 520200 114481 520228 124063
rect 520186 114472 520242 114481
rect 520186 114407 520242 114416
rect 520830 109032 520886 109041
rect 520830 108967 520886 108976
rect 520094 106040 520150 106049
rect 520094 105975 520150 105984
rect 520278 106040 520334 106049
rect 520278 105975 520334 105984
rect 519726 104816 519782 104825
rect 519726 104751 519782 104760
rect 519634 103456 519690 103465
rect 519634 103391 519690 103400
rect 519542 102096 519598 102105
rect 519542 102031 519598 102040
rect 116950 101552 117006 101561
rect 116950 101487 117006 101496
rect 116858 99376 116914 99385
rect 116858 99311 116914 99320
rect 520292 97889 520320 105975
rect 520738 103048 520794 103057
rect 520738 102983 520794 102992
rect 520278 97880 520334 97889
rect 520278 97815 520334 97824
rect 116766 97744 116822 97753
rect 116766 97679 116822 97688
rect 116674 95840 116730 95849
rect 116674 95775 116730 95784
rect 520278 95568 520334 95577
rect 520278 95503 520334 95512
rect 116582 93664 116638 93673
rect 116582 93599 116638 93608
rect 115940 92472 115992 92478
rect 115940 92414 115992 92420
rect 115952 91905 115980 92414
rect 519726 92304 519782 92313
rect 519726 92239 519782 92248
rect 115938 91896 115994 91905
rect 115938 91831 115994 91840
rect 116124 89684 116176 89690
rect 116124 89626 116176 89632
rect 116136 89593 116164 89626
rect 116122 89584 116178 89593
rect 116122 89519 116178 89528
rect 115940 88324 115992 88330
rect 115940 88266 115992 88272
rect 115952 88097 115980 88266
rect 115938 88088 115994 88097
rect 115938 88023 115994 88032
rect 114468 87032 114520 87038
rect 114466 87000 114468 87009
rect 116676 87032 116728 87038
rect 114520 87000 114522 87009
rect 116676 86974 116728 86980
rect 114466 86935 114522 86944
rect 116032 86964 116084 86970
rect 116032 86906 116084 86912
rect 116044 86193 116072 86906
rect 116030 86184 116086 86193
rect 116030 86119 116086 86128
rect 116584 83972 116636 83978
rect 116584 83914 116636 83920
rect 116596 83881 116624 83914
rect 116582 83872 116638 83881
rect 116582 83807 116638 83816
rect 116124 82816 116176 82822
rect 116124 82758 116176 82764
rect 116136 82385 116164 82758
rect 116122 82376 116178 82385
rect 116122 82311 116178 82320
rect 115938 80064 115994 80073
rect 114192 80028 114244 80034
rect 115938 79999 115940 80008
rect 114192 79970 114244 79976
rect 115992 79999 115994 80008
rect 115940 79970 115992 79976
rect 116688 78577 116716 86974
rect 519634 86456 519690 86465
rect 519634 86391 519690 86400
rect 519266 81968 519322 81977
rect 519266 81903 519322 81912
rect 116674 78568 116730 78577
rect 116674 78503 116730 78512
rect 519280 76537 519308 81903
rect 519648 80073 519676 86391
rect 519740 85513 519768 92239
rect 520094 90944 520150 90953
rect 520094 90879 520150 90888
rect 520002 89448 520058 89457
rect 520002 89383 520058 89392
rect 519818 87952 519874 87961
rect 519818 87887 519874 87896
rect 519726 85504 519782 85513
rect 519726 85439 519782 85448
rect 519726 84960 519782 84969
rect 519726 84895 519782 84904
rect 519634 80064 519690 80073
rect 519634 79999 519690 80008
rect 519740 78305 519768 84895
rect 519832 81433 519860 87887
rect 520016 82793 520044 89383
rect 520108 84153 520136 90879
rect 520292 88233 520320 95503
rect 520752 95169 520780 102983
rect 520844 100745 520872 108967
rect 520922 107536 520978 107545
rect 520922 107471 520978 107480
rect 520830 100736 520886 100745
rect 520830 100671 520886 100680
rect 520936 99385 520964 107471
rect 521014 104544 521070 104553
rect 521014 104479 521070 104488
rect 520922 99376 520978 99385
rect 520922 99311 520978 99320
rect 521028 96393 521056 104479
rect 521198 101552 521254 101561
rect 521198 101487 521254 101496
rect 521014 96384 521070 96393
rect 521014 96319 521070 96328
rect 520738 95160 520794 95169
rect 520738 95095 520794 95104
rect 520922 93936 520978 93945
rect 520922 93871 520978 93880
rect 520278 88224 520334 88233
rect 520278 88159 520334 88168
rect 520936 86873 520964 93871
rect 521212 93809 521240 101487
rect 521474 100056 521530 100065
rect 521474 99991 521530 100000
rect 521382 98560 521438 98569
rect 521382 98495 521438 98504
rect 521198 93800 521254 93809
rect 521198 93735 521254 93744
rect 521396 91089 521424 98495
rect 521488 92449 521516 99991
rect 521566 97064 521622 97073
rect 521566 96999 521622 97008
rect 521474 92440 521530 92449
rect 521474 92375 521530 92384
rect 521382 91080 521438 91089
rect 521382 91015 521438 91024
rect 521580 89729 521608 96999
rect 521566 89720 521622 89729
rect 521566 89655 521622 89664
rect 520922 86864 520978 86873
rect 520922 86799 520978 86808
rect 520094 84144 520150 84153
rect 520094 84079 520150 84088
rect 520094 83464 520150 83473
rect 520094 83399 520150 83408
rect 520002 82784 520058 82793
rect 520002 82719 520058 82728
rect 519818 81424 519874 81433
rect 519818 81359 519874 81368
rect 519910 78976 519966 78985
rect 519910 78911 519966 78920
rect 519726 78296 519782 78305
rect 519726 78231 519782 78240
rect 519818 77480 519874 77489
rect 519818 77415 519874 77424
rect 519266 76528 519322 76537
rect 519266 76463 519322 76472
rect 519726 75984 519782 75993
rect 519726 75919 519782 75928
rect 116674 73536 116730 73545
rect 116674 73471 116730 73480
rect 116030 71904 116086 71913
rect 116030 71839 116086 71848
rect 116044 71806 116072 71839
rect 114192 71800 114244 71806
rect 114192 71742 114244 71748
rect 116032 71800 116084 71806
rect 116032 71742 116084 71748
rect 114100 69080 114152 69086
rect 114100 69022 114152 69028
rect 114008 67652 114060 67658
rect 114008 67594 114060 67600
rect 113916 66292 113968 66298
rect 113916 66234 113968 66240
rect 113824 63572 113876 63578
rect 113824 63514 113876 63520
rect 109684 41472 109736 41478
rect 109684 41414 109736 41420
rect 109592 3052 109644 3058
rect 109592 2994 109644 3000
rect 2504 2916 2556 2922
rect 2504 2858 2556 2864
rect 2516 2666 2544 2858
rect 109604 2689 109632 2994
rect 45650 2680 45706 2689
rect 2516 2638 2714 2666
rect 40684 2644 40736 2650
rect 40684 2586 40736 2592
rect 43628 2644 43680 2650
rect 49974 2680 50030 2689
rect 49358 2650 49648 2666
rect 49358 2644 49660 2650
rect 49358 2638 49608 2644
rect 45650 2615 45652 2624
rect 43628 2586 43680 2592
rect 45704 2615 45706 2624
rect 45652 2586 45704 2592
rect 49608 2586 49660 2592
rect 49792 2644 49844 2650
rect 49792 2586 49844 2592
rect 49884 2644 49936 2650
rect 66258 2680 66314 2689
rect 59386 2650 59768 2666
rect 53932 2644 53984 2650
rect 49974 2615 49976 2624
rect 49884 2586 49936 2592
rect 50028 2615 50030 2624
rect 49976 2586 50028 2592
rect 53668 2604 53932 2632
rect 32772 2576 32824 2582
rect 32772 2518 32824 2524
rect 6012 1426 6040 2108
rect 9324 1465 9352 2108
rect 12636 1601 12664 2108
rect 15948 1737 15976 2108
rect 19352 1873 19380 2108
rect 19338 1864 19394 1873
rect 19338 1799 19394 1808
rect 15934 1728 15990 1737
rect 15934 1663 15990 1672
rect 12622 1592 12678 1601
rect 12622 1527 12678 1536
rect 22664 1494 22692 2108
rect 25976 1562 26004 2108
rect 29288 1630 29316 2108
rect 32692 1698 32720 2108
rect 32680 1692 32732 1698
rect 32680 1634 32732 1640
rect 29276 1624 29328 1630
rect 29276 1566 29328 1572
rect 25964 1556 26016 1562
rect 25964 1498 26016 1504
rect 22652 1488 22704 1494
rect 9310 1456 9366 1465
rect 6000 1420 6052 1426
rect 22652 1430 22704 1436
rect 9310 1391 9366 1400
rect 6000 1362 6052 1368
rect 32784 800 32812 2518
rect 40696 2514 40724 2586
rect 40684 2508 40736 2514
rect 40684 2450 40736 2456
rect 39672 2440 39724 2446
rect 36018 2378 36400 2394
rect 39330 2388 39672 2394
rect 39330 2382 39724 2388
rect 36018 2372 36412 2378
rect 36018 2366 36360 2372
rect 39330 2366 39712 2382
rect 43640 2378 43668 2586
rect 46046 2378 46336 2394
rect 49804 2378 49832 2586
rect 43628 2372 43680 2378
rect 36360 2314 36412 2320
rect 46046 2372 46348 2378
rect 46046 2366 46296 2372
rect 43628 2314 43680 2320
rect 46296 2314 46348 2320
rect 49792 2372 49844 2378
rect 49792 2314 49844 2320
rect 49896 2310 49924 2586
rect 53668 2446 53696 2604
rect 53932 2586 53984 2592
rect 58992 2644 59044 2650
rect 59386 2644 59780 2650
rect 59386 2638 59728 2644
rect 58992 2586 59044 2592
rect 59728 2586 59780 2592
rect 59820 2644 59872 2650
rect 84566 2680 84622 2689
rect 66258 2615 66314 2624
rect 67548 2644 67600 2650
rect 59820 2586 59872 2592
rect 53656 2440 53708 2446
rect 56232 2440 56284 2446
rect 53656 2382 53708 2388
rect 55982 2388 56232 2394
rect 55982 2382 56284 2388
rect 55982 2366 56272 2382
rect 59004 2310 59032 2586
rect 59832 2378 59860 2586
rect 64878 2544 64934 2553
rect 64878 2479 64880 2488
rect 64932 2479 64934 2488
rect 64880 2450 64932 2456
rect 59820 2372 59872 2378
rect 59820 2314 59872 2320
rect 42984 2304 43036 2310
rect 42642 2252 42984 2258
rect 42642 2246 43036 2252
rect 49884 2304 49936 2310
rect 52920 2304 52972 2310
rect 49884 2246 49936 2252
rect 52670 2252 52920 2258
rect 52670 2246 52972 2252
rect 58992 2304 59044 2310
rect 66272 2258 66300 2615
rect 67548 2586 67600 2592
rect 68836 2644 68888 2650
rect 68836 2586 68888 2592
rect 68928 2644 68980 2650
rect 68928 2586 68980 2592
rect 69020 2644 69072 2650
rect 69020 2586 69072 2592
rect 69848 2644 69900 2650
rect 69848 2586 69900 2592
rect 70676 2644 70728 2650
rect 70676 2586 70728 2592
rect 72424 2644 72476 2650
rect 72424 2586 72476 2592
rect 72516 2644 72568 2650
rect 72516 2586 72568 2592
rect 75000 2644 75052 2650
rect 75000 2586 75052 2592
rect 76288 2644 76340 2650
rect 76288 2586 76340 2592
rect 76472 2644 76524 2650
rect 76472 2586 76524 2592
rect 84016 2644 84068 2650
rect 84016 2586 84068 2592
rect 84476 2644 84528 2650
rect 106094 2680 106150 2689
rect 84566 2615 84568 2624
rect 84476 2586 84528 2592
rect 84620 2615 84622 2624
rect 84752 2644 84804 2650
rect 84568 2586 84620 2592
rect 84752 2586 84804 2592
rect 85304 2644 85356 2650
rect 85304 2586 85356 2592
rect 85856 2644 85908 2650
rect 85856 2586 85908 2592
rect 98276 2644 98328 2650
rect 106094 2615 106096 2624
rect 98276 2586 98328 2592
rect 106148 2615 106150 2624
rect 109590 2680 109646 2689
rect 109590 2615 109646 2624
rect 106096 2586 106148 2592
rect 67560 2417 67588 2586
rect 68848 2446 68876 2586
rect 68836 2440 68888 2446
rect 67546 2408 67602 2417
rect 68836 2382 68888 2388
rect 67546 2343 67602 2352
rect 68940 2310 68968 2586
rect 58992 2246 59044 2252
rect 42642 2230 43024 2246
rect 52670 2230 52960 2246
rect 66010 2230 66300 2258
rect 68928 2304 68980 2310
rect 69032 2281 69060 2586
rect 68928 2246 68980 2252
rect 69018 2272 69074 2281
rect 69322 2242 69704 2258
rect 69322 2236 69716 2242
rect 69322 2230 69664 2236
rect 69018 2207 69074 2216
rect 69664 2178 69716 2184
rect 69860 2174 69888 2586
rect 63040 2168 63092 2174
rect 62698 2116 63040 2122
rect 62698 2110 63092 2116
rect 69848 2168 69900 2174
rect 69848 2110 69900 2116
rect 62698 2094 63080 2110
rect 70688 2106 70716 2586
rect 70676 2100 70728 2106
rect 70676 2042 70728 2048
rect 72436 2038 72464 2586
rect 72528 2514 72556 2586
rect 72516 2508 72568 2514
rect 72516 2450 72568 2456
rect 72424 2032 72476 2038
rect 72424 1974 72476 1980
rect 72712 1834 72740 2108
rect 75012 2106 75040 2586
rect 76300 2174 76328 2586
rect 76484 2281 76512 2586
rect 76564 2576 76616 2582
rect 76564 2518 76616 2524
rect 76576 2378 76604 2518
rect 84028 2446 84056 2586
rect 84016 2440 84068 2446
rect 84016 2382 84068 2388
rect 76564 2372 76616 2378
rect 76564 2314 76616 2320
rect 84488 2310 84516 2586
rect 84476 2304 84528 2310
rect 76470 2272 76526 2281
rect 84476 2246 84528 2252
rect 84764 2242 84792 2586
rect 85316 2417 85344 2586
rect 85868 2553 85896 2586
rect 85854 2544 85910 2553
rect 85854 2479 85910 2488
rect 85302 2408 85358 2417
rect 85302 2343 85358 2352
rect 96002 2242 96384 2258
rect 76470 2207 76526 2216
rect 84752 2236 84804 2242
rect 96002 2236 96396 2242
rect 96002 2230 96344 2236
rect 84752 2178 84804 2184
rect 96344 2178 96396 2184
rect 76288 2168 76340 2174
rect 93032 2168 93084 2174
rect 76288 2110 76340 2116
rect 75000 2100 75052 2106
rect 75000 2042 75052 2048
rect 72700 1828 72752 1834
rect 72700 1770 72752 1776
rect 76024 1766 76052 2108
rect 79336 1902 79364 2108
rect 82648 1970 82676 2108
rect 86066 2094 86448 2122
rect 89378 2106 89668 2122
rect 92690 2116 93032 2122
rect 92690 2110 93084 2116
rect 89378 2100 89680 2106
rect 89378 2094 89628 2100
rect 86420 2038 86448 2094
rect 92690 2094 93072 2110
rect 89628 2042 89680 2048
rect 86408 2032 86460 2038
rect 86408 1974 86460 1980
rect 82636 1964 82688 1970
rect 82636 1906 82688 1912
rect 79324 1896 79376 1902
rect 79324 1838 79376 1844
rect 76012 1760 76064 1766
rect 76012 1702 76064 1708
rect 98288 800 98316 2586
rect 109342 2514 109632 2530
rect 109342 2508 109644 2514
rect 109342 2502 109592 2508
rect 109592 2450 109644 2456
rect 106188 2440 106240 2446
rect 102718 2378 103008 2394
rect 106030 2388 106188 2394
rect 106030 2382 106240 2388
rect 102718 2372 103020 2378
rect 102718 2366 102968 2372
rect 106030 2366 106228 2382
rect 102968 2314 103020 2320
rect 99656 2304 99708 2310
rect 99406 2252 99656 2258
rect 99406 2246 99708 2252
rect 99406 2230 99696 2246
rect 109696 1834 109724 41414
rect 111064 34536 111116 34542
rect 111064 34478 111116 34484
rect 109776 4208 109828 4214
rect 109776 4150 109828 4156
rect 109684 1828 109736 1834
rect 109684 1770 109736 1776
rect 109788 1426 109816 4150
rect 111076 3942 111104 34478
rect 112444 33176 112496 33182
rect 112444 33118 112496 33124
rect 111156 23520 111208 23526
rect 111156 23462 111208 23468
rect 111064 3936 111116 3942
rect 111064 3878 111116 3884
rect 111168 3534 111196 23462
rect 111248 22160 111300 22166
rect 111248 22102 111300 22108
rect 111156 3528 111208 3534
rect 111156 3470 111208 3476
rect 111260 3466 111288 22102
rect 112456 3874 112484 33118
rect 112536 31816 112588 31822
rect 112536 31758 112588 31764
rect 112444 3868 112496 3874
rect 112444 3810 112496 3816
rect 112548 3806 112576 31758
rect 112628 29028 112680 29034
rect 112628 28970 112680 28976
rect 112536 3800 112588 3806
rect 112536 3742 112588 3748
rect 112640 3738 112668 28970
rect 112720 27668 112772 27674
rect 112720 27610 112772 27616
rect 112628 3732 112680 3738
rect 112628 3674 112680 3680
rect 112732 3670 112760 27610
rect 112812 24880 112864 24886
rect 112812 24822 112864 24828
rect 112720 3664 112772 3670
rect 112720 3606 112772 3612
rect 112824 3602 112852 24822
rect 113836 8265 113864 63514
rect 113928 19145 113956 66234
rect 114020 30977 114048 67594
rect 114112 42401 114140 69022
rect 114204 53689 114232 71742
rect 116214 69728 116270 69737
rect 116214 69663 116270 69672
rect 116228 69086 116256 69663
rect 116216 69080 116268 69086
rect 116216 69022 116268 69028
rect 115938 67824 115994 67833
rect 115938 67759 115994 67768
rect 115952 67658 115980 67759
rect 115940 67652 115992 67658
rect 115940 67594 115992 67600
rect 116582 66600 116638 66609
rect 116582 66535 116638 66544
rect 116596 66298 116624 66535
rect 116584 66292 116636 66298
rect 116584 66234 116636 66240
rect 116688 64874 116716 73471
rect 519740 71097 519768 75919
rect 519832 72457 519860 77415
rect 519924 73817 519952 78911
rect 520108 76945 520136 83399
rect 520186 80472 520242 80481
rect 520186 80407 520242 80416
rect 520094 76936 520150 76945
rect 520094 76871 520150 76880
rect 520200 75177 520228 80407
rect 520186 75168 520242 75177
rect 520186 75103 520242 75112
rect 521198 74488 521254 74497
rect 521198 74423 521254 74432
rect 519910 73808 519966 73817
rect 519910 73743 519966 73752
rect 521014 72992 521070 73001
rect 521014 72927 521070 72936
rect 519818 72448 519874 72457
rect 519818 72383 519874 72392
rect 519726 71088 519782 71097
rect 519726 71023 519782 71032
rect 520738 69864 520794 69873
rect 520738 69799 520794 69808
rect 520462 66872 520518 66881
rect 520462 66807 520518 66816
rect 520370 65376 520426 65385
rect 520370 65311 520426 65320
rect 116596 64846 116716 64874
rect 116596 64734 116624 64846
rect 114468 64728 114520 64734
rect 114466 64696 114468 64705
rect 116584 64728 116636 64734
rect 114520 64696 114522 64705
rect 116584 64670 116636 64676
rect 114466 64631 114522 64640
rect 116030 64016 116086 64025
rect 116030 63951 116086 63960
rect 116044 63578 116072 63951
rect 116032 63572 116084 63578
rect 116032 63514 116084 63520
rect 116582 62248 116638 62257
rect 116582 62183 116638 62192
rect 114190 53680 114246 53689
rect 114190 53615 114246 53624
rect 116490 47288 116546 47297
rect 116490 47223 116546 47232
rect 116214 44704 116270 44713
rect 116214 44639 116270 44648
rect 114098 42392 114154 42401
rect 114098 42327 114154 42336
rect 116122 41576 116178 41585
rect 116122 41511 116178 41520
rect 116136 41478 116164 41511
rect 116124 41472 116176 41478
rect 116124 41414 116176 41420
rect 114100 38684 114152 38690
rect 114100 38626 114152 38632
rect 114006 30968 114062 30977
rect 114006 30903 114062 30912
rect 113914 19136 113970 19145
rect 113914 19071 113970 19080
rect 113822 8256 113878 8265
rect 113822 8191 113878 8200
rect 112812 3596 112864 3602
rect 112812 3538 112864 3544
rect 111248 3460 111300 3466
rect 111248 3402 111300 3408
rect 114112 3330 114140 38626
rect 116228 38554 116256 44639
rect 116306 42936 116362 42945
rect 116306 42871 116362 42880
rect 116216 38548 116268 38554
rect 116216 38490 116268 38496
rect 115938 37360 115994 37369
rect 114192 37324 114244 37330
rect 115938 37295 115940 37304
rect 114192 37266 114244 37272
rect 115992 37295 115994 37304
rect 115940 37266 115992 37272
rect 114204 3398 114232 37266
rect 116122 35184 116178 35193
rect 116122 35119 116178 35128
rect 116136 34542 116164 35119
rect 116124 34536 116176 34542
rect 116124 34478 116176 34484
rect 116122 33280 116178 33289
rect 116122 33215 116178 33224
rect 116136 33182 116164 33215
rect 116124 33176 116176 33182
rect 116124 33118 116176 33124
rect 116122 31920 116178 31929
rect 116122 31855 116178 31864
rect 116136 31822 116164 31855
rect 116124 31816 116176 31822
rect 116124 31758 116176 31764
rect 116122 29336 116178 29345
rect 116122 29271 116178 29280
rect 116136 29034 116164 29271
rect 116124 29028 116176 29034
rect 116124 28970 116176 28976
rect 116122 27704 116178 27713
rect 116122 27639 116124 27648
rect 116176 27639 116178 27648
rect 116124 27610 116176 27616
rect 116122 25528 116178 25537
rect 116122 25463 116178 25472
rect 116136 24886 116164 25463
rect 116124 24880 116176 24886
rect 116124 24822 116176 24828
rect 116122 23624 116178 23633
rect 116122 23559 116178 23568
rect 116136 23526 116164 23559
rect 116124 23520 116176 23526
rect 116124 23462 116176 23468
rect 116122 22400 116178 22409
rect 116122 22335 116178 22344
rect 116136 22166 116164 22335
rect 116124 22160 116176 22166
rect 116124 22102 116176 22108
rect 116214 19816 116270 19825
rect 116214 19751 116270 19760
rect 116122 18048 116178 18057
rect 116122 17983 116178 17992
rect 116136 16574 116164 17983
rect 116044 16546 116164 16574
rect 115938 13968 115994 13977
rect 115938 13903 115994 13912
rect 115952 4706 115980 13903
rect 115860 4678 115980 4706
rect 115860 4026 115888 4678
rect 115938 4584 115994 4593
rect 115938 4519 115994 4528
rect 115952 4214 115980 4519
rect 115940 4208 115992 4214
rect 115940 4150 115992 4156
rect 115860 3998 115980 4026
rect 114192 3392 114244 3398
rect 114192 3334 114244 3340
rect 114100 3324 114152 3330
rect 114100 3266 114152 3272
rect 115848 2916 115900 2922
rect 115848 2858 115900 2864
rect 115860 2825 115888 2858
rect 115846 2816 115902 2825
rect 115846 2751 115902 2760
rect 115952 1494 115980 3998
rect 116044 1630 116072 16546
rect 116122 15872 116178 15881
rect 116122 15807 116178 15816
rect 116032 1624 116084 1630
rect 116032 1566 116084 1572
rect 116136 1562 116164 15807
rect 116228 1698 116256 19751
rect 116320 1766 116348 42871
rect 116398 38992 116454 39001
rect 116398 38927 116454 38936
rect 116412 38690 116440 38927
rect 116400 38684 116452 38690
rect 116400 38626 116452 38632
rect 116400 38548 116452 38554
rect 116400 38490 116452 38496
rect 116412 1902 116440 38490
rect 116504 1970 116532 47223
rect 116596 2514 116624 62183
rect 520384 61577 520412 65311
rect 520476 62937 520504 66807
rect 520752 65657 520780 69799
rect 521028 68377 521056 72927
rect 521106 71496 521162 71505
rect 521106 71431 521162 71440
rect 521014 68368 521070 68377
rect 521014 68303 521070 68312
rect 521120 67017 521148 71431
rect 521212 69737 521240 74423
rect 521198 69728 521254 69737
rect 521198 69663 521254 69672
rect 521198 68368 521254 68377
rect 521198 68303 521254 68312
rect 521106 67008 521162 67017
rect 521106 66943 521162 66952
rect 520738 65648 520794 65657
rect 520738 65583 520794 65592
rect 521212 64297 521240 68303
rect 521198 64288 521254 64297
rect 521198 64223 521254 64232
rect 521198 63880 521254 63889
rect 521198 63815 521254 63824
rect 520462 62928 520518 62937
rect 520462 62863 520518 62872
rect 521014 62384 521070 62393
rect 521014 62319 521070 62328
rect 520370 61568 520426 61577
rect 520370 61503 520426 61512
rect 116674 60072 116730 60081
rect 116674 60007 116730 60016
rect 116584 2508 116636 2514
rect 116584 2450 116636 2456
rect 116688 2446 116716 60007
rect 520554 59392 520610 59401
rect 520554 59327 520610 59336
rect 116766 58168 116822 58177
rect 116766 58103 116822 58112
rect 116676 2440 116728 2446
rect 116676 2382 116728 2388
rect 116780 2378 116808 58103
rect 519910 57896 519966 57905
rect 519910 57831 519966 57840
rect 116858 56944 116914 56953
rect 116858 56879 116914 56888
rect 116768 2372 116820 2378
rect 116768 2314 116820 2320
rect 116872 2310 116900 56879
rect 519266 56400 519322 56409
rect 519266 56335 519322 56344
rect 519082 54904 519138 54913
rect 519082 54839 519138 54848
rect 116950 54360 117006 54369
rect 116950 54295 117006 54304
rect 116860 2304 116912 2310
rect 116860 2246 116912 2252
rect 116964 2242 116992 54295
rect 117042 52592 117098 52601
rect 117042 52527 117098 52536
rect 116952 2236 117004 2242
rect 116952 2178 117004 2184
rect 117056 2174 117084 52527
rect 519096 52057 519124 54839
rect 519280 53417 519308 56335
rect 519924 54777 519952 57831
rect 520568 56137 520596 59327
rect 521028 58857 521056 62319
rect 521106 60888 521162 60897
rect 521106 60823 521162 60832
rect 521014 58848 521070 58857
rect 521014 58783 521070 58792
rect 521120 57497 521148 60823
rect 521212 60217 521240 63815
rect 521198 60208 521254 60217
rect 521198 60143 521254 60152
rect 521106 57488 521162 57497
rect 521106 57423 521162 57432
rect 520554 56128 520610 56137
rect 520554 56063 520610 56072
rect 519910 54768 519966 54777
rect 519910 54703 519966 54712
rect 519266 53408 519322 53417
rect 519266 53343 519322 53352
rect 520002 53408 520058 53417
rect 520002 53343 520058 53352
rect 519082 52048 519138 52057
rect 519082 51983 519138 51992
rect 117134 51232 117190 51241
rect 117134 51167 117190 51176
rect 117044 2168 117096 2174
rect 117044 2110 117096 2116
rect 117148 2106 117176 51167
rect 520016 50697 520044 53343
rect 520186 51912 520242 51921
rect 520186 51847 520242 51856
rect 520002 50688 520058 50697
rect 520002 50623 520058 50632
rect 520094 50416 520150 50425
rect 520094 50351 520150 50360
rect 117226 48648 117282 48657
rect 117226 48583 117282 48592
rect 117136 2100 117188 2106
rect 117136 2042 117188 2048
rect 117240 2038 117268 48583
rect 520108 47841 520136 50351
rect 520200 49337 520228 51847
rect 520186 49328 520242 49337
rect 520186 49263 520242 49272
rect 520186 48920 520242 48929
rect 520186 48855 520242 48864
rect 520094 47832 520150 47841
rect 520094 47767 520150 47776
rect 519910 47288 519966 47297
rect 519910 47223 519966 47232
rect 519818 45792 519874 45801
rect 519818 45727 519874 45736
rect 519832 43897 519860 45727
rect 519924 45257 519952 47223
rect 520200 46617 520228 48855
rect 520186 46608 520242 46617
rect 520186 46543 520242 46552
rect 519910 45248 519966 45257
rect 519910 45183 519966 45192
rect 520186 44296 520242 44305
rect 520186 44231 520242 44240
rect 519818 43888 519874 43897
rect 519818 43823 519874 43832
rect 520200 42537 520228 44231
rect 520738 42800 520794 42809
rect 520738 42735 520794 42744
rect 520186 42528 520242 42537
rect 520186 42463 520242 42472
rect 520752 41313 520780 42735
rect 520738 41304 520794 41313
rect 520738 41239 520794 41248
rect 520922 41304 520978 41313
rect 520922 41239 520978 41248
rect 520936 39953 520964 41239
rect 520922 39944 520978 39953
rect 520922 39879 520978 39888
rect 520370 39808 520426 39817
rect 520370 39743 520426 39752
rect 520384 38321 520412 39743
rect 520370 38312 520426 38321
rect 520370 38247 520426 38256
rect 520554 38312 520610 38321
rect 520554 38247 520610 38256
rect 520568 37233 520596 38247
rect 520554 37224 520610 37233
rect 520554 37159 520610 37168
rect 521566 36816 521622 36825
rect 521566 36751 521622 36760
rect 521580 36009 521608 36751
rect 521566 36000 521622 36009
rect 521566 35935 521622 35944
rect 520922 35320 520978 35329
rect 520922 35255 520978 35264
rect 520936 34513 520964 35255
rect 520922 34504 520978 34513
rect 520922 34439 520978 34448
rect 521106 33824 521162 33833
rect 521106 33759 521162 33768
rect 521120 33153 521148 33759
rect 521106 33144 521162 33153
rect 521106 33079 521162 33088
rect 521106 32328 521162 32337
rect 521106 32263 521162 32272
rect 521120 31657 521148 32263
rect 521106 31648 521162 31657
rect 521106 31583 521162 31592
rect 521106 29336 521162 29345
rect 521106 29271 521162 29280
rect 521120 28665 521148 29271
rect 521106 28656 521162 28665
rect 521106 28591 521162 28600
rect 521106 24848 521162 24857
rect 521106 24783 521162 24792
rect 521120 23633 521148 24783
rect 521106 23624 521162 23633
rect 521106 23559 521162 23568
rect 520922 23216 520978 23225
rect 520922 23151 520978 23160
rect 520936 22273 520964 23151
rect 520922 22264 520978 22273
rect 520922 22199 520978 22208
rect 520922 21720 520978 21729
rect 520922 21655 520978 21664
rect 520936 20913 520964 21655
rect 520922 20904 520978 20913
rect 520922 20839 520978 20848
rect 521106 20224 521162 20233
rect 521106 20159 521162 20168
rect 521120 19553 521148 20159
rect 521106 19544 521162 19553
rect 521106 19479 521162 19488
rect 520370 7440 520426 7449
rect 520370 7375 520426 7384
rect 520384 6769 520412 7375
rect 520370 6760 520426 6769
rect 520370 6695 520426 6704
rect 521106 6080 521162 6089
rect 521106 6015 521162 6024
rect 521120 5273 521148 6015
rect 521106 5264 521162 5273
rect 521106 5199 521162 5208
rect 521106 4720 521162 4729
rect 521106 4655 521162 4664
rect 521120 3777 521148 4655
rect 521106 3768 521162 3777
rect 521106 3703 521162 3712
rect 520922 3360 520978 3369
rect 520922 3295 520978 3304
rect 117964 3052 118016 3058
rect 117964 2994 118016 3000
rect 117688 2984 117740 2990
rect 117688 2926 117740 2932
rect 117228 2032 117280 2038
rect 117228 1974 117280 1980
rect 116492 1964 116544 1970
rect 116492 1906 116544 1912
rect 116400 1896 116452 1902
rect 116400 1838 116452 1844
rect 116308 1760 116360 1766
rect 116308 1702 116360 1708
rect 116216 1692 116268 1698
rect 116216 1634 116268 1640
rect 116124 1556 116176 1562
rect 116124 1498 116176 1504
rect 117700 1494 117728 2926
rect 115940 1488 115992 1494
rect 115940 1430 115992 1436
rect 117688 1488 117740 1494
rect 117688 1430 117740 1436
rect 117976 1426 118004 2994
rect 443656 2514 443992 2530
rect 294788 2508 294840 2514
rect 294788 2450 294840 2456
rect 425796 2508 425848 2514
rect 425796 2450 425848 2456
rect 443644 2508 443992 2514
rect 443696 2502 443992 2508
rect 443644 2450 443696 2456
rect 143644 2094 143980 2122
rect 193600 2094 193936 2122
rect 243648 2094 243984 2122
rect 293604 2094 293940 2122
rect 143644 1494 143672 2094
rect 143632 1488 143684 1494
rect 143632 1430 143684 1436
rect 163778 1456 163834 1465
rect 109776 1420 109828 1426
rect 109776 1362 109828 1368
rect 117964 1420 118016 1426
rect 193600 1426 193628 2094
rect 229282 1592 229338 1601
rect 229282 1527 229338 1536
rect 163778 1391 163834 1400
rect 193588 1420 193640 1426
rect 117964 1362 118016 1368
rect 163792 800 163820 1391
rect 193588 1362 193640 1368
rect 229296 800 229324 1527
rect 243648 1465 243676 2094
rect 293604 1601 293632 2094
rect 293590 1592 293646 1601
rect 293590 1527 293646 1536
rect 243634 1456 243690 1465
rect 294800 1426 294828 2450
rect 343652 2094 343988 2122
rect 393608 2094 393944 2122
rect 343652 1426 343680 2094
rect 393608 1465 393636 2094
rect 360290 1456 360346 1465
rect 243634 1391 243690 1400
rect 294788 1420 294840 1426
rect 294788 1362 294840 1368
rect 343640 1420 343692 1426
rect 360290 1391 360346 1400
rect 393594 1456 393650 1465
rect 393594 1391 393650 1400
rect 343640 1362 343692 1368
rect 294800 800 294828 1362
rect 360304 800 360332 1391
rect 425808 800 425836 2450
rect 520936 2281 520964 3295
rect 520922 2272 520978 2281
rect 520922 2207 520978 2216
rect 521106 2136 521162 2145
rect 493612 2094 493948 2122
rect 493612 1426 493640 2094
rect 521106 2071 521162 2080
rect 491300 1420 491352 1426
rect 491300 1362 491352 1368
rect 493600 1420 493652 1426
rect 493600 1362 493652 1368
rect 491312 800 491340 1362
rect 32770 -400 32826 800
rect 98274 -400 98330 800
rect 163778 -400 163834 800
rect 229282 -400 229338 800
rect 294786 -400 294842 800
rect 360290 -400 360346 800
rect 425794 -400 425850 800
rect 491298 -400 491354 800
rect 521120 785 521148 2071
rect 521106 776 521162 785
rect 521106 711 521162 720
<< via2 >>
rect 16302 159432 16358 159488
rect 16578 153720 16634 153776
rect 19890 153856 19946 153912
rect 23018 159296 23074 159352
rect 28078 156576 28134 156632
rect 29826 159568 29882 159624
rect 31482 156712 31538 156768
rect 33966 157936 34022 157992
rect 40682 158072 40738 158128
rect 44086 158208 44142 158264
rect 42430 156848 42486 156904
rect 27250 153992 27306 154048
rect 49146 156984 49202 157040
rect 57518 158344 57574 158400
rect 54298 154264 54354 154320
rect 51078 154128 51134 154184
rect 12438 152496 12494 152552
rect 8850 152360 8906 152416
rect 61750 155216 61806 155272
rect 65982 157120 66038 157176
rect 69294 155488 69350 155544
rect 68466 155352 68522 155408
rect 76010 155624 76066 155680
rect 85302 155760 85358 155816
rect 89718 154400 89774 154456
rect 92018 155896 92074 155952
rect 104622 158480 104678 158536
rect 113086 157256 113142 157312
rect 118606 153332 118662 153368
rect 118606 153312 118608 153332
rect 118608 153312 118660 153332
rect 118660 153312 118662 153332
rect 102598 149504 102654 149560
rect 109682 149504 109738 149560
rect 99286 149368 99342 149424
rect 105266 149368 105322 149424
rect 113822 143656 113878 143712
rect 116122 148688 116178 148744
rect 116122 147328 116178 147384
rect 116030 145696 116086 145752
rect 116214 143384 116270 143440
rect 116490 141752 116546 141808
rect 116398 139984 116454 140040
rect 116214 137808 116270 137864
rect 116398 136040 116454 136096
rect 116122 133728 116178 133784
rect 113914 132504 113970 132560
rect 116122 132232 116178 132288
rect 116122 130328 116178 130384
rect 116122 128016 116178 128072
rect 116122 126384 116178 126440
rect 116122 123800 116178 123856
rect 116122 122576 116178 122632
rect 114006 120808 114062 120864
rect 116122 120672 116178 120728
rect 116122 118360 116178 118416
rect 116122 116728 116178 116784
rect 116122 114144 116178 114200
rect 116122 112920 116178 112976
rect 116122 111152 116178 111208
rect 114098 109520 114154 109576
rect 116122 108840 116178 108896
rect 114190 98096 114246 98152
rect 119986 153332 120042 153368
rect 119986 153312 119988 153332
rect 119988 153312 120040 153332
rect 120040 153312 120042 153332
rect 127806 159432 127862 159488
rect 126242 152632 126298 152688
rect 126242 152360 126298 152416
rect 127806 153040 127862 153096
rect 128818 152496 128874 152552
rect 132038 153720 132094 153776
rect 131394 153040 131450 153096
rect 134614 153856 134670 153912
rect 137374 159452 137430 159488
rect 137374 159432 137376 159452
rect 137376 159432 137428 159452
rect 137428 159432 137430 159452
rect 136546 159296 136602 159352
rect 138570 159432 138626 159488
rect 139398 159568 139454 159624
rect 139858 159588 139914 159624
rect 139858 159568 139860 159588
rect 139860 159568 139912 159588
rect 139912 159568 139914 159588
rect 139950 156576 140006 156632
rect 139766 153992 139822 154048
rect 144918 159568 144974 159624
rect 142710 156712 142766 156768
rect 143630 152632 143686 152688
rect 144918 157936 144974 157992
rect 149610 158072 149666 158128
rect 150990 156848 151046 156904
rect 152554 158208 152610 158264
rect 157246 159588 157302 159624
rect 157246 159568 157248 159588
rect 157248 159568 157300 159588
rect 157300 159568 157302 159588
rect 157338 159432 157394 159488
rect 156418 156984 156474 157040
rect 158350 154128 158406 154184
rect 160926 154264 160982 154320
rect 162858 158344 162914 158400
rect 166078 155216 166134 155272
rect 169298 157120 169354 157176
rect 171138 155488 171194 155544
rect 171230 155352 171286 155408
rect 177026 155624 177082 155680
rect 184018 155760 184074 155816
rect 185214 154284 185270 154320
rect 185214 154264 185216 154284
rect 185216 154264 185268 154284
rect 185268 154264 185270 154284
rect 186226 154980 186228 155000
rect 186228 154980 186280 155000
rect 186280 154980 186282 155000
rect 186226 154944 186282 154980
rect 186594 154980 186596 155000
rect 186596 154980 186648 155000
rect 186648 154980 186650 155000
rect 186594 154944 186650 154980
rect 187238 154400 187294 154456
rect 188342 153448 188398 153504
rect 189170 155896 189226 155952
rect 191470 154264 191526 154320
rect 192390 153448 192446 153504
rect 198738 158480 198794 158536
rect 204718 159296 204774 159352
rect 203890 155352 203946 155408
rect 205270 157256 205326 157312
rect 209686 156612 209688 156632
rect 209688 156612 209740 156632
rect 209740 156612 209742 156632
rect 209686 156576 209742 156612
rect 210790 156612 210792 156632
rect 210792 156612 210844 156632
rect 210844 156612 210846 156632
rect 210790 156576 210846 156612
rect 209134 155352 209190 155408
rect 211526 153720 211582 153776
rect 227442 152360 227498 152416
rect 274546 159432 274602 159488
rect 275190 159296 275246 159352
rect 280986 153720 281042 153776
rect 283010 153856 283066 153912
rect 286230 153876 286286 153912
rect 286230 153856 286232 153876
rect 286232 153856 286284 153876
rect 286284 153856 286286 153876
rect 292578 152360 292634 152416
rect 313462 152360 313518 152416
rect 328550 159432 328606 159488
rect 357438 152360 357494 152416
rect 407670 152360 407726 152416
rect 427634 150184 427690 150240
rect 428048 150184 428104 150240
rect 431222 152496 431278 152552
rect 430578 152360 430634 152416
rect 444654 152632 444710 152688
rect 445574 152632 445630 152688
rect 448610 152496 448666 152552
rect 519726 163104 519782 163160
rect 519542 161608 519598 161664
rect 519358 158616 519414 158672
rect 519634 160112 519690 160168
rect 519542 148416 519598 148472
rect 520002 157120 520058 157176
rect 519818 151136 519874 151192
rect 519726 149776 519782 149832
rect 519726 148144 519782 148200
rect 519634 147056 519690 147112
rect 519358 145696 519414 145752
rect 519542 145152 519598 145208
rect 519266 140528 519322 140584
rect 519358 139032 519414 139088
rect 519266 129376 519322 129432
rect 519450 137400 519506 137456
rect 519358 128016 519414 128072
rect 519634 142160 519690 142216
rect 519542 133456 519598 133512
rect 519542 131552 519598 131608
rect 519450 126656 519506 126712
rect 519266 122440 519322 122496
rect 519910 149640 519966 149696
rect 519818 138896 519874 138952
rect 520094 155624 520150 155680
rect 520002 144336 520058 144392
rect 520186 154128 520242 154184
rect 520094 142976 520150 143032
rect 521106 152632 521162 152688
rect 521014 146648 521070 146704
rect 520922 143656 520978 143712
rect 520186 141616 520242 141672
rect 519910 137536 519966 137592
rect 519726 136176 519782 136232
rect 520186 136040 520242 136096
rect 520002 134544 520058 134600
rect 519634 130736 519690 130792
rect 519818 130056 519874 130112
rect 519634 128560 519690 128616
rect 519542 121216 519598 121272
rect 519358 121080 519414 121136
rect 519266 113056 519322 113112
rect 519450 119584 519506 119640
rect 519358 111696 519414 111752
rect 519726 127064 519782 127120
rect 519634 118496 519690 118552
rect 519910 125568 519966 125624
rect 519818 119856 519874 119912
rect 519818 118088 519874 118144
rect 519726 117136 519782 117192
rect 519726 113464 519782 113520
rect 519634 111968 519690 112024
rect 519542 110472 519598 110528
rect 519450 110336 519506 110392
rect 117226 107344 117282 107400
rect 117134 104488 117190 104544
rect 117042 103128 117098 103184
rect 520094 133048 520150 133104
rect 520002 123936 520058 123992
rect 521106 140256 521162 140312
rect 521014 134680 521070 134736
rect 520922 132096 520978 132152
rect 520186 125160 520242 125216
rect 520186 124072 520242 124128
rect 520094 122576 520150 122632
rect 520002 116456 520058 116512
rect 519910 115504 519966 115560
rect 519818 108976 519874 109032
rect 520094 114960 520150 115016
rect 520002 107480 520058 107536
rect 520186 114416 520242 114472
rect 520830 108976 520886 109032
rect 520094 105984 520150 106040
rect 520278 105984 520334 106040
rect 519726 104760 519782 104816
rect 519634 103400 519690 103456
rect 519542 102040 519598 102096
rect 116950 101496 117006 101552
rect 116858 99320 116914 99376
rect 520738 102992 520794 103048
rect 520278 97824 520334 97880
rect 116766 97688 116822 97744
rect 116674 95784 116730 95840
rect 520278 95512 520334 95568
rect 116582 93608 116638 93664
rect 519726 92248 519782 92304
rect 115938 91840 115994 91896
rect 116122 89528 116178 89584
rect 115938 88032 115994 88088
rect 114466 86980 114468 87000
rect 114468 86980 114520 87000
rect 114520 86980 114522 87000
rect 114466 86944 114522 86980
rect 116030 86128 116086 86184
rect 116582 83816 116638 83872
rect 116122 82320 116178 82376
rect 115938 80028 115994 80064
rect 115938 80008 115940 80028
rect 115940 80008 115992 80028
rect 115992 80008 115994 80028
rect 519634 86400 519690 86456
rect 519266 81912 519322 81968
rect 116674 78512 116730 78568
rect 520094 90888 520150 90944
rect 520002 89392 520058 89448
rect 519818 87896 519874 87952
rect 519726 85448 519782 85504
rect 519726 84904 519782 84960
rect 519634 80008 519690 80064
rect 520922 107480 520978 107536
rect 520830 100680 520886 100736
rect 521014 104488 521070 104544
rect 520922 99320 520978 99376
rect 521198 101496 521254 101552
rect 521014 96328 521070 96384
rect 520738 95104 520794 95160
rect 520922 93880 520978 93936
rect 520278 88168 520334 88224
rect 521474 100000 521530 100056
rect 521382 98504 521438 98560
rect 521198 93744 521254 93800
rect 521566 97008 521622 97064
rect 521474 92384 521530 92440
rect 521382 91024 521438 91080
rect 521566 89664 521622 89720
rect 520922 86808 520978 86864
rect 520094 84088 520150 84144
rect 520094 83408 520150 83464
rect 520002 82728 520058 82784
rect 519818 81368 519874 81424
rect 519910 78920 519966 78976
rect 519726 78240 519782 78296
rect 519818 77424 519874 77480
rect 519266 76472 519322 76528
rect 519726 75928 519782 75984
rect 116674 73480 116730 73536
rect 116030 71848 116086 71904
rect 45650 2644 45706 2680
rect 45650 2624 45652 2644
rect 45652 2624 45704 2644
rect 45704 2624 45706 2644
rect 49974 2644 50030 2680
rect 49974 2624 49976 2644
rect 49976 2624 50028 2644
rect 50028 2624 50030 2644
rect 19338 1808 19394 1864
rect 15934 1672 15990 1728
rect 12622 1536 12678 1592
rect 9310 1400 9366 1456
rect 66258 2624 66314 2680
rect 64878 2508 64934 2544
rect 64878 2488 64880 2508
rect 64880 2488 64932 2508
rect 64932 2488 64934 2508
rect 84566 2644 84622 2680
rect 84566 2624 84568 2644
rect 84568 2624 84620 2644
rect 84620 2624 84622 2644
rect 106094 2644 106150 2680
rect 106094 2624 106096 2644
rect 106096 2624 106148 2644
rect 106148 2624 106150 2644
rect 109590 2624 109646 2680
rect 67546 2352 67602 2408
rect 69018 2216 69074 2272
rect 76470 2216 76526 2272
rect 85854 2488 85910 2544
rect 85302 2352 85358 2408
rect 116214 69672 116270 69728
rect 115938 67768 115994 67824
rect 116582 66544 116638 66600
rect 520186 80416 520242 80472
rect 520094 76880 520150 76936
rect 520186 75112 520242 75168
rect 521198 74432 521254 74488
rect 519910 73752 519966 73808
rect 521014 72936 521070 72992
rect 519818 72392 519874 72448
rect 519726 71032 519782 71088
rect 520738 69808 520794 69864
rect 520462 66816 520518 66872
rect 520370 65320 520426 65376
rect 114466 64676 114468 64696
rect 114468 64676 114520 64696
rect 114520 64676 114522 64696
rect 114466 64640 114522 64676
rect 116030 63960 116086 64016
rect 116582 62192 116638 62248
rect 114190 53624 114246 53680
rect 116490 47232 116546 47288
rect 116214 44648 116270 44704
rect 114098 42336 114154 42392
rect 116122 41520 116178 41576
rect 114006 30912 114062 30968
rect 113914 19080 113970 19136
rect 113822 8200 113878 8256
rect 116306 42880 116362 42936
rect 115938 37324 115994 37360
rect 115938 37304 115940 37324
rect 115940 37304 115992 37324
rect 115992 37304 115994 37324
rect 116122 35128 116178 35184
rect 116122 33224 116178 33280
rect 116122 31864 116178 31920
rect 116122 29280 116178 29336
rect 116122 27668 116178 27704
rect 116122 27648 116124 27668
rect 116124 27648 116176 27668
rect 116176 27648 116178 27668
rect 116122 25472 116178 25528
rect 116122 23568 116178 23624
rect 116122 22344 116178 22400
rect 116214 19760 116270 19816
rect 116122 17992 116178 18048
rect 115938 13912 115994 13968
rect 115938 4528 115994 4584
rect 115846 2760 115902 2816
rect 116122 15816 116178 15872
rect 116398 38936 116454 38992
rect 521106 71440 521162 71496
rect 521014 68312 521070 68368
rect 521198 69672 521254 69728
rect 521198 68312 521254 68368
rect 521106 66952 521162 67008
rect 520738 65592 520794 65648
rect 521198 64232 521254 64288
rect 521198 63824 521254 63880
rect 520462 62872 520518 62928
rect 521014 62328 521070 62384
rect 520370 61512 520426 61568
rect 116674 60016 116730 60072
rect 520554 59336 520610 59392
rect 116766 58112 116822 58168
rect 519910 57840 519966 57896
rect 116858 56888 116914 56944
rect 519266 56344 519322 56400
rect 519082 54848 519138 54904
rect 116950 54304 117006 54360
rect 117042 52536 117098 52592
rect 521106 60832 521162 60888
rect 521014 58792 521070 58848
rect 521198 60152 521254 60208
rect 521106 57432 521162 57488
rect 520554 56072 520610 56128
rect 519910 54712 519966 54768
rect 519266 53352 519322 53408
rect 520002 53352 520058 53408
rect 519082 51992 519138 52048
rect 117134 51176 117190 51232
rect 520186 51856 520242 51912
rect 520002 50632 520058 50688
rect 520094 50360 520150 50416
rect 117226 48592 117282 48648
rect 520186 49272 520242 49328
rect 520186 48864 520242 48920
rect 520094 47776 520150 47832
rect 519910 47232 519966 47288
rect 519818 45736 519874 45792
rect 520186 46552 520242 46608
rect 519910 45192 519966 45248
rect 520186 44240 520242 44296
rect 519818 43832 519874 43888
rect 520738 42744 520794 42800
rect 520186 42472 520242 42528
rect 520738 41248 520794 41304
rect 520922 41248 520978 41304
rect 520922 39888 520978 39944
rect 520370 39752 520426 39808
rect 520370 38256 520426 38312
rect 520554 38256 520610 38312
rect 520554 37168 520610 37224
rect 521566 36760 521622 36816
rect 521566 35944 521622 36000
rect 520922 35264 520978 35320
rect 520922 34448 520978 34504
rect 521106 33768 521162 33824
rect 521106 33088 521162 33144
rect 521106 32272 521162 32328
rect 521106 31592 521162 31648
rect 521106 29280 521162 29336
rect 521106 28600 521162 28656
rect 521106 24792 521162 24848
rect 521106 23568 521162 23624
rect 520922 23160 520978 23216
rect 520922 22208 520978 22264
rect 520922 21664 520978 21720
rect 520922 20848 520978 20904
rect 521106 20168 521162 20224
rect 521106 19488 521162 19544
rect 520370 7384 520426 7440
rect 520370 6704 520426 6760
rect 521106 6024 521162 6080
rect 521106 5208 521162 5264
rect 521106 4664 521162 4720
rect 521106 3712 521162 3768
rect 520922 3304 520978 3360
rect 163778 1400 163834 1456
rect 229282 1536 229338 1592
rect 293590 1536 293646 1592
rect 243634 1400 243690 1456
rect 360290 1400 360346 1456
rect 393594 1400 393650 1456
rect 520922 2216 520978 2272
rect 521106 2080 521162 2136
rect 521106 720 521162 776
<< metal3 >>
rect 519721 163162 519787 163165
rect 523200 163162 524400 163192
rect 519721 163160 524400 163162
rect 519721 163104 519726 163160
rect 519782 163104 524400 163160
rect 519721 163102 524400 163104
rect 519721 163099 519787 163102
rect 523200 163072 524400 163102
rect 519537 161666 519603 161669
rect 523200 161666 524400 161696
rect 519537 161664 524400 161666
rect 519537 161608 519542 161664
rect 519598 161608 524400 161664
rect 519537 161606 524400 161608
rect 519537 161603 519603 161606
rect 523200 161576 524400 161606
rect 519629 160170 519695 160173
rect 523200 160170 524400 160200
rect 519629 160168 524400 160170
rect 519629 160112 519634 160168
rect 519690 160112 524400 160168
rect 519629 160110 524400 160112
rect 519629 160107 519695 160110
rect 523200 160080 524400 160110
rect 29821 159626 29887 159629
rect 139393 159626 139459 159629
rect 29821 159624 139459 159626
rect 29821 159568 29826 159624
rect 29882 159568 139398 159624
rect 139454 159568 139459 159624
rect 29821 159566 139459 159568
rect 29821 159563 29887 159566
rect 139393 159563 139459 159566
rect 139853 159626 139919 159629
rect 144913 159626 144979 159629
rect 139853 159624 144979 159626
rect 139853 159568 139858 159624
rect 139914 159568 144918 159624
rect 144974 159568 144979 159624
rect 139853 159566 144979 159568
rect 139853 159563 139919 159566
rect 144913 159563 144979 159566
rect 157241 159626 157307 159629
rect 157241 159624 157350 159626
rect 157241 159568 157246 159624
rect 157302 159568 157350 159624
rect 157241 159563 157350 159568
rect 157290 159493 157350 159563
rect 16297 159490 16363 159493
rect 127801 159490 127867 159493
rect 16297 159488 127867 159490
rect 16297 159432 16302 159488
rect 16358 159432 127806 159488
rect 127862 159432 127867 159488
rect 16297 159430 127867 159432
rect 16297 159427 16363 159430
rect 127801 159427 127867 159430
rect 137369 159490 137435 159493
rect 138565 159490 138631 159493
rect 137369 159488 138631 159490
rect 137369 159432 137374 159488
rect 137430 159432 138570 159488
rect 138626 159432 138631 159488
rect 137369 159430 138631 159432
rect 157290 159488 157399 159493
rect 157290 159432 157338 159488
rect 157394 159432 157399 159488
rect 157290 159430 157399 159432
rect 137369 159427 137435 159430
rect 138565 159427 138631 159430
rect 157333 159427 157399 159430
rect 274541 159490 274607 159493
rect 328545 159490 328611 159493
rect 274541 159488 328611 159490
rect 274541 159432 274546 159488
rect 274602 159432 328550 159488
rect 328606 159432 328611 159488
rect 274541 159430 328611 159432
rect 274541 159427 274607 159430
rect 328545 159427 328611 159430
rect 23013 159354 23079 159357
rect 136541 159354 136607 159357
rect 23013 159352 136607 159354
rect 23013 159296 23018 159352
rect 23074 159296 136546 159352
rect 136602 159296 136607 159352
rect 23013 159294 136607 159296
rect 23013 159291 23079 159294
rect 136541 159291 136607 159294
rect 204713 159354 204779 159357
rect 275185 159354 275251 159357
rect 204713 159352 275251 159354
rect 204713 159296 204718 159352
rect 204774 159296 275190 159352
rect 275246 159296 275251 159352
rect 204713 159294 275251 159296
rect 204713 159291 204779 159294
rect 275185 159291 275251 159294
rect 519353 158674 519419 158677
rect 523200 158674 524400 158704
rect 519353 158672 524400 158674
rect 519353 158616 519358 158672
rect 519414 158616 524400 158672
rect 519353 158614 524400 158616
rect 519353 158611 519419 158614
rect 523200 158584 524400 158614
rect 104617 158538 104683 158541
rect 198733 158538 198799 158541
rect 104617 158536 198799 158538
rect 104617 158480 104622 158536
rect 104678 158480 198738 158536
rect 198794 158480 198799 158536
rect 104617 158478 198799 158480
rect 104617 158475 104683 158478
rect 198733 158475 198799 158478
rect 57513 158402 57579 158405
rect 162853 158402 162919 158405
rect 57513 158400 162919 158402
rect 57513 158344 57518 158400
rect 57574 158344 162858 158400
rect 162914 158344 162919 158400
rect 57513 158342 162919 158344
rect 57513 158339 57579 158342
rect 162853 158339 162919 158342
rect 44081 158266 44147 158269
rect 152549 158266 152615 158269
rect 44081 158264 152615 158266
rect 44081 158208 44086 158264
rect 44142 158208 152554 158264
rect 152610 158208 152615 158264
rect 44081 158206 152615 158208
rect 44081 158203 44147 158206
rect 152549 158203 152615 158206
rect 40677 158130 40743 158133
rect 149605 158130 149671 158133
rect 40677 158128 149671 158130
rect 40677 158072 40682 158128
rect 40738 158072 149610 158128
rect 149666 158072 149671 158128
rect 40677 158070 149671 158072
rect 40677 158067 40743 158070
rect 149605 158067 149671 158070
rect 33961 157994 34027 157997
rect 144913 157994 144979 157997
rect 33961 157992 144979 157994
rect 33961 157936 33966 157992
rect 34022 157936 144918 157992
rect 144974 157936 144979 157992
rect 33961 157934 144979 157936
rect 33961 157931 34027 157934
rect 144913 157931 144979 157934
rect 113081 157314 113147 157317
rect 205265 157314 205331 157317
rect 113081 157312 205331 157314
rect 113081 157256 113086 157312
rect 113142 157256 205270 157312
rect 205326 157256 205331 157312
rect 113081 157254 205331 157256
rect 113081 157251 113147 157254
rect 205265 157251 205331 157254
rect 65977 157178 66043 157181
rect 169293 157178 169359 157181
rect 65977 157176 169359 157178
rect 65977 157120 65982 157176
rect 66038 157120 169298 157176
rect 169354 157120 169359 157176
rect 65977 157118 169359 157120
rect 65977 157115 66043 157118
rect 169293 157115 169359 157118
rect 519997 157178 520063 157181
rect 523200 157178 524400 157208
rect 519997 157176 524400 157178
rect 519997 157120 520002 157176
rect 520058 157120 524400 157176
rect 519997 157118 524400 157120
rect 519997 157115 520063 157118
rect 523200 157088 524400 157118
rect 49141 157042 49207 157045
rect 156413 157042 156479 157045
rect 49141 157040 156479 157042
rect 49141 156984 49146 157040
rect 49202 156984 156418 157040
rect 156474 156984 156479 157040
rect 49141 156982 156479 156984
rect 49141 156979 49207 156982
rect 156413 156979 156479 156982
rect 42425 156906 42491 156909
rect 150985 156906 151051 156909
rect 42425 156904 151051 156906
rect 42425 156848 42430 156904
rect 42486 156848 150990 156904
rect 151046 156848 151051 156904
rect 42425 156846 151051 156848
rect 42425 156843 42491 156846
rect 150985 156843 151051 156846
rect 31477 156770 31543 156773
rect 142705 156770 142771 156773
rect 31477 156768 142771 156770
rect 31477 156712 31482 156768
rect 31538 156712 142710 156768
rect 142766 156712 142771 156768
rect 31477 156710 142771 156712
rect 31477 156707 31543 156710
rect 142705 156707 142771 156710
rect 28073 156634 28139 156637
rect 139945 156634 140011 156637
rect 28073 156632 140011 156634
rect 28073 156576 28078 156632
rect 28134 156576 139950 156632
rect 140006 156576 140011 156632
rect 28073 156574 140011 156576
rect 28073 156571 28139 156574
rect 139945 156571 140011 156574
rect 209681 156634 209747 156637
rect 210785 156634 210851 156637
rect 209681 156632 210851 156634
rect 209681 156576 209686 156632
rect 209742 156576 210790 156632
rect 210846 156576 210851 156632
rect 209681 156574 210851 156576
rect 209681 156571 209747 156574
rect 210785 156571 210851 156574
rect 92013 155954 92079 155957
rect 189165 155954 189231 155957
rect 92013 155952 189231 155954
rect 92013 155896 92018 155952
rect 92074 155896 189170 155952
rect 189226 155896 189231 155952
rect 92013 155894 189231 155896
rect 92013 155891 92079 155894
rect 189165 155891 189231 155894
rect 85297 155818 85363 155821
rect 184013 155818 184079 155821
rect 85297 155816 184079 155818
rect 85297 155760 85302 155816
rect 85358 155760 184018 155816
rect 184074 155760 184079 155816
rect 85297 155758 184079 155760
rect 85297 155755 85363 155758
rect 184013 155755 184079 155758
rect 76005 155682 76071 155685
rect 177021 155682 177087 155685
rect 76005 155680 177087 155682
rect 76005 155624 76010 155680
rect 76066 155624 177026 155680
rect 177082 155624 177087 155680
rect 76005 155622 177087 155624
rect 76005 155619 76071 155622
rect 177021 155619 177087 155622
rect 520089 155682 520155 155685
rect 523200 155682 524400 155712
rect 520089 155680 524400 155682
rect 520089 155624 520094 155680
rect 520150 155624 524400 155680
rect 520089 155622 524400 155624
rect 520089 155619 520155 155622
rect 523200 155592 524400 155622
rect 69289 155546 69355 155549
rect 171133 155546 171199 155549
rect 69289 155544 171199 155546
rect 69289 155488 69294 155544
rect 69350 155488 171138 155544
rect 171194 155488 171199 155544
rect 69289 155486 171199 155488
rect 69289 155483 69355 155486
rect 171133 155483 171199 155486
rect 68461 155410 68527 155413
rect 171225 155410 171291 155413
rect 68461 155408 171291 155410
rect 68461 155352 68466 155408
rect 68522 155352 171230 155408
rect 171286 155352 171291 155408
rect 68461 155350 171291 155352
rect 68461 155347 68527 155350
rect 171225 155347 171291 155350
rect 203885 155410 203951 155413
rect 209129 155410 209195 155413
rect 203885 155408 209195 155410
rect 203885 155352 203890 155408
rect 203946 155352 209134 155408
rect 209190 155352 209195 155408
rect 203885 155350 209195 155352
rect 203885 155347 203951 155350
rect 209129 155347 209195 155350
rect 61745 155274 61811 155277
rect 166073 155274 166139 155277
rect 61745 155272 166139 155274
rect 61745 155216 61750 155272
rect 61806 155216 166078 155272
rect 166134 155216 166139 155272
rect 61745 155214 166139 155216
rect 61745 155211 61811 155214
rect 166073 155211 166139 155214
rect 186221 155002 186287 155005
rect 186589 155002 186655 155005
rect 186221 155000 186655 155002
rect 186221 154944 186226 155000
rect 186282 154944 186594 155000
rect 186650 154944 186655 155000
rect 186221 154942 186655 154944
rect 186221 154939 186287 154942
rect 186589 154939 186655 154942
rect 89713 154458 89779 154461
rect 187233 154458 187299 154461
rect 89713 154456 187299 154458
rect 89713 154400 89718 154456
rect 89774 154400 187238 154456
rect 187294 154400 187299 154456
rect 89713 154398 187299 154400
rect 89713 154395 89779 154398
rect 187233 154395 187299 154398
rect 54293 154322 54359 154325
rect 160921 154322 160987 154325
rect 54293 154320 160987 154322
rect 54293 154264 54298 154320
rect 54354 154264 160926 154320
rect 160982 154264 160987 154320
rect 54293 154262 160987 154264
rect 54293 154259 54359 154262
rect 160921 154259 160987 154262
rect 185209 154322 185275 154325
rect 191465 154322 191531 154325
rect 185209 154320 191531 154322
rect 185209 154264 185214 154320
rect 185270 154264 191470 154320
rect 191526 154264 191531 154320
rect 185209 154262 191531 154264
rect 185209 154259 185275 154262
rect 191465 154259 191531 154262
rect 51073 154186 51139 154189
rect 158345 154186 158411 154189
rect 51073 154184 158411 154186
rect 51073 154128 51078 154184
rect 51134 154128 158350 154184
rect 158406 154128 158411 154184
rect 51073 154126 158411 154128
rect 51073 154123 51139 154126
rect 158345 154123 158411 154126
rect 520181 154186 520247 154189
rect 523200 154186 524400 154216
rect 520181 154184 524400 154186
rect 520181 154128 520186 154184
rect 520242 154128 524400 154184
rect 520181 154126 524400 154128
rect 520181 154123 520247 154126
rect 523200 154096 524400 154126
rect 27245 154050 27311 154053
rect 139761 154050 139827 154053
rect 27245 154048 139827 154050
rect 27245 153992 27250 154048
rect 27306 153992 139766 154048
rect 139822 153992 139827 154048
rect 27245 153990 139827 153992
rect 27245 153987 27311 153990
rect 139761 153987 139827 153990
rect 19885 153914 19951 153917
rect 134609 153914 134675 153917
rect 19885 153912 134675 153914
rect 19885 153856 19890 153912
rect 19946 153856 134614 153912
rect 134670 153856 134675 153912
rect 19885 153854 134675 153856
rect 19885 153851 19951 153854
rect 134609 153851 134675 153854
rect 283005 153914 283071 153917
rect 286225 153914 286291 153917
rect 283005 153912 286291 153914
rect 283005 153856 283010 153912
rect 283066 153856 286230 153912
rect 286286 153856 286291 153912
rect 283005 153854 286291 153856
rect 283005 153851 283071 153854
rect 286225 153851 286291 153854
rect 16573 153778 16639 153781
rect 132033 153778 132099 153781
rect 16573 153776 132099 153778
rect 16573 153720 16578 153776
rect 16634 153720 132038 153776
rect 132094 153720 132099 153776
rect 16573 153718 132099 153720
rect 16573 153715 16639 153718
rect 132033 153715 132099 153718
rect 211521 153778 211587 153781
rect 280981 153778 281047 153781
rect 211521 153776 281047 153778
rect 211521 153720 211526 153776
rect 211582 153720 280986 153776
rect 281042 153720 281047 153776
rect 211521 153718 281047 153720
rect 211521 153715 211587 153718
rect 280981 153715 281047 153718
rect 188337 153506 188403 153509
rect 192385 153506 192451 153509
rect 188337 153504 192451 153506
rect 188337 153448 188342 153504
rect 188398 153448 192390 153504
rect 192446 153448 192451 153504
rect 188337 153446 192451 153448
rect 188337 153443 188403 153446
rect 192385 153443 192451 153446
rect 118601 153370 118667 153373
rect 119981 153370 120047 153373
rect 118601 153368 120047 153370
rect 118601 153312 118606 153368
rect 118662 153312 119986 153368
rect 120042 153312 120047 153368
rect 118601 153310 120047 153312
rect 118601 153307 118667 153310
rect 119981 153307 120047 153310
rect 127801 153098 127867 153101
rect 131389 153098 131455 153101
rect 127801 153096 131455 153098
rect 127801 153040 127806 153096
rect 127862 153040 131394 153096
rect 131450 153040 131455 153096
rect 127801 153038 131455 153040
rect 127801 153035 127867 153038
rect 131389 153035 131455 153038
rect 126237 152690 126303 152693
rect 143625 152690 143691 152693
rect 126237 152688 143691 152690
rect 126237 152632 126242 152688
rect 126298 152632 143630 152688
rect 143686 152632 143691 152688
rect 126237 152630 143691 152632
rect 126237 152627 126303 152630
rect 143625 152627 143691 152630
rect 444649 152690 444715 152693
rect 445569 152690 445635 152693
rect 444649 152688 445635 152690
rect 444649 152632 444654 152688
rect 444710 152632 445574 152688
rect 445630 152632 445635 152688
rect 444649 152630 445635 152632
rect 444649 152627 444715 152630
rect 445569 152627 445635 152630
rect 521101 152690 521167 152693
rect 523200 152690 524400 152720
rect 521101 152688 524400 152690
rect 521101 152632 521106 152688
rect 521162 152632 524400 152688
rect 521101 152630 524400 152632
rect 521101 152627 521167 152630
rect 523200 152600 524400 152630
rect 12433 152554 12499 152557
rect 128813 152554 128879 152557
rect 12433 152552 128879 152554
rect 12433 152496 12438 152552
rect 12494 152496 128818 152552
rect 128874 152496 128879 152552
rect 12433 152494 128879 152496
rect 12433 152491 12499 152494
rect 128813 152491 128879 152494
rect 431217 152554 431283 152557
rect 448605 152554 448671 152557
rect 431217 152552 448671 152554
rect 431217 152496 431222 152552
rect 431278 152496 448610 152552
rect 448666 152496 448671 152552
rect 431217 152494 448671 152496
rect 431217 152491 431283 152494
rect 448605 152491 448671 152494
rect 8845 152418 8911 152421
rect 126237 152418 126303 152421
rect 8845 152416 126303 152418
rect 8845 152360 8850 152416
rect 8906 152360 126242 152416
rect 126298 152360 126303 152416
rect 8845 152358 126303 152360
rect 8845 152355 8911 152358
rect 126237 152355 126303 152358
rect 227437 152418 227503 152421
rect 292573 152418 292639 152421
rect 227437 152416 292639 152418
rect 227437 152360 227442 152416
rect 227498 152360 292578 152416
rect 292634 152360 292639 152416
rect 227437 152358 292639 152360
rect 227437 152355 227503 152358
rect 292573 152355 292639 152358
rect 313457 152418 313523 152421
rect 357433 152418 357499 152421
rect 313457 152416 357499 152418
rect 313457 152360 313462 152416
rect 313518 152360 357438 152416
rect 357494 152360 357499 152416
rect 313457 152358 357499 152360
rect 313457 152355 313523 152358
rect 357433 152355 357499 152358
rect 407665 152418 407731 152421
rect 430573 152418 430639 152421
rect 407665 152416 430639 152418
rect 407665 152360 407670 152416
rect 407726 152360 430578 152416
rect 430634 152360 430639 152416
rect 407665 152358 430639 152360
rect 407665 152355 407731 152358
rect 430573 152355 430639 152358
rect 519813 151194 519879 151197
rect 523200 151194 524400 151224
rect 519813 151192 524400 151194
rect 519813 151136 519818 151192
rect 519874 151136 524400 151192
rect 519813 151134 524400 151136
rect 519813 151131 519879 151134
rect 523200 151104 524400 151134
rect 427629 150242 427695 150245
rect 428043 150242 428109 150245
rect 427629 150240 428109 150242
rect 427629 150184 427634 150240
rect 427690 150184 428048 150240
rect 428104 150184 428109 150240
rect 427629 150182 428109 150184
rect 427629 150179 427695 150182
rect 428043 150179 428109 150182
rect 519721 149834 519787 149837
rect 518758 149832 519787 149834
rect 518758 149776 519726 149832
rect 519782 149776 519787 149832
rect 518758 149774 519787 149776
rect 102593 149562 102659 149565
rect 109677 149562 109743 149565
rect 102593 149560 109743 149562
rect 102593 149504 102598 149560
rect 102654 149504 109682 149560
rect 109738 149504 109743 149560
rect 102593 149502 109743 149504
rect 102593 149499 102659 149502
rect 109677 149499 109743 149502
rect 99281 149426 99347 149429
rect 105261 149426 105327 149429
rect 99281 149424 105327 149426
rect 99281 149368 99286 149424
rect 99342 149368 105266 149424
rect 105322 149368 105327 149424
rect 99281 149366 105327 149368
rect 99281 149363 99347 149366
rect 105261 149363 105327 149366
rect 518758 149260 518818 149774
rect 519721 149771 519787 149774
rect 519905 149698 519971 149701
rect 523200 149698 524400 149728
rect 519905 149696 524400 149698
rect 519905 149640 519910 149696
rect 519966 149640 524400 149696
rect 519905 149638 524400 149640
rect 519905 149635 519971 149638
rect 523200 149608 524400 149638
rect 116117 148746 116183 148749
rect 119110 148746 119170 148988
rect 116117 148744 119170 148746
rect 116117 148688 116122 148744
rect 116178 148688 119170 148744
rect 116117 148686 119170 148688
rect 116117 148683 116183 148686
rect 519537 148474 519603 148477
rect 518758 148472 519603 148474
rect 518758 148416 519542 148472
rect 519598 148416 519603 148472
rect 518758 148414 519603 148416
rect 518758 147900 518818 148414
rect 519537 148411 519603 148414
rect 519721 148202 519787 148205
rect 523200 148202 524400 148232
rect 519721 148200 524400 148202
rect 519721 148144 519726 148200
rect 519782 148144 524400 148200
rect 519721 148142 524400 148144
rect 519721 148139 519787 148142
rect 523200 148112 524400 148142
rect 116117 147386 116183 147389
rect 116117 147384 119170 147386
rect 116117 147328 116122 147384
rect 116178 147328 119170 147384
rect 116117 147326 119170 147328
rect 116117 147323 116183 147326
rect 119110 147084 119170 147326
rect 519629 147114 519695 147117
rect 518758 147112 519695 147114
rect 518758 147056 519634 147112
rect 519690 147056 519695 147112
rect 518758 147054 519695 147056
rect 518758 146540 518818 147054
rect 519629 147051 519695 147054
rect 521009 146706 521075 146709
rect 523200 146706 524400 146736
rect 521009 146704 524400 146706
rect 521009 146648 521014 146704
rect 521070 146648 524400 146704
rect 521009 146646 524400 146648
rect 521009 146643 521075 146646
rect 523200 146616 524400 146646
rect 116025 145754 116091 145757
rect 519353 145754 519419 145757
rect 116025 145752 119170 145754
rect 116025 145696 116030 145752
rect 116086 145696 119170 145752
rect 116025 145694 119170 145696
rect 116025 145691 116091 145694
rect 119110 145180 119170 145694
rect 518758 145752 519419 145754
rect 518758 145696 519358 145752
rect 519414 145696 519419 145752
rect 518758 145694 519419 145696
rect 518758 145180 518818 145694
rect 519353 145691 519419 145694
rect 519537 145210 519603 145213
rect 523200 145210 524400 145240
rect 519537 145208 524400 145210
rect 519537 145152 519542 145208
rect 519598 145152 524400 145208
rect 519537 145150 524400 145152
rect 519537 145147 519603 145150
rect 523200 145120 524400 145150
rect 519997 144394 520063 144397
rect 518758 144392 520063 144394
rect 518758 144336 520002 144392
rect 520058 144336 520063 144392
rect 518758 144334 520063 144336
rect 110830 143714 110890 144228
rect 518758 143820 518818 144334
rect 519997 144331 520063 144334
rect 113817 143714 113883 143717
rect 110830 143712 113883 143714
rect 110830 143656 113822 143712
rect 113878 143656 113883 143712
rect 110830 143654 113883 143656
rect 113817 143651 113883 143654
rect 520917 143714 520983 143717
rect 523200 143714 524400 143744
rect 520917 143712 524400 143714
rect 520917 143656 520922 143712
rect 520978 143656 524400 143712
rect 520917 143654 524400 143656
rect 520917 143651 520983 143654
rect 523200 143624 524400 143654
rect 116209 143442 116275 143445
rect 116209 143440 119170 143442
rect 116209 143384 116214 143440
rect 116270 143384 119170 143440
rect 116209 143382 119170 143384
rect 116209 143379 116275 143382
rect 119110 143276 119170 143382
rect 520089 143034 520155 143037
rect 518758 143032 520155 143034
rect 518758 142976 520094 143032
rect 520150 142976 520155 143032
rect 518758 142974 520155 142976
rect 518758 142460 518818 142974
rect 520089 142971 520155 142974
rect 519629 142218 519695 142221
rect 523200 142218 524400 142248
rect 519629 142216 524400 142218
rect 519629 142160 519634 142216
rect 519690 142160 524400 142216
rect 519629 142158 524400 142160
rect 519629 142155 519695 142158
rect 523200 142128 524400 142158
rect 116485 141810 116551 141813
rect 116485 141808 119170 141810
rect 116485 141752 116490 141808
rect 116546 141752 119170 141808
rect 116485 141750 119170 141752
rect 116485 141747 116551 141750
rect 119110 141372 119170 141750
rect 520181 141674 520247 141677
rect 518758 141672 520247 141674
rect 518758 141616 520186 141672
rect 520242 141616 520247 141672
rect 518758 141614 520247 141616
rect 518758 141100 518818 141614
rect 520181 141611 520247 141614
rect 519261 140586 519327 140589
rect 523200 140586 524400 140616
rect 519261 140584 524400 140586
rect 519261 140528 519266 140584
rect 519322 140528 524400 140584
rect 519261 140526 524400 140528
rect 519261 140523 519327 140526
rect 523200 140496 524400 140526
rect 521101 140314 521167 140317
rect 518758 140312 521167 140314
rect 518758 140256 521106 140312
rect 521162 140256 521167 140312
rect 518758 140254 521167 140256
rect 116393 140042 116459 140045
rect 116393 140040 119170 140042
rect 116393 139984 116398 140040
rect 116454 139984 119170 140040
rect 116393 139982 119170 139984
rect 116393 139979 116459 139982
rect 119110 139468 119170 139982
rect 518758 139740 518818 140254
rect 521101 140251 521167 140254
rect 519353 139090 519419 139093
rect 523200 139090 524400 139120
rect 519353 139088 524400 139090
rect 519353 139032 519358 139088
rect 519414 139032 524400 139088
rect 519353 139030 524400 139032
rect 519353 139027 519419 139030
rect 523200 139000 524400 139030
rect 519813 138954 519879 138957
rect 518758 138952 519879 138954
rect 518758 138896 519818 138952
rect 519874 138896 519879 138952
rect 518758 138894 519879 138896
rect 518758 138380 518818 138894
rect 519813 138891 519879 138894
rect 116209 137866 116275 137869
rect 116209 137864 119170 137866
rect 116209 137808 116214 137864
rect 116270 137808 119170 137864
rect 116209 137806 119170 137808
rect 116209 137803 116275 137806
rect 119110 137564 119170 137806
rect 519905 137594 519971 137597
rect 523200 137594 524400 137624
rect 518758 137592 519971 137594
rect 518758 137536 519910 137592
rect 519966 137536 519971 137592
rect 518758 137534 519971 137536
rect 518758 137020 518818 137534
rect 519905 137531 519971 137534
rect 520046 137534 524400 137594
rect 519445 137458 519511 137461
rect 520046 137458 520106 137534
rect 523200 137504 524400 137534
rect 519445 137456 520106 137458
rect 519445 137400 519450 137456
rect 519506 137400 520106 137456
rect 519445 137398 520106 137400
rect 519445 137395 519511 137398
rect 519721 136234 519787 136237
rect 518758 136232 519787 136234
rect 518758 136176 519726 136232
rect 519782 136176 519787 136232
rect 518758 136174 519787 136176
rect 116393 136098 116459 136101
rect 116393 136096 119170 136098
rect 116393 136040 116398 136096
rect 116454 136040 119170 136096
rect 116393 136038 119170 136040
rect 116393 136035 116459 136038
rect 119110 135524 119170 136038
rect 518758 135660 518818 136174
rect 519721 136171 519787 136174
rect 520181 136098 520247 136101
rect 523200 136098 524400 136128
rect 520181 136096 524400 136098
rect 520181 136040 520186 136096
rect 520242 136040 524400 136096
rect 520181 136038 524400 136040
rect 520181 136035 520247 136038
rect 523200 136008 524400 136038
rect 521009 134738 521075 134741
rect 518758 134736 521075 134738
rect 518758 134680 521014 134736
rect 521070 134680 521075 134736
rect 518758 134678 521075 134680
rect 518758 134300 518818 134678
rect 521009 134675 521075 134678
rect 519997 134602 520063 134605
rect 523200 134602 524400 134632
rect 519997 134600 524400 134602
rect 519997 134544 520002 134600
rect 520058 134544 524400 134600
rect 519997 134542 524400 134544
rect 519997 134539 520063 134542
rect 523200 134512 524400 134542
rect 116117 133786 116183 133789
rect 116117 133784 119170 133786
rect 116117 133728 116122 133784
rect 116178 133728 119170 133784
rect 116117 133726 119170 133728
rect 116117 133723 116183 133726
rect 119110 133620 119170 133726
rect 519537 133514 519603 133517
rect 518758 133512 519603 133514
rect 518758 133456 519542 133512
rect 519598 133456 519603 133512
rect 518758 133454 519603 133456
rect 518758 132940 518818 133454
rect 519537 133451 519603 133454
rect 520089 133106 520155 133109
rect 523200 133106 524400 133136
rect 520089 133104 524400 133106
rect 520089 133048 520094 133104
rect 520150 133048 524400 133104
rect 520089 133046 524400 133048
rect 520089 133043 520155 133046
rect 523200 133016 524400 133046
rect 110830 132562 110890 132804
rect 113909 132562 113975 132565
rect 110830 132560 113975 132562
rect 110830 132504 113914 132560
rect 113970 132504 113975 132560
rect 110830 132502 113975 132504
rect 113909 132499 113975 132502
rect 116117 132290 116183 132293
rect 116117 132288 119170 132290
rect 116117 132232 116122 132288
rect 116178 132232 119170 132288
rect 116117 132230 119170 132232
rect 116117 132227 116183 132230
rect 119110 131716 119170 132230
rect 520917 132154 520983 132157
rect 518758 132152 520983 132154
rect 518758 132096 520922 132152
rect 520978 132096 520983 132152
rect 518758 132094 520983 132096
rect 518758 131580 518818 132094
rect 520917 132091 520983 132094
rect 519537 131610 519603 131613
rect 523200 131610 524400 131640
rect 519537 131608 524400 131610
rect 519537 131552 519542 131608
rect 519598 131552 524400 131608
rect 519537 131550 524400 131552
rect 519537 131547 519603 131550
rect 523200 131520 524400 131550
rect 519629 130794 519695 130797
rect 518758 130792 519695 130794
rect 518758 130736 519634 130792
rect 519690 130736 519695 130792
rect 518758 130734 519695 130736
rect 116117 130386 116183 130389
rect 116117 130384 119170 130386
rect 116117 130328 116122 130384
rect 116178 130328 119170 130384
rect 116117 130326 119170 130328
rect 116117 130323 116183 130326
rect 119110 129812 119170 130326
rect 518758 130220 518818 130734
rect 519629 130731 519695 130734
rect 519813 130114 519879 130117
rect 523200 130114 524400 130144
rect 519813 130112 524400 130114
rect 519813 130056 519818 130112
rect 519874 130056 524400 130112
rect 519813 130054 524400 130056
rect 519813 130051 519879 130054
rect 523200 130024 524400 130054
rect 519261 129434 519327 129437
rect 518758 129432 519327 129434
rect 518758 129376 519266 129432
rect 519322 129376 519327 129432
rect 518758 129374 519327 129376
rect 518758 128860 518818 129374
rect 519261 129371 519327 129374
rect 519629 128618 519695 128621
rect 523200 128618 524400 128648
rect 519629 128616 524400 128618
rect 519629 128560 519634 128616
rect 519690 128560 524400 128616
rect 519629 128558 524400 128560
rect 519629 128555 519695 128558
rect 523200 128528 524400 128558
rect 116117 128074 116183 128077
rect 519353 128074 519419 128077
rect 116117 128072 119170 128074
rect 116117 128016 116122 128072
rect 116178 128016 119170 128072
rect 116117 128014 119170 128016
rect 116117 128011 116183 128014
rect 119110 127908 119170 128014
rect 518758 128072 519419 128074
rect 518758 128016 519358 128072
rect 519414 128016 519419 128072
rect 518758 128014 519419 128016
rect 518758 127500 518818 128014
rect 519353 128011 519419 128014
rect 519721 127122 519787 127125
rect 523200 127122 524400 127152
rect 519721 127120 524400 127122
rect 519721 127064 519726 127120
rect 519782 127064 524400 127120
rect 519721 127062 524400 127064
rect 519721 127059 519787 127062
rect 523200 127032 524400 127062
rect 519445 126714 519511 126717
rect 518758 126712 519511 126714
rect 518758 126656 519450 126712
rect 519506 126656 519511 126712
rect 518758 126654 519511 126656
rect 116117 126442 116183 126445
rect 116117 126440 119170 126442
rect 116117 126384 116122 126440
rect 116178 126384 119170 126440
rect 116117 126382 119170 126384
rect 116117 126379 116183 126382
rect 119110 126004 119170 126382
rect 518758 126140 518818 126654
rect 519445 126651 519511 126654
rect 519905 125626 519971 125629
rect 523200 125626 524400 125656
rect 519905 125624 524400 125626
rect 519905 125568 519910 125624
rect 519966 125568 524400 125624
rect 519905 125566 524400 125568
rect 519905 125563 519971 125566
rect 523200 125536 524400 125566
rect 520181 125218 520247 125221
rect 518758 125216 520247 125218
rect 518758 125160 520186 125216
rect 520242 125160 520247 125216
rect 518758 125158 520247 125160
rect 518758 124780 518818 125158
rect 520181 125155 520247 125158
rect 520181 124130 520247 124133
rect 523200 124130 524400 124160
rect 520181 124128 524400 124130
rect 116117 123858 116183 123861
rect 119110 123858 119170 124100
rect 520181 124072 520186 124128
rect 520242 124072 524400 124128
rect 520181 124070 524400 124072
rect 520181 124067 520247 124070
rect 523200 124040 524400 124070
rect 519997 123994 520063 123997
rect 116117 123856 119170 123858
rect 116117 123800 116122 123856
rect 116178 123800 119170 123856
rect 116117 123798 119170 123800
rect 518758 123992 520063 123994
rect 518758 123936 520002 123992
rect 520058 123936 520063 123992
rect 518758 123934 520063 123936
rect 116117 123795 116183 123798
rect 518758 123420 518818 123934
rect 519997 123931 520063 123934
rect 116117 122634 116183 122637
rect 520089 122634 520155 122637
rect 523200 122634 524400 122664
rect 116117 122632 119170 122634
rect 116117 122576 116122 122632
rect 116178 122576 119170 122632
rect 116117 122574 119170 122576
rect 116117 122571 116183 122574
rect 119110 122196 119170 122574
rect 518758 122632 520155 122634
rect 518758 122576 520094 122632
rect 520150 122576 520155 122632
rect 518758 122574 520155 122576
rect 518758 122060 518818 122574
rect 520089 122571 520155 122574
rect 520230 122574 524400 122634
rect 519261 122498 519327 122501
rect 520230 122498 520290 122574
rect 523200 122544 524400 122574
rect 519261 122496 520290 122498
rect 519261 122440 519266 122496
rect 519322 122440 520290 122496
rect 519261 122438 520290 122440
rect 519261 122435 519327 122438
rect 110830 120866 110890 121380
rect 519537 121274 519603 121277
rect 518758 121272 519603 121274
rect 518758 121216 519542 121272
rect 519598 121216 519603 121272
rect 518758 121214 519603 121216
rect 114001 120866 114067 120869
rect 110830 120864 114067 120866
rect 110830 120808 114006 120864
rect 114062 120808 114067 120864
rect 110830 120806 114067 120808
rect 114001 120803 114067 120806
rect 116117 120730 116183 120733
rect 116117 120728 119170 120730
rect 116117 120672 116122 120728
rect 116178 120672 119170 120728
rect 518758 120700 518818 121214
rect 519537 121211 519603 121214
rect 519353 121138 519419 121141
rect 523200 121138 524400 121168
rect 519353 121136 524400 121138
rect 519353 121080 519358 121136
rect 519414 121080 524400 121136
rect 519353 121078 524400 121080
rect 519353 121075 519419 121078
rect 523200 121048 524400 121078
rect 116117 120670 119170 120672
rect 116117 120667 116183 120670
rect 119110 120156 119170 120670
rect 519813 119914 519879 119917
rect 518758 119912 519879 119914
rect 518758 119856 519818 119912
rect 519874 119856 519879 119912
rect 518758 119854 519879 119856
rect 518758 119340 518818 119854
rect 519813 119851 519879 119854
rect 519445 119642 519511 119645
rect 523200 119642 524400 119672
rect 519445 119640 524400 119642
rect 519445 119584 519450 119640
rect 519506 119584 524400 119640
rect 519445 119582 524400 119584
rect 519445 119579 519511 119582
rect 523200 119552 524400 119582
rect 519629 118554 519695 118557
rect 518758 118552 519695 118554
rect 518758 118496 519634 118552
rect 519690 118496 519695 118552
rect 518758 118494 519695 118496
rect 116117 118418 116183 118421
rect 116117 118416 119170 118418
rect 116117 118360 116122 118416
rect 116178 118360 119170 118416
rect 116117 118358 119170 118360
rect 116117 118355 116183 118358
rect 119110 118252 119170 118358
rect 518758 117980 518818 118494
rect 519629 118491 519695 118494
rect 519813 118146 519879 118149
rect 523200 118146 524400 118176
rect 519813 118144 524400 118146
rect 519813 118088 519818 118144
rect 519874 118088 524400 118144
rect 519813 118086 524400 118088
rect 519813 118083 519879 118086
rect 523200 118056 524400 118086
rect 519721 117194 519787 117197
rect 518758 117192 519787 117194
rect 518758 117136 519726 117192
rect 519782 117136 519787 117192
rect 518758 117134 519787 117136
rect 116117 116786 116183 116789
rect 116117 116784 119170 116786
rect 116117 116728 116122 116784
rect 116178 116728 119170 116784
rect 116117 116726 119170 116728
rect 116117 116723 116183 116726
rect 119110 116348 119170 116726
rect 518758 116620 518818 117134
rect 519721 117131 519787 117134
rect 519997 116514 520063 116517
rect 523200 116514 524400 116544
rect 519997 116512 524400 116514
rect 519997 116456 520002 116512
rect 520058 116456 524400 116512
rect 519997 116454 524400 116456
rect 519997 116451 520063 116454
rect 523200 116424 524400 116454
rect 519905 115562 519971 115565
rect 518758 115560 519971 115562
rect 518758 115504 519910 115560
rect 519966 115504 519971 115560
rect 518758 115502 519971 115504
rect 518758 115260 518818 115502
rect 519905 115499 519971 115502
rect 520089 115018 520155 115021
rect 523200 115018 524400 115048
rect 520089 115016 524400 115018
rect 520089 114960 520094 115016
rect 520150 114960 524400 115016
rect 520089 114958 524400 114960
rect 520089 114955 520155 114958
rect 523200 114928 524400 114958
rect 520181 114474 520247 114477
rect 518758 114472 520247 114474
rect 116117 114202 116183 114205
rect 119110 114202 119170 114444
rect 116117 114200 119170 114202
rect 116117 114144 116122 114200
rect 116178 114144 119170 114200
rect 116117 114142 119170 114144
rect 518758 114416 520186 114472
rect 520242 114416 520247 114472
rect 518758 114414 520247 114416
rect 116117 114139 116183 114142
rect 518758 113900 518818 114414
rect 520181 114411 520247 114414
rect 519721 113522 519787 113525
rect 523200 113522 524400 113552
rect 519721 113520 524400 113522
rect 519721 113464 519726 113520
rect 519782 113464 524400 113520
rect 519721 113462 524400 113464
rect 519721 113459 519787 113462
rect 523200 113432 524400 113462
rect 519261 113114 519327 113117
rect 518758 113112 519327 113114
rect 518758 113056 519266 113112
rect 519322 113056 519327 113112
rect 518758 113054 519327 113056
rect 116117 112978 116183 112981
rect 116117 112976 119170 112978
rect 116117 112920 116122 112976
rect 116178 112920 119170 112976
rect 116117 112918 119170 112920
rect 116117 112915 116183 112918
rect 119110 112540 119170 112918
rect 518758 112540 518818 113054
rect 519261 113051 519327 113054
rect 519629 112026 519695 112029
rect 523200 112026 524400 112056
rect 519629 112024 524400 112026
rect 519629 111968 519634 112024
rect 519690 111968 524400 112024
rect 519629 111966 524400 111968
rect 519629 111963 519695 111966
rect 523200 111936 524400 111966
rect 519353 111754 519419 111757
rect 518758 111752 519419 111754
rect 518758 111696 519358 111752
rect 519414 111696 519419 111752
rect 518758 111694 519419 111696
rect 116117 111210 116183 111213
rect 116117 111208 119170 111210
rect 116117 111152 116122 111208
rect 116178 111152 119170 111208
rect 518758 111180 518818 111694
rect 519353 111691 519419 111694
rect 116117 111150 119170 111152
rect 116117 111147 116183 111150
rect 119110 110636 119170 111150
rect 519537 110530 519603 110533
rect 523200 110530 524400 110560
rect 519537 110528 524400 110530
rect 519537 110472 519542 110528
rect 519598 110472 524400 110528
rect 519537 110470 524400 110472
rect 519537 110467 519603 110470
rect 523200 110440 524400 110470
rect 519445 110394 519511 110397
rect 518758 110392 519511 110394
rect 518758 110336 519450 110392
rect 519506 110336 519511 110392
rect 518758 110334 519511 110336
rect 110830 109578 110890 110092
rect 518758 109820 518818 110334
rect 519445 110331 519511 110334
rect 114093 109578 114159 109581
rect 110830 109576 114159 109578
rect 110830 109520 114098 109576
rect 114154 109520 114159 109576
rect 110830 109518 114159 109520
rect 114093 109515 114159 109518
rect 519813 109034 519879 109037
rect 518758 109032 519879 109034
rect 518758 108976 519818 109032
rect 519874 108976 519879 109032
rect 518758 108974 519879 108976
rect 116117 108898 116183 108901
rect 116117 108896 119170 108898
rect 116117 108840 116122 108896
rect 116178 108840 119170 108896
rect 116117 108838 119170 108840
rect 116117 108835 116183 108838
rect 119110 108732 119170 108838
rect 518758 108460 518818 108974
rect 519813 108971 519879 108974
rect 520825 109034 520891 109037
rect 523200 109034 524400 109064
rect 520825 109032 524400 109034
rect 520825 108976 520830 109032
rect 520886 108976 524400 109032
rect 520825 108974 524400 108976
rect 520825 108971 520891 108974
rect 523200 108944 524400 108974
rect 519997 107538 520063 107541
rect 518758 107536 520063 107538
rect 518758 107480 520002 107536
rect 520058 107480 520063 107536
rect 518758 107478 520063 107480
rect 117221 107402 117287 107405
rect 117221 107400 119170 107402
rect 117221 107344 117226 107400
rect 117282 107344 119170 107400
rect 117221 107342 119170 107344
rect 117221 107339 117287 107342
rect 119110 106828 119170 107342
rect 518758 107100 518818 107478
rect 519997 107475 520063 107478
rect 520917 107538 520983 107541
rect 523200 107538 524400 107568
rect 520917 107536 524400 107538
rect 520917 107480 520922 107536
rect 520978 107480 524400 107536
rect 520917 107478 524400 107480
rect 520917 107475 520983 107478
rect 523200 107448 524400 107478
rect 520089 106042 520155 106045
rect 518758 106040 520155 106042
rect 518758 105984 520094 106040
rect 520150 105984 520155 106040
rect 518758 105982 520155 105984
rect 518758 105740 518818 105982
rect 520089 105979 520155 105982
rect 520273 106042 520339 106045
rect 523200 106042 524400 106072
rect 520273 106040 524400 106042
rect 520273 105984 520278 106040
rect 520334 105984 524400 106040
rect 520273 105982 524400 105984
rect 520273 105979 520339 105982
rect 523200 105952 524400 105982
rect 519721 104818 519787 104821
rect 518758 104816 519787 104818
rect 117129 104546 117195 104549
rect 119110 104546 119170 104788
rect 117129 104544 119170 104546
rect 117129 104488 117134 104544
rect 117190 104488 119170 104544
rect 117129 104486 119170 104488
rect 518758 104760 519726 104816
rect 519782 104760 519787 104816
rect 518758 104758 519787 104760
rect 117129 104483 117195 104486
rect 518758 104380 518818 104758
rect 519721 104755 519787 104758
rect 521009 104546 521075 104549
rect 523200 104546 524400 104576
rect 521009 104544 524400 104546
rect 521009 104488 521014 104544
rect 521070 104488 524400 104544
rect 521009 104486 524400 104488
rect 521009 104483 521075 104486
rect 523200 104456 524400 104486
rect 519629 103458 519695 103461
rect 518758 103456 519695 103458
rect 518758 103400 519634 103456
rect 519690 103400 519695 103456
rect 518758 103398 519695 103400
rect 117037 103186 117103 103189
rect 117037 103184 119170 103186
rect 117037 103128 117042 103184
rect 117098 103128 119170 103184
rect 117037 103126 119170 103128
rect 117037 103123 117103 103126
rect 119110 102884 119170 103126
rect 518758 103020 518818 103398
rect 519629 103395 519695 103398
rect 520733 103050 520799 103053
rect 523200 103050 524400 103080
rect 520733 103048 524400 103050
rect 520733 102992 520738 103048
rect 520794 102992 524400 103048
rect 520733 102990 524400 102992
rect 520733 102987 520799 102990
rect 523200 102960 524400 102990
rect 519537 102098 519603 102101
rect 518758 102096 519603 102098
rect 518758 102040 519542 102096
rect 519598 102040 519603 102096
rect 518758 102038 519603 102040
rect 518758 101660 518818 102038
rect 519537 102035 519603 102038
rect 116945 101554 117011 101557
rect 521193 101554 521259 101557
rect 523200 101554 524400 101584
rect 116945 101552 119170 101554
rect 116945 101496 116950 101552
rect 117006 101496 119170 101552
rect 116945 101494 119170 101496
rect 116945 101491 117011 101494
rect 119110 100980 119170 101494
rect 521193 101552 524400 101554
rect 521193 101496 521198 101552
rect 521254 101496 524400 101552
rect 521193 101494 524400 101496
rect 521193 101491 521259 101494
rect 523200 101464 524400 101494
rect 520825 100738 520891 100741
rect 518758 100736 520891 100738
rect 518758 100680 520830 100736
rect 520886 100680 520891 100736
rect 518758 100678 520891 100680
rect 518758 100300 518818 100678
rect 520825 100675 520891 100678
rect 521469 100058 521535 100061
rect 523200 100058 524400 100088
rect 521469 100056 524400 100058
rect 521469 100000 521474 100056
rect 521530 100000 524400 100056
rect 521469 99998 524400 100000
rect 521469 99995 521535 99998
rect 523200 99968 524400 99998
rect 116853 99378 116919 99381
rect 520917 99378 520983 99381
rect 116853 99376 119170 99378
rect 116853 99320 116858 99376
rect 116914 99320 119170 99376
rect 116853 99318 119170 99320
rect 116853 99315 116919 99318
rect 119110 99076 119170 99318
rect 518758 99376 520983 99378
rect 518758 99320 520922 99376
rect 520978 99320 520983 99376
rect 518758 99318 520983 99320
rect 518758 98940 518818 99318
rect 520917 99315 520983 99318
rect 110830 98154 110890 98668
rect 521377 98562 521443 98565
rect 523200 98562 524400 98592
rect 521377 98560 524400 98562
rect 521377 98504 521382 98560
rect 521438 98504 524400 98560
rect 521377 98502 524400 98504
rect 521377 98499 521443 98502
rect 523200 98472 524400 98502
rect 114185 98154 114251 98157
rect 110830 98152 114251 98154
rect 110830 98096 114190 98152
rect 114246 98096 114251 98152
rect 110830 98094 114251 98096
rect 114185 98091 114251 98094
rect 520273 97882 520339 97885
rect 518758 97880 520339 97882
rect 518758 97824 520278 97880
rect 520334 97824 520339 97880
rect 518758 97822 520339 97824
rect 116761 97746 116827 97749
rect 116761 97744 119170 97746
rect 116761 97688 116766 97744
rect 116822 97688 119170 97744
rect 116761 97686 119170 97688
rect 116761 97683 116827 97686
rect 119110 97172 119170 97686
rect 518758 97580 518818 97822
rect 520273 97819 520339 97822
rect 521561 97066 521627 97069
rect 523200 97066 524400 97096
rect 521561 97064 524400 97066
rect 521561 97008 521566 97064
rect 521622 97008 524400 97064
rect 521561 97006 524400 97008
rect 521561 97003 521627 97006
rect 523200 96976 524400 97006
rect 521009 96386 521075 96389
rect 518758 96384 521075 96386
rect 518758 96328 521014 96384
rect 521070 96328 521075 96384
rect 518758 96326 521075 96328
rect 518758 96220 518818 96326
rect 521009 96323 521075 96326
rect 116669 95842 116735 95845
rect 116669 95840 119170 95842
rect 116669 95784 116674 95840
rect 116730 95784 119170 95840
rect 116669 95782 119170 95784
rect 116669 95779 116735 95782
rect 119110 95268 119170 95782
rect 520273 95570 520339 95573
rect 523200 95570 524400 95600
rect 520273 95568 524400 95570
rect 520273 95512 520278 95568
rect 520334 95512 524400 95568
rect 520273 95510 524400 95512
rect 520273 95507 520339 95510
rect 523200 95480 524400 95510
rect 520733 95162 520799 95165
rect 518758 95160 520799 95162
rect 518758 95104 520738 95160
rect 520794 95104 520799 95160
rect 518758 95102 520799 95104
rect 518758 94860 518818 95102
rect 520733 95099 520799 95102
rect 520917 93938 520983 93941
rect 523200 93938 524400 93968
rect 520917 93936 524400 93938
rect 520917 93880 520922 93936
rect 520978 93880 524400 93936
rect 520917 93878 524400 93880
rect 520917 93875 520983 93878
rect 523200 93848 524400 93878
rect 521193 93802 521259 93805
rect 518758 93800 521259 93802
rect 518758 93744 521198 93800
rect 521254 93744 521259 93800
rect 518758 93742 521259 93744
rect 116577 93666 116643 93669
rect 116577 93664 119170 93666
rect 116577 93608 116582 93664
rect 116638 93608 119170 93664
rect 116577 93606 119170 93608
rect 116577 93603 116643 93606
rect 119110 93364 119170 93606
rect 518758 93500 518818 93742
rect 521193 93739 521259 93742
rect 521469 92442 521535 92445
rect 523200 92442 524400 92472
rect 518758 92440 521535 92442
rect 518758 92384 521474 92440
rect 521530 92384 521535 92440
rect 518758 92382 521535 92384
rect 518758 92140 518818 92382
rect 521469 92379 521535 92382
rect 521702 92382 524400 92442
rect 519721 92306 519787 92309
rect 521702 92306 521762 92382
rect 523200 92352 524400 92382
rect 519721 92304 521762 92306
rect 519721 92248 519726 92304
rect 519782 92248 521762 92304
rect 519721 92246 521762 92248
rect 519721 92243 519787 92246
rect 115933 91898 115999 91901
rect 115933 91896 119170 91898
rect 115933 91840 115938 91896
rect 115994 91840 119170 91896
rect 115933 91838 119170 91840
rect 115933 91835 115999 91838
rect 119110 91324 119170 91838
rect 521377 91082 521443 91085
rect 518758 91080 521443 91082
rect 518758 91024 521382 91080
rect 521438 91024 521443 91080
rect 518758 91022 521443 91024
rect 518758 90780 518818 91022
rect 521377 91019 521443 91022
rect 520089 90946 520155 90949
rect 523200 90946 524400 90976
rect 520089 90944 524400 90946
rect 520089 90888 520094 90944
rect 520150 90888 524400 90944
rect 520089 90886 524400 90888
rect 520089 90883 520155 90886
rect 523200 90856 524400 90886
rect 521561 89722 521627 89725
rect 518758 89720 521627 89722
rect 518758 89664 521566 89720
rect 521622 89664 521627 89720
rect 518758 89662 521627 89664
rect 116117 89586 116183 89589
rect 116117 89584 119170 89586
rect 116117 89528 116122 89584
rect 116178 89528 119170 89584
rect 116117 89526 119170 89528
rect 116117 89523 116183 89526
rect 119110 89420 119170 89526
rect 518758 89420 518818 89662
rect 521561 89659 521627 89662
rect 519997 89450 520063 89453
rect 523200 89450 524400 89480
rect 519997 89448 524400 89450
rect 519997 89392 520002 89448
rect 520058 89392 524400 89448
rect 519997 89390 524400 89392
rect 519997 89387 520063 89390
rect 523200 89360 524400 89390
rect 520273 88226 520339 88229
rect 518758 88224 520339 88226
rect 518758 88168 520278 88224
rect 520334 88168 520339 88224
rect 518758 88166 520339 88168
rect 115933 88090 115999 88093
rect 115933 88088 119170 88090
rect 115933 88032 115938 88088
rect 115994 88032 119170 88088
rect 518758 88060 518818 88166
rect 520273 88163 520339 88166
rect 115933 88030 119170 88032
rect 115933 88027 115999 88030
rect 119110 87516 119170 88030
rect 519813 87954 519879 87957
rect 523200 87954 524400 87984
rect 519813 87952 524400 87954
rect 519813 87896 519818 87952
rect 519874 87896 524400 87952
rect 519813 87894 524400 87896
rect 519813 87891 519879 87894
rect 523200 87864 524400 87894
rect 110830 87002 110890 87244
rect 114461 87002 114527 87005
rect 110830 87000 114527 87002
rect 110830 86944 114466 87000
rect 114522 86944 114527 87000
rect 110830 86942 114527 86944
rect 114461 86939 114527 86942
rect 520917 86866 520983 86869
rect 518758 86864 520983 86866
rect 518758 86808 520922 86864
rect 520978 86808 520983 86864
rect 518758 86806 520983 86808
rect 518758 86700 518818 86806
rect 520917 86803 520983 86806
rect 519629 86458 519695 86461
rect 523200 86458 524400 86488
rect 519629 86456 524400 86458
rect 519629 86400 519634 86456
rect 519690 86400 524400 86456
rect 519629 86398 524400 86400
rect 519629 86395 519695 86398
rect 523200 86368 524400 86398
rect 116025 86186 116091 86189
rect 116025 86184 119170 86186
rect 116025 86128 116030 86184
rect 116086 86128 119170 86184
rect 116025 86126 119170 86128
rect 116025 86123 116091 86126
rect 119110 85612 119170 86126
rect 519721 85506 519787 85509
rect 518758 85504 519787 85506
rect 518758 85448 519726 85504
rect 519782 85448 519787 85504
rect 518758 85446 519787 85448
rect 518758 85340 518818 85446
rect 519721 85443 519787 85446
rect 519721 84962 519787 84965
rect 523200 84962 524400 84992
rect 519721 84960 524400 84962
rect 519721 84904 519726 84960
rect 519782 84904 524400 84960
rect 519721 84902 524400 84904
rect 519721 84899 519787 84902
rect 523200 84872 524400 84902
rect 520089 84146 520155 84149
rect 518758 84144 520155 84146
rect 518758 84088 520094 84144
rect 520150 84088 520155 84144
rect 518758 84086 520155 84088
rect 518758 83980 518818 84086
rect 520089 84083 520155 84086
rect 116577 83874 116643 83877
rect 116577 83872 119170 83874
rect 116577 83816 116582 83872
rect 116638 83816 119170 83872
rect 116577 83814 119170 83816
rect 116577 83811 116643 83814
rect 119110 83708 119170 83814
rect 520089 83466 520155 83469
rect 523200 83466 524400 83496
rect 520089 83464 524400 83466
rect 520089 83408 520094 83464
rect 520150 83408 524400 83464
rect 520089 83406 524400 83408
rect 520089 83403 520155 83406
rect 523200 83376 524400 83406
rect 519997 82786 520063 82789
rect 518758 82784 520063 82786
rect 518758 82728 520002 82784
rect 520058 82728 520063 82784
rect 518758 82726 520063 82728
rect 518758 82620 518818 82726
rect 519997 82723 520063 82726
rect 116117 82378 116183 82381
rect 116117 82376 119170 82378
rect 116117 82320 116122 82376
rect 116178 82320 119170 82376
rect 116117 82318 119170 82320
rect 116117 82315 116183 82318
rect 119110 81804 119170 82318
rect 519261 81970 519327 81973
rect 523200 81970 524400 82000
rect 519261 81968 524400 81970
rect 519261 81912 519266 81968
rect 519322 81912 524400 81968
rect 519261 81910 524400 81912
rect 519261 81907 519327 81910
rect 523200 81880 524400 81910
rect 519813 81426 519879 81429
rect 518758 81424 519879 81426
rect 518758 81368 519818 81424
rect 519874 81368 519879 81424
rect 518758 81366 519879 81368
rect 518758 81260 518818 81366
rect 519813 81363 519879 81366
rect 520181 80474 520247 80477
rect 523200 80474 524400 80504
rect 520181 80472 524400 80474
rect 520181 80416 520186 80472
rect 520242 80416 524400 80472
rect 520181 80414 524400 80416
rect 520181 80411 520247 80414
rect 523200 80384 524400 80414
rect 115933 80066 115999 80069
rect 519629 80066 519695 80069
rect 115933 80064 119170 80066
rect 115933 80008 115938 80064
rect 115994 80008 119170 80064
rect 115933 80006 119170 80008
rect 115933 80003 115999 80006
rect 119110 79900 119170 80006
rect 518758 80064 519695 80066
rect 518758 80008 519634 80064
rect 519690 80008 519695 80064
rect 518758 80006 519695 80008
rect 518758 79900 518818 80006
rect 519629 80003 519695 80006
rect 519905 78978 519971 78981
rect 523200 78978 524400 79008
rect 519905 78976 524400 78978
rect 519905 78920 519910 78976
rect 519966 78920 524400 78976
rect 519905 78918 524400 78920
rect 519905 78915 519971 78918
rect 523200 78888 524400 78918
rect 116669 78570 116735 78573
rect 116669 78568 119170 78570
rect 116669 78512 116674 78568
rect 116730 78512 119170 78568
rect 116669 78510 119170 78512
rect 116669 78507 116735 78510
rect 119110 77996 119170 78510
rect 518758 78298 518818 78540
rect 519721 78298 519787 78301
rect 518758 78296 519787 78298
rect 518758 78240 519726 78296
rect 519782 78240 519787 78296
rect 518758 78238 519787 78240
rect 519721 78235 519787 78238
rect 519813 77482 519879 77485
rect 523200 77482 524400 77512
rect 519813 77480 524400 77482
rect 519813 77424 519818 77480
rect 519874 77424 524400 77480
rect 519813 77422 524400 77424
rect 519813 77419 519879 77422
rect 523200 77392 524400 77422
rect 518758 76938 518818 77180
rect 520089 76938 520155 76941
rect 518758 76936 520155 76938
rect 518758 76880 520094 76936
rect 520150 76880 520155 76936
rect 518758 76878 520155 76880
rect 520089 76875 520155 76878
rect 519261 76530 519327 76533
rect 518758 76528 519327 76530
rect 518758 76472 519266 76528
rect 519322 76472 519327 76528
rect 518758 76470 519327 76472
rect 110830 76198 119170 76258
rect 110830 75956 110890 76198
rect 119110 75956 119170 76198
rect 518758 75956 518818 76470
rect 519261 76467 519327 76470
rect 519721 75986 519787 75989
rect 523200 75986 524400 76016
rect 519721 75984 524400 75986
rect 519721 75928 519726 75984
rect 519782 75928 524400 75984
rect 519721 75926 524400 75928
rect 519721 75923 519787 75926
rect 523200 75896 524400 75926
rect 520181 75170 520247 75173
rect 518758 75168 520247 75170
rect 518758 75112 520186 75168
rect 520242 75112 520247 75168
rect 518758 75110 520247 75112
rect 518758 74596 518818 75110
rect 520181 75107 520247 75110
rect 521193 74490 521259 74493
rect 523200 74490 524400 74520
rect 521193 74488 524400 74490
rect 521193 74432 521198 74488
rect 521254 74432 524400 74488
rect 521193 74430 524400 74432
rect 521193 74427 521259 74430
rect 523200 74400 524400 74430
rect 116669 73538 116735 73541
rect 119110 73538 119170 74052
rect 519905 73810 519971 73813
rect 116669 73536 119170 73538
rect 116669 73480 116674 73536
rect 116730 73480 119170 73536
rect 116669 73478 119170 73480
rect 518758 73808 519971 73810
rect 518758 73752 519910 73808
rect 519966 73752 519971 73808
rect 518758 73750 519971 73752
rect 116669 73475 116735 73478
rect 518758 73236 518818 73750
rect 519905 73747 519971 73750
rect 521009 72994 521075 72997
rect 523200 72994 524400 73024
rect 521009 72992 524400 72994
rect 521009 72936 521014 72992
rect 521070 72936 524400 72992
rect 521009 72934 524400 72936
rect 521009 72931 521075 72934
rect 523200 72904 524400 72934
rect 519813 72450 519879 72453
rect 518758 72448 519879 72450
rect 518758 72392 519818 72448
rect 519874 72392 519879 72448
rect 518758 72390 519879 72392
rect 116025 71906 116091 71909
rect 119110 71906 119170 72148
rect 116025 71904 119170 71906
rect 116025 71848 116030 71904
rect 116086 71848 119170 71904
rect 518758 71876 518818 72390
rect 519813 72387 519879 72390
rect 116025 71846 119170 71848
rect 116025 71843 116091 71846
rect 521101 71498 521167 71501
rect 523200 71498 524400 71528
rect 521101 71496 524400 71498
rect 521101 71440 521106 71496
rect 521162 71440 524400 71496
rect 521101 71438 524400 71440
rect 521101 71435 521167 71438
rect 523200 71408 524400 71438
rect 519721 71090 519787 71093
rect 518758 71088 519787 71090
rect 518758 71032 519726 71088
rect 519782 71032 519787 71088
rect 518758 71030 519787 71032
rect 518758 70516 518818 71030
rect 519721 71027 519787 71030
rect 116209 69730 116275 69733
rect 119110 69730 119170 70244
rect 520733 69866 520799 69869
rect 523200 69866 524400 69896
rect 520733 69864 524400 69866
rect 520733 69808 520738 69864
rect 520794 69808 524400 69864
rect 520733 69806 524400 69808
rect 520733 69803 520799 69806
rect 523200 69776 524400 69806
rect 521193 69730 521259 69733
rect 116209 69728 119170 69730
rect 116209 69672 116214 69728
rect 116270 69672 119170 69728
rect 116209 69670 119170 69672
rect 518758 69728 521259 69730
rect 518758 69672 521198 69728
rect 521254 69672 521259 69728
rect 518758 69670 521259 69672
rect 116209 69667 116275 69670
rect 518758 69156 518818 69670
rect 521193 69667 521259 69670
rect 521009 68370 521075 68373
rect 518758 68368 521075 68370
rect 115933 67826 115999 67829
rect 119110 67826 119170 68340
rect 115933 67824 119170 67826
rect 115933 67768 115938 67824
rect 115994 67768 119170 67824
rect 518758 68312 521014 68368
rect 521070 68312 521075 68368
rect 518758 68310 521075 68312
rect 518758 67796 518818 68310
rect 521009 68307 521075 68310
rect 521193 68370 521259 68373
rect 523200 68370 524400 68400
rect 521193 68368 524400 68370
rect 521193 68312 521198 68368
rect 521254 68312 524400 68368
rect 521193 68310 524400 68312
rect 521193 68307 521259 68310
rect 523200 68280 524400 68310
rect 115933 67766 119170 67768
rect 115933 67763 115999 67766
rect 521101 67010 521167 67013
rect 518758 67008 521167 67010
rect 518758 66952 521106 67008
rect 521162 66952 521167 67008
rect 518758 66950 521167 66952
rect 116577 66602 116643 66605
rect 116577 66600 119170 66602
rect 116577 66544 116582 66600
rect 116638 66544 119170 66600
rect 116577 66542 119170 66544
rect 116577 66539 116643 66542
rect 119110 66436 119170 66542
rect 518758 66436 518818 66950
rect 521101 66947 521167 66950
rect 520457 66874 520523 66877
rect 523200 66874 524400 66904
rect 520457 66872 524400 66874
rect 520457 66816 520462 66872
rect 520518 66816 524400 66872
rect 520457 66814 524400 66816
rect 520457 66811 520523 66814
rect 523200 66784 524400 66814
rect 520733 65650 520799 65653
rect 518758 65648 520799 65650
rect 518758 65592 520738 65648
rect 520794 65592 520799 65648
rect 518758 65590 520799 65592
rect 518758 65076 518818 65590
rect 520733 65587 520799 65590
rect 520365 65378 520431 65381
rect 523200 65378 524400 65408
rect 520365 65376 524400 65378
rect 520365 65320 520370 65376
rect 520426 65320 524400 65376
rect 520365 65318 524400 65320
rect 520365 65315 520431 65318
rect 523200 65288 524400 65318
rect 114461 64698 114527 64701
rect 110830 64696 114527 64698
rect 110830 64640 114466 64696
rect 114522 64640 114527 64696
rect 110830 64638 114527 64640
rect 110830 64532 110890 64638
rect 114461 64635 114527 64638
rect 116025 64018 116091 64021
rect 119110 64018 119170 64532
rect 521193 64290 521259 64293
rect 116025 64016 119170 64018
rect 116025 63960 116030 64016
rect 116086 63960 119170 64016
rect 116025 63958 119170 63960
rect 518758 64288 521259 64290
rect 518758 64232 521198 64288
rect 521254 64232 521259 64288
rect 518758 64230 521259 64232
rect 116025 63955 116091 63958
rect 518758 63716 518818 64230
rect 521193 64227 521259 64230
rect 521193 63882 521259 63885
rect 523200 63882 524400 63912
rect 521193 63880 524400 63882
rect 521193 63824 521198 63880
rect 521254 63824 524400 63880
rect 521193 63822 524400 63824
rect 521193 63819 521259 63822
rect 523200 63792 524400 63822
rect 520457 62930 520523 62933
rect 518758 62928 520523 62930
rect 518758 62872 520462 62928
rect 520518 62872 520523 62928
rect 518758 62870 520523 62872
rect 116577 62250 116643 62253
rect 119110 62250 119170 62628
rect 518758 62356 518818 62870
rect 520457 62867 520523 62870
rect 521009 62386 521075 62389
rect 523200 62386 524400 62416
rect 521009 62384 524400 62386
rect 521009 62328 521014 62384
rect 521070 62328 524400 62384
rect 521009 62326 524400 62328
rect 521009 62323 521075 62326
rect 523200 62296 524400 62326
rect 116577 62248 119170 62250
rect 116577 62192 116582 62248
rect 116638 62192 119170 62248
rect 116577 62190 119170 62192
rect 116577 62187 116643 62190
rect 520365 61570 520431 61573
rect 518758 61568 520431 61570
rect 518758 61512 520370 61568
rect 520426 61512 520431 61568
rect 518758 61510 520431 61512
rect 518758 60996 518818 61510
rect 520365 61507 520431 61510
rect 521101 60890 521167 60893
rect 523200 60890 524400 60920
rect 521101 60888 524400 60890
rect 521101 60832 521106 60888
rect 521162 60832 524400 60888
rect 521101 60830 524400 60832
rect 521101 60827 521167 60830
rect 523200 60800 524400 60830
rect 116669 60074 116735 60077
rect 119110 60074 119170 60588
rect 521193 60210 521259 60213
rect 116669 60072 119170 60074
rect 116669 60016 116674 60072
rect 116730 60016 119170 60072
rect 116669 60014 119170 60016
rect 518758 60208 521259 60210
rect 518758 60152 521198 60208
rect 521254 60152 521259 60208
rect 518758 60150 521259 60152
rect 116669 60011 116735 60014
rect 518758 59636 518818 60150
rect 521193 60147 521259 60150
rect 520549 59394 520615 59397
rect 523200 59394 524400 59424
rect 520549 59392 524400 59394
rect 520549 59336 520554 59392
rect 520610 59336 524400 59392
rect 520549 59334 524400 59336
rect 520549 59331 520615 59334
rect 523200 59304 524400 59334
rect 521009 58850 521075 58853
rect 518758 58848 521075 58850
rect 518758 58792 521014 58848
rect 521070 58792 521075 58848
rect 518758 58790 521075 58792
rect 116761 58170 116827 58173
rect 119110 58170 119170 58684
rect 518758 58276 518818 58790
rect 521009 58787 521075 58790
rect 116761 58168 119170 58170
rect 116761 58112 116766 58168
rect 116822 58112 119170 58168
rect 116761 58110 119170 58112
rect 116761 58107 116827 58110
rect 519905 57898 519971 57901
rect 523200 57898 524400 57928
rect 519905 57896 524400 57898
rect 519905 57840 519910 57896
rect 519966 57840 524400 57896
rect 519905 57838 524400 57840
rect 519905 57835 519971 57838
rect 523200 57808 524400 57838
rect 521101 57490 521167 57493
rect 518758 57488 521167 57490
rect 518758 57432 521106 57488
rect 521162 57432 521167 57488
rect 518758 57430 521167 57432
rect 116853 56946 116919 56949
rect 116853 56944 119170 56946
rect 116853 56888 116858 56944
rect 116914 56888 119170 56944
rect 518758 56916 518818 57430
rect 521101 57427 521167 57430
rect 116853 56886 119170 56888
rect 116853 56883 116919 56886
rect 119110 56780 119170 56886
rect 519261 56402 519327 56405
rect 523200 56402 524400 56432
rect 519261 56400 524400 56402
rect 519261 56344 519266 56400
rect 519322 56344 524400 56400
rect 519261 56342 524400 56344
rect 519261 56339 519327 56342
rect 523200 56312 524400 56342
rect 520549 56130 520615 56133
rect 518758 56128 520615 56130
rect 518758 56072 520554 56128
rect 520610 56072 520615 56128
rect 518758 56070 520615 56072
rect 518758 55556 518818 56070
rect 520549 56067 520615 56070
rect 519077 54906 519143 54909
rect 523200 54906 524400 54936
rect 519077 54904 524400 54906
rect 116945 54362 117011 54365
rect 119110 54362 119170 54876
rect 519077 54848 519082 54904
rect 519138 54848 524400 54904
rect 519077 54846 524400 54848
rect 519077 54843 519143 54846
rect 523200 54816 524400 54846
rect 519905 54770 519971 54773
rect 116945 54360 119170 54362
rect 116945 54304 116950 54360
rect 117006 54304 119170 54360
rect 116945 54302 119170 54304
rect 518758 54768 519971 54770
rect 518758 54712 519910 54768
rect 519966 54712 519971 54768
rect 518758 54710 519971 54712
rect 116945 54299 117011 54302
rect 518758 54196 518818 54710
rect 519905 54707 519971 54710
rect 114185 53682 114251 53685
rect 110830 53680 114251 53682
rect 110830 53624 114190 53680
rect 114246 53624 114251 53680
rect 110830 53622 114251 53624
rect 110830 53108 110890 53622
rect 114185 53619 114251 53622
rect 519261 53410 519327 53413
rect 518758 53408 519327 53410
rect 518758 53352 519266 53408
rect 519322 53352 519327 53408
rect 518758 53350 519327 53352
rect 117037 52594 117103 52597
rect 119110 52594 119170 52972
rect 518758 52836 518818 53350
rect 519261 53347 519327 53350
rect 519997 53410 520063 53413
rect 523200 53410 524400 53440
rect 519997 53408 524400 53410
rect 519997 53352 520002 53408
rect 520058 53352 524400 53408
rect 519997 53350 524400 53352
rect 519997 53347 520063 53350
rect 523200 53320 524400 53350
rect 117037 52592 119170 52594
rect 117037 52536 117042 52592
rect 117098 52536 119170 52592
rect 117037 52534 119170 52536
rect 117037 52531 117103 52534
rect 519077 52050 519143 52053
rect 518758 52048 519143 52050
rect 518758 51992 519082 52048
rect 519138 51992 519143 52048
rect 518758 51990 519143 51992
rect 518758 51476 518818 51990
rect 519077 51987 519143 51990
rect 520181 51914 520247 51917
rect 523200 51914 524400 51944
rect 520181 51912 524400 51914
rect 520181 51856 520186 51912
rect 520242 51856 524400 51912
rect 520181 51854 524400 51856
rect 520181 51851 520247 51854
rect 523200 51824 524400 51854
rect 117129 51234 117195 51237
rect 117129 51232 119170 51234
rect 117129 51176 117134 51232
rect 117190 51176 119170 51232
rect 117129 51174 119170 51176
rect 117129 51171 117195 51174
rect 119110 51068 119170 51174
rect 519997 50690 520063 50693
rect 518758 50688 520063 50690
rect 518758 50632 520002 50688
rect 520058 50632 520063 50688
rect 518758 50630 520063 50632
rect 518758 50116 518818 50630
rect 519997 50627 520063 50630
rect 520089 50418 520155 50421
rect 523200 50418 524400 50448
rect 520089 50416 524400 50418
rect 520089 50360 520094 50416
rect 520150 50360 524400 50416
rect 520089 50358 524400 50360
rect 520089 50355 520155 50358
rect 523200 50328 524400 50358
rect 520181 49330 520247 49333
rect 518758 49328 520247 49330
rect 518758 49272 520186 49328
rect 520242 49272 520247 49328
rect 518758 49270 520247 49272
rect 117221 48650 117287 48653
rect 119110 48650 119170 49164
rect 518758 48756 518818 49270
rect 520181 49267 520247 49270
rect 520181 48922 520247 48925
rect 523200 48922 524400 48952
rect 520181 48920 524400 48922
rect 520181 48864 520186 48920
rect 520242 48864 524400 48920
rect 520181 48862 524400 48864
rect 520181 48859 520247 48862
rect 523200 48832 524400 48862
rect 117221 48648 119170 48650
rect 117221 48592 117226 48648
rect 117282 48592 119170 48648
rect 117221 48590 119170 48592
rect 117221 48587 117287 48590
rect 520089 47834 520155 47837
rect 518758 47832 520155 47834
rect 518758 47776 520094 47832
rect 520150 47776 520155 47832
rect 518758 47774 520155 47776
rect 518758 47396 518818 47774
rect 520089 47771 520155 47774
rect 116485 47290 116551 47293
rect 519905 47290 519971 47293
rect 523200 47290 524400 47320
rect 116485 47288 119170 47290
rect 116485 47232 116490 47288
rect 116546 47232 119170 47288
rect 116485 47230 119170 47232
rect 116485 47227 116551 47230
rect 119110 47124 119170 47230
rect 519905 47288 524400 47290
rect 519905 47232 519910 47288
rect 519966 47232 524400 47288
rect 519905 47230 524400 47232
rect 519905 47227 519971 47230
rect 523200 47200 524400 47230
rect 520181 46610 520247 46613
rect 518758 46608 520247 46610
rect 518758 46552 520186 46608
rect 520242 46552 520247 46608
rect 518758 46550 520247 46552
rect 518758 46036 518818 46550
rect 520181 46547 520247 46550
rect 519813 45794 519879 45797
rect 523200 45794 524400 45824
rect 519813 45792 524400 45794
rect 519813 45736 519818 45792
rect 519874 45736 524400 45792
rect 519813 45734 524400 45736
rect 519813 45731 519879 45734
rect 523200 45704 524400 45734
rect 519905 45250 519971 45253
rect 518758 45248 519971 45250
rect 116209 44706 116275 44709
rect 119110 44706 119170 45220
rect 116209 44704 119170 44706
rect 116209 44648 116214 44704
rect 116270 44648 119170 44704
rect 518758 45192 519910 45248
rect 519966 45192 519971 45248
rect 518758 45190 519971 45192
rect 518758 44676 518818 45190
rect 519905 45187 519971 45190
rect 116209 44646 119170 44648
rect 116209 44643 116275 44646
rect 520181 44298 520247 44301
rect 523200 44298 524400 44328
rect 520181 44296 524400 44298
rect 520181 44240 520186 44296
rect 520242 44240 524400 44296
rect 520181 44238 524400 44240
rect 520181 44235 520247 44238
rect 523200 44208 524400 44238
rect 519813 43890 519879 43893
rect 518758 43888 519879 43890
rect 518758 43832 519818 43888
rect 519874 43832 519879 43888
rect 518758 43830 519879 43832
rect 518758 43316 518818 43830
rect 519813 43827 519879 43830
rect 116301 42938 116367 42941
rect 119110 42938 119170 43316
rect 116301 42936 119170 42938
rect 116301 42880 116306 42936
rect 116362 42880 119170 42936
rect 116301 42878 119170 42880
rect 116301 42875 116367 42878
rect 520733 42802 520799 42805
rect 523200 42802 524400 42832
rect 520733 42800 524400 42802
rect 520733 42744 520738 42800
rect 520794 42744 524400 42800
rect 520733 42742 524400 42744
rect 520733 42739 520799 42742
rect 523200 42712 524400 42742
rect 520181 42530 520247 42533
rect 518758 42528 520247 42530
rect 518758 42472 520186 42528
rect 520242 42472 520247 42528
rect 518758 42470 520247 42472
rect 114093 42394 114159 42397
rect 110830 42392 114159 42394
rect 110830 42336 114098 42392
rect 114154 42336 114159 42392
rect 110830 42334 114159 42336
rect 110830 41820 110890 42334
rect 114093 42331 114159 42334
rect 518758 41956 518818 42470
rect 520181 42467 520247 42470
rect 116117 41578 116183 41581
rect 116117 41576 119170 41578
rect 116117 41520 116122 41576
rect 116178 41520 119170 41576
rect 116117 41518 119170 41520
rect 116117 41515 116183 41518
rect 119110 41412 119170 41518
rect 520733 41306 520799 41309
rect 518758 41304 520799 41306
rect 518758 41248 520738 41304
rect 520794 41248 520799 41304
rect 518758 41246 520799 41248
rect 518758 40596 518818 41246
rect 520733 41243 520799 41246
rect 520917 41306 520983 41309
rect 523200 41306 524400 41336
rect 520917 41304 524400 41306
rect 520917 41248 520922 41304
rect 520978 41248 524400 41304
rect 520917 41246 524400 41248
rect 520917 41243 520983 41246
rect 523200 41216 524400 41246
rect 520917 39946 520983 39949
rect 518758 39944 520983 39946
rect 518758 39888 520922 39944
rect 520978 39888 520983 39944
rect 518758 39886 520983 39888
rect 116393 38994 116459 38997
rect 119110 38994 119170 39508
rect 518758 39236 518818 39886
rect 520917 39883 520983 39886
rect 520365 39810 520431 39813
rect 523200 39810 524400 39840
rect 520365 39808 524400 39810
rect 520365 39752 520370 39808
rect 520426 39752 524400 39808
rect 520365 39750 524400 39752
rect 520365 39747 520431 39750
rect 523200 39720 524400 39750
rect 116393 38992 119170 38994
rect 116393 38936 116398 38992
rect 116454 38936 119170 38992
rect 116393 38934 119170 38936
rect 116393 38931 116459 38934
rect 520365 38314 520431 38317
rect 518758 38312 520431 38314
rect 518758 38256 520370 38312
rect 520426 38256 520431 38312
rect 518758 38254 520431 38256
rect 518758 37876 518818 38254
rect 520365 38251 520431 38254
rect 520549 38314 520615 38317
rect 523200 38314 524400 38344
rect 520549 38312 524400 38314
rect 520549 38256 520554 38312
rect 520610 38256 524400 38312
rect 520549 38254 524400 38256
rect 520549 38251 520615 38254
rect 523200 38224 524400 38254
rect 115933 37362 115999 37365
rect 119110 37362 119170 37604
rect 115933 37360 119170 37362
rect 115933 37304 115938 37360
rect 115994 37304 119170 37360
rect 115933 37302 119170 37304
rect 115933 37299 115999 37302
rect 520549 37226 520615 37229
rect 518758 37224 520615 37226
rect 518758 37168 520554 37224
rect 520610 37168 520615 37224
rect 518758 37166 520615 37168
rect 518758 36516 518818 37166
rect 520549 37163 520615 37166
rect 521561 36818 521627 36821
rect 523200 36818 524400 36848
rect 521561 36816 524400 36818
rect 521561 36760 521566 36816
rect 521622 36760 524400 36816
rect 521561 36758 524400 36760
rect 521561 36755 521627 36758
rect 523200 36728 524400 36758
rect 521561 36002 521627 36005
rect 521561 36000 521670 36002
rect 521561 35944 521566 36000
rect 521622 35944 521670 36000
rect 521561 35939 521670 35944
rect 521610 35866 521670 35939
rect 518758 35806 521670 35866
rect 116117 35186 116183 35189
rect 119110 35186 119170 35700
rect 116117 35184 119170 35186
rect 116117 35128 116122 35184
rect 116178 35128 119170 35184
rect 518758 35156 518818 35806
rect 520917 35322 520983 35325
rect 523200 35322 524400 35352
rect 520917 35320 524400 35322
rect 520917 35264 520922 35320
rect 520978 35264 524400 35320
rect 520917 35262 524400 35264
rect 520917 35259 520983 35262
rect 523200 35232 524400 35262
rect 116117 35126 119170 35128
rect 116117 35123 116183 35126
rect 520917 34506 520983 34509
rect 518758 34504 520983 34506
rect 518758 34448 520922 34504
rect 520978 34448 520983 34504
rect 518758 34446 520983 34448
rect 518758 33796 518818 34446
rect 520917 34443 520983 34446
rect 521101 33826 521167 33829
rect 523200 33826 524400 33856
rect 521101 33824 524400 33826
rect 116117 33282 116183 33285
rect 119110 33282 119170 33796
rect 521101 33768 521106 33824
rect 521162 33768 524400 33824
rect 521101 33766 524400 33768
rect 521101 33763 521167 33766
rect 523200 33736 524400 33766
rect 116117 33280 119170 33282
rect 116117 33224 116122 33280
rect 116178 33224 119170 33280
rect 116117 33222 119170 33224
rect 116117 33219 116183 33222
rect 521101 33146 521167 33149
rect 518758 33144 521167 33146
rect 518758 33088 521106 33144
rect 521162 33088 521167 33144
rect 518758 33086 521167 33088
rect 518758 32436 518818 33086
rect 521101 33083 521167 33086
rect 521101 32330 521167 32333
rect 523200 32330 524400 32360
rect 521101 32328 524400 32330
rect 521101 32272 521106 32328
rect 521162 32272 524400 32328
rect 521101 32270 524400 32272
rect 521101 32267 521167 32270
rect 523200 32240 524400 32270
rect 116117 31922 116183 31925
rect 116117 31920 119170 31922
rect 116117 31864 116122 31920
rect 116178 31864 119170 31920
rect 116117 31862 119170 31864
rect 116117 31859 116183 31862
rect 119110 31756 119170 31862
rect 521101 31650 521167 31653
rect 518758 31648 521167 31650
rect 518758 31592 521106 31648
rect 521162 31592 521167 31648
rect 518758 31590 521167 31592
rect 518758 31076 518818 31590
rect 521101 31587 521167 31590
rect 114001 30970 114067 30973
rect 110830 30968 114067 30970
rect 110830 30912 114006 30968
rect 114062 30912 114067 30968
rect 110830 30910 114067 30912
rect 110830 30396 110890 30910
rect 114001 30907 114067 30910
rect 523200 30834 524400 30864
rect 518850 30774 524400 30834
rect 518850 30290 518910 30774
rect 523200 30744 524400 30774
rect 518758 30230 518910 30290
rect 116117 29338 116183 29341
rect 119110 29338 119170 29852
rect 518758 29716 518818 30230
rect 116117 29336 119170 29338
rect 116117 29280 116122 29336
rect 116178 29280 119170 29336
rect 116117 29278 119170 29280
rect 521101 29338 521167 29341
rect 523200 29338 524400 29368
rect 521101 29336 524400 29338
rect 521101 29280 521106 29336
rect 521162 29280 524400 29336
rect 521101 29278 524400 29280
rect 116117 29275 116183 29278
rect 521101 29275 521167 29278
rect 523200 29248 524400 29278
rect 521101 28658 521167 28661
rect 518758 28656 521167 28658
rect 518758 28600 521106 28656
rect 521162 28600 521167 28656
rect 518758 28598 521167 28600
rect 518758 28356 518818 28598
rect 521101 28595 521167 28598
rect 116117 27706 116183 27709
rect 119110 27706 119170 27948
rect 523200 27842 524400 27872
rect 116117 27704 119170 27706
rect 116117 27648 116122 27704
rect 116178 27648 119170 27704
rect 116117 27646 119170 27648
rect 518850 27782 524400 27842
rect 116117 27643 116183 27646
rect 518850 27570 518910 27782
rect 523200 27752 524400 27782
rect 518758 27510 518910 27570
rect 518758 26996 518818 27510
rect 523200 26346 524400 26376
rect 521610 26286 524400 26346
rect 521610 26210 521670 26286
rect 523200 26256 524400 26286
rect 518758 26150 521670 26210
rect 116117 25530 116183 25533
rect 119110 25530 119170 26044
rect 518758 25636 518818 26150
rect 116117 25528 119170 25530
rect 116117 25472 116122 25528
rect 116178 25472 119170 25528
rect 116117 25470 119170 25472
rect 116117 25467 116183 25470
rect 521101 24850 521167 24853
rect 523200 24850 524400 24880
rect 521101 24848 524400 24850
rect 521101 24792 521106 24848
rect 521162 24792 524400 24848
rect 521101 24790 524400 24792
rect 521101 24787 521167 24790
rect 523200 24760 524400 24790
rect 116117 23626 116183 23629
rect 119110 23626 119170 24140
rect 116117 23624 119170 23626
rect 116117 23568 116122 23624
rect 116178 23568 119170 23624
rect 116117 23566 119170 23568
rect 518758 23626 518818 24276
rect 521101 23626 521167 23629
rect 518758 23624 521167 23626
rect 518758 23568 521106 23624
rect 521162 23568 521167 23624
rect 518758 23566 521167 23568
rect 116117 23563 116183 23566
rect 521101 23563 521167 23566
rect 520917 23218 520983 23221
rect 523200 23218 524400 23248
rect 520917 23216 524400 23218
rect 520917 23160 520922 23216
rect 520978 23160 524400 23216
rect 520917 23158 524400 23160
rect 520917 23155 520983 23158
rect 523200 23128 524400 23158
rect 116117 22402 116183 22405
rect 116117 22400 119170 22402
rect 116117 22344 116122 22400
rect 116178 22344 119170 22400
rect 116117 22342 119170 22344
rect 116117 22339 116183 22342
rect 119110 22236 119170 22342
rect 518758 22266 518818 22916
rect 520917 22266 520983 22269
rect 518758 22264 520983 22266
rect 518758 22208 520922 22264
rect 520978 22208 520983 22264
rect 518758 22206 520983 22208
rect 520917 22203 520983 22206
rect 520917 21722 520983 21725
rect 523200 21722 524400 21752
rect 520917 21720 524400 21722
rect 520917 21664 520922 21720
rect 520978 21664 524400 21720
rect 520917 21662 524400 21664
rect 520917 21659 520983 21662
rect 523200 21632 524400 21662
rect 518758 20906 518818 21556
rect 520917 20906 520983 20909
rect 518758 20904 520983 20906
rect 518758 20848 520922 20904
rect 520978 20848 520983 20904
rect 518758 20846 520983 20848
rect 520917 20843 520983 20846
rect 116209 19818 116275 19821
rect 119110 19818 119170 20332
rect 521101 20226 521167 20229
rect 523200 20226 524400 20256
rect 521101 20224 524400 20226
rect 116209 19816 119170 19818
rect 116209 19760 116214 19816
rect 116270 19760 119170 19816
rect 116209 19758 119170 19760
rect 116209 19755 116275 19758
rect 518758 19546 518818 20196
rect 521101 20168 521106 20224
rect 521162 20168 524400 20224
rect 521101 20166 524400 20168
rect 521101 20163 521167 20166
rect 523200 20136 524400 20166
rect 521101 19546 521167 19549
rect 518758 19544 521167 19546
rect 518758 19488 521106 19544
rect 521162 19488 521167 19544
rect 518758 19486 521167 19488
rect 521101 19483 521167 19486
rect 113909 19138 113975 19141
rect 110830 19136 113975 19138
rect 110830 19080 113914 19136
rect 113970 19080 113975 19136
rect 110830 19078 113975 19080
rect 110830 18972 110890 19078
rect 113909 19075 113975 19078
rect 116117 18050 116183 18053
rect 119110 18050 119170 18428
rect 518758 18186 518818 18836
rect 523200 18730 524400 18760
rect 521150 18670 524400 18730
rect 521150 18186 521210 18670
rect 523200 18640 524400 18670
rect 518758 18126 521210 18186
rect 116117 18048 119170 18050
rect 116117 17992 116122 18048
rect 116178 17992 119170 18048
rect 116117 17990 119170 17992
rect 116117 17987 116183 17990
rect 518758 16826 518818 17476
rect 523200 17234 524400 17264
rect 521150 17174 524400 17234
rect 521150 16826 521210 17174
rect 523200 17144 524400 17174
rect 518758 16766 521210 16826
rect 116117 15874 116183 15877
rect 119110 15874 119170 16388
rect 116117 15872 119170 15874
rect 116117 15816 116122 15872
rect 116178 15816 119170 15872
rect 116117 15814 119170 15816
rect 116117 15811 116183 15814
rect 518758 15466 518818 16116
rect 523200 15738 524400 15768
rect 521150 15678 524400 15738
rect 521150 15466 521210 15678
rect 523200 15648 524400 15678
rect 518758 15406 521210 15466
rect 115933 13970 115999 13973
rect 119110 13970 119170 14484
rect 518758 14106 518818 14756
rect 523200 14242 524400 14272
rect 521150 14182 524400 14242
rect 521150 14106 521210 14182
rect 523200 14152 524400 14182
rect 518758 14046 521210 14106
rect 115933 13968 119170 13970
rect 115933 13912 115938 13968
rect 115994 13912 119170 13968
rect 115933 13910 119170 13912
rect 115933 13907 115999 13910
rect 116526 12684 116532 12748
rect 116596 12746 116602 12748
rect 518758 12746 518818 13396
rect 523200 12746 524400 12776
rect 116596 12686 119170 12746
rect 518758 12686 524400 12746
rect 116596 12684 116602 12686
rect 119110 12580 119170 12686
rect 523200 12656 524400 12686
rect 518758 11386 518818 12036
rect 518758 11326 518910 11386
rect 518850 11250 518910 11326
rect 523200 11250 524400 11280
rect 518850 11190 524400 11250
rect 523200 11160 524400 11190
rect 116710 10100 116716 10164
rect 116780 10162 116786 10164
rect 119110 10162 119170 10676
rect 116780 10102 119170 10162
rect 116780 10100 116786 10102
rect 518758 10026 518818 10676
rect 518758 9966 518910 10026
rect 518850 9754 518910 9966
rect 523200 9754 524400 9784
rect 518850 9694 524400 9754
rect 523200 9664 524400 9694
rect 117262 8332 117268 8396
rect 117332 8394 117338 8396
rect 119110 8394 119170 8772
rect 518758 8666 518818 9316
rect 518758 8606 518910 8666
rect 117332 8334 119170 8394
rect 117332 8332 117338 8334
rect 113817 8258 113883 8261
rect 110830 8256 113883 8258
rect 110830 8200 113822 8256
rect 113878 8200 113883 8256
rect 110830 8198 113883 8200
rect 518850 8258 518910 8606
rect 523200 8258 524400 8288
rect 518850 8198 524400 8258
rect 110830 7684 110890 8198
rect 113817 8195 113883 8198
rect 523200 8168 524400 8198
rect 518758 7442 518818 7956
rect 520365 7442 520431 7445
rect 518758 7440 520431 7442
rect 518758 7384 520370 7440
rect 520426 7384 520431 7440
rect 518758 7382 520431 7384
rect 520365 7379 520431 7382
rect 116158 6292 116164 6356
rect 116228 6354 116234 6356
rect 119110 6354 119170 6868
rect 520365 6762 520431 6765
rect 523200 6762 524400 6792
rect 520365 6760 524400 6762
rect 520365 6704 520370 6760
rect 520426 6704 524400 6760
rect 520365 6702 524400 6704
rect 520365 6699 520431 6702
rect 523200 6672 524400 6702
rect 116228 6294 119170 6354
rect 116228 6292 116234 6294
rect 518758 6082 518818 6596
rect 521101 6082 521167 6085
rect 518758 6080 521167 6082
rect 518758 6024 521106 6080
rect 521162 6024 521167 6080
rect 518758 6022 521167 6024
rect 521101 6019 521167 6022
rect 521101 5266 521167 5269
rect 523200 5266 524400 5296
rect 521101 5264 524400 5266
rect 115933 4586 115999 4589
rect 119110 4586 119170 4964
rect 518758 4722 518818 5236
rect 521101 5208 521106 5264
rect 521162 5208 524400 5264
rect 521101 5206 524400 5208
rect 521101 5203 521167 5206
rect 523200 5176 524400 5206
rect 521101 4722 521167 4725
rect 518758 4720 521167 4722
rect 518758 4664 521106 4720
rect 521162 4664 521167 4720
rect 518758 4662 521167 4664
rect 521101 4659 521167 4662
rect 115933 4584 119170 4586
rect 115933 4528 115938 4584
rect 115994 4528 119170 4584
rect 115933 4526 119170 4528
rect 115933 4523 115999 4526
rect 518758 3362 518818 3876
rect 521101 3770 521167 3773
rect 523200 3770 524400 3800
rect 521101 3768 524400 3770
rect 521101 3712 521106 3768
rect 521162 3712 524400 3768
rect 521101 3710 524400 3712
rect 521101 3707 521167 3710
rect 523200 3680 524400 3710
rect 520917 3362 520983 3365
rect 518758 3360 520983 3362
rect 518758 3304 520922 3360
rect 520978 3304 520983 3360
rect 518758 3302 520983 3304
rect 520917 3299 520983 3302
rect 115841 2818 115907 2821
rect 119110 2818 119170 3060
rect 115841 2816 119170 2818
rect 115841 2760 115846 2816
rect 115902 2760 119170 2816
rect 115841 2758 119170 2760
rect 115841 2755 115907 2758
rect 45645 2682 45711 2685
rect 49969 2682 50035 2685
rect 45645 2680 50035 2682
rect 45645 2624 45650 2680
rect 45706 2624 49974 2680
rect 50030 2624 50035 2680
rect 45645 2622 50035 2624
rect 45645 2619 45711 2622
rect 49969 2619 50035 2622
rect 66253 2682 66319 2685
rect 84561 2682 84627 2685
rect 66253 2680 84627 2682
rect 66253 2624 66258 2680
rect 66314 2624 84566 2680
rect 84622 2624 84627 2680
rect 66253 2622 84627 2624
rect 66253 2619 66319 2622
rect 84561 2619 84627 2622
rect 106089 2682 106155 2685
rect 109585 2682 109651 2685
rect 106089 2680 109651 2682
rect 106089 2624 106094 2680
rect 106150 2624 109590 2680
rect 109646 2624 109651 2680
rect 106089 2622 109651 2624
rect 106089 2619 106155 2622
rect 109585 2619 109651 2622
rect 64873 2546 64939 2549
rect 85849 2546 85915 2549
rect 64873 2544 85915 2546
rect 64873 2488 64878 2544
rect 64934 2488 85854 2544
rect 85910 2488 85915 2544
rect 64873 2486 85915 2488
rect 64873 2483 64939 2486
rect 85849 2483 85915 2486
rect 67541 2410 67607 2413
rect 85297 2410 85363 2413
rect 67541 2408 85363 2410
rect 67541 2352 67546 2408
rect 67602 2352 85302 2408
rect 85358 2352 85363 2408
rect 67541 2350 85363 2352
rect 67541 2347 67607 2350
rect 85297 2347 85363 2350
rect 69013 2274 69079 2277
rect 76465 2274 76531 2277
rect 69013 2272 76531 2274
rect 69013 2216 69018 2272
rect 69074 2216 76470 2272
rect 76526 2216 76531 2272
rect 69013 2214 76531 2216
rect 69013 2211 69079 2214
rect 76465 2211 76531 2214
rect 518758 2138 518818 2652
rect 520917 2274 520983 2277
rect 523200 2274 524400 2304
rect 520917 2272 524400 2274
rect 520917 2216 520922 2272
rect 520978 2216 524400 2272
rect 520917 2214 524400 2216
rect 520917 2211 520983 2214
rect 523200 2184 524400 2214
rect 521101 2138 521167 2141
rect 518758 2136 521167 2138
rect 518758 2080 521106 2136
rect 521162 2080 521167 2136
rect 518758 2078 521167 2080
rect 521101 2075 521167 2078
rect 19333 1866 19399 1869
rect 116526 1866 116532 1868
rect 19333 1864 116532 1866
rect 19333 1808 19338 1864
rect 19394 1808 116532 1864
rect 19333 1806 116532 1808
rect 19333 1803 19399 1806
rect 116526 1804 116532 1806
rect 116596 1804 116602 1868
rect 15929 1730 15995 1733
rect 116710 1730 116716 1732
rect 15929 1728 116716 1730
rect 15929 1672 15934 1728
rect 15990 1672 116716 1728
rect 15929 1670 116716 1672
rect 15929 1667 15995 1670
rect 116710 1668 116716 1670
rect 116780 1668 116786 1732
rect 12617 1594 12683 1597
rect 117262 1594 117268 1596
rect 12617 1592 117268 1594
rect 12617 1536 12622 1592
rect 12678 1536 117268 1592
rect 12617 1534 117268 1536
rect 12617 1531 12683 1534
rect 117262 1532 117268 1534
rect 117332 1532 117338 1596
rect 229277 1594 229343 1597
rect 293585 1594 293651 1597
rect 229277 1592 293651 1594
rect 229277 1536 229282 1592
rect 229338 1536 293590 1592
rect 293646 1536 293651 1592
rect 229277 1534 293651 1536
rect 229277 1531 229343 1534
rect 293585 1531 293651 1534
rect 9305 1458 9371 1461
rect 116158 1458 116164 1460
rect 9305 1456 116164 1458
rect 9305 1400 9310 1456
rect 9366 1400 116164 1456
rect 9305 1398 116164 1400
rect 9305 1395 9371 1398
rect 116158 1396 116164 1398
rect 116228 1396 116234 1460
rect 163773 1458 163839 1461
rect 243629 1458 243695 1461
rect 163773 1456 243695 1458
rect 163773 1400 163778 1456
rect 163834 1400 243634 1456
rect 243690 1400 243695 1456
rect 163773 1398 243695 1400
rect 163773 1395 163839 1398
rect 243629 1395 243695 1398
rect 360285 1458 360351 1461
rect 393589 1458 393655 1461
rect 360285 1456 393655 1458
rect 360285 1400 360290 1456
rect 360346 1400 393594 1456
rect 393650 1400 393655 1456
rect 360285 1398 393655 1400
rect 360285 1395 360351 1398
rect 393589 1395 393655 1398
rect 521101 778 521167 781
rect 523200 778 524400 808
rect 521101 776 524400 778
rect 521101 720 521106 776
rect 521162 720 524400 776
rect 521101 718 524400 720
rect 521101 715 521167 718
rect 523200 688 524400 718
<< via3 >>
rect 116532 12684 116596 12748
rect 116716 10100 116780 10164
rect 117268 8332 117332 8396
rect 116164 6292 116228 6356
rect 116532 1804 116596 1868
rect 116716 1668 116780 1732
rect 117268 1532 117332 1596
rect 116164 1396 116228 1460
<< metal4 >>
rect 1664 144454 1984 144496
rect 1664 144218 1706 144454
rect 1942 144218 1984 144454
rect 1664 144134 1984 144218
rect 1664 143898 1706 144134
rect 1942 143898 1984 144134
rect 1664 143856 1984 143898
rect 109956 144454 110276 144496
rect 109956 144218 109998 144454
rect 110234 144218 110276 144454
rect 109956 144134 110276 144218
rect 109956 143898 109998 144134
rect 110234 143898 110276 144134
rect 109956 143856 110276 143898
rect 119664 144454 119984 144496
rect 119664 144218 119706 144454
rect 119942 144218 119984 144454
rect 119664 144134 119984 144218
rect 119664 143898 119706 144134
rect 119942 143898 119984 144134
rect 119664 143856 119984 143898
rect 517940 144454 518260 144496
rect 517940 144218 517982 144454
rect 518218 144218 518260 144454
rect 517940 144134 518260 144218
rect 517940 143898 517982 144134
rect 518218 143898 518260 144134
rect 517940 143856 518260 143898
rect 1096 131454 1332 131496
rect 1096 131134 1332 131218
rect 1096 130856 1332 130898
rect 110616 131454 110936 131496
rect 110616 131218 110658 131454
rect 110894 131218 110936 131454
rect 110616 131134 110936 131218
rect 110616 130898 110658 131134
rect 110894 130898 110936 131134
rect 110616 130856 110936 130898
rect 119004 131454 119324 131496
rect 119004 131218 119046 131454
rect 119282 131218 119324 131454
rect 119004 131134 119324 131218
rect 119004 130898 119046 131134
rect 119282 130898 119324 131134
rect 119004 130856 119324 130898
rect 518600 131454 518920 131496
rect 518600 131218 518642 131454
rect 518878 131218 518920 131454
rect 518600 131134 518920 131218
rect 518600 130898 518642 131134
rect 518878 130898 518920 131134
rect 518600 130856 518920 130898
rect 1664 118454 1984 118496
rect 1664 118218 1706 118454
rect 1942 118218 1984 118454
rect 1664 118134 1984 118218
rect 1664 117898 1706 118134
rect 1942 117898 1984 118134
rect 1664 117856 1984 117898
rect 109956 118454 110276 118496
rect 109956 118218 109998 118454
rect 110234 118218 110276 118454
rect 109956 118134 110276 118218
rect 109956 117898 109998 118134
rect 110234 117898 110276 118134
rect 109956 117856 110276 117898
rect 119664 118454 119984 118496
rect 119664 118218 119706 118454
rect 119942 118218 119984 118454
rect 119664 118134 119984 118218
rect 119664 117898 119706 118134
rect 119942 117898 119984 118134
rect 119664 117856 119984 117898
rect 517940 118454 518260 118496
rect 517940 118218 517982 118454
rect 518218 118218 518260 118454
rect 517940 118134 518260 118218
rect 517940 117898 517982 118134
rect 518218 117898 518260 118134
rect 517940 117856 518260 117898
rect 1096 105454 1332 105496
rect 1096 105134 1332 105218
rect 1096 104856 1332 104898
rect 110616 105454 110936 105496
rect 110616 105218 110658 105454
rect 110894 105218 110936 105454
rect 110616 105134 110936 105218
rect 110616 104898 110658 105134
rect 110894 104898 110936 105134
rect 110616 104856 110936 104898
rect 119004 105454 119324 105496
rect 119004 105218 119046 105454
rect 119282 105218 119324 105454
rect 119004 105134 119324 105218
rect 119004 104898 119046 105134
rect 119282 104898 119324 105134
rect 119004 104856 119324 104898
rect 518600 105454 518920 105496
rect 518600 105218 518642 105454
rect 518878 105218 518920 105454
rect 518600 105134 518920 105218
rect 518600 104898 518642 105134
rect 518878 104898 518920 105134
rect 518600 104856 518920 104898
rect 1664 92454 1984 92496
rect 1664 92218 1706 92454
rect 1942 92218 1984 92454
rect 1664 92134 1984 92218
rect 1664 91898 1706 92134
rect 1942 91898 1984 92134
rect 1664 91856 1984 91898
rect 109956 92454 110276 92496
rect 109956 92218 109998 92454
rect 110234 92218 110276 92454
rect 109956 92134 110276 92218
rect 109956 91898 109998 92134
rect 110234 91898 110276 92134
rect 109956 91856 110276 91898
rect 119664 92454 119984 92496
rect 119664 92218 119706 92454
rect 119942 92218 119984 92454
rect 119664 92134 119984 92218
rect 119664 91898 119706 92134
rect 119942 91898 119984 92134
rect 119664 91856 119984 91898
rect 517940 92454 518260 92496
rect 517940 92218 517982 92454
rect 518218 92218 518260 92454
rect 517940 92134 518260 92218
rect 517940 91898 517982 92134
rect 518218 91898 518260 92134
rect 517940 91856 518260 91898
rect 1096 79454 1332 79496
rect 1096 79134 1332 79218
rect 1096 78856 1332 78898
rect 110616 79454 110936 79496
rect 110616 79218 110658 79454
rect 110894 79218 110936 79454
rect 110616 79134 110936 79218
rect 110616 78898 110658 79134
rect 110894 78898 110936 79134
rect 110616 78856 110936 78898
rect 119004 79454 119324 79496
rect 119004 79218 119046 79454
rect 119282 79218 119324 79454
rect 119004 79134 119324 79218
rect 119004 78898 119046 79134
rect 119282 78898 119324 79134
rect 119004 78856 119324 78898
rect 518600 79454 518920 79496
rect 518600 79218 518642 79454
rect 518878 79218 518920 79454
rect 518600 79134 518920 79218
rect 518600 78898 518642 79134
rect 518878 78898 518920 79134
rect 518600 78856 518920 78898
rect 1664 66454 1984 66496
rect 1664 66218 1706 66454
rect 1942 66218 1984 66454
rect 1664 66134 1984 66218
rect 1664 65898 1706 66134
rect 1942 65898 1984 66134
rect 1664 65856 1984 65898
rect 109956 66454 110276 66496
rect 109956 66218 109998 66454
rect 110234 66218 110276 66454
rect 109956 66134 110276 66218
rect 109956 65898 109998 66134
rect 110234 65898 110276 66134
rect 109956 65856 110276 65898
rect 119664 66454 119984 66496
rect 119664 66218 119706 66454
rect 119942 66218 119984 66454
rect 119664 66134 119984 66218
rect 119664 65898 119706 66134
rect 119942 65898 119984 66134
rect 119664 65856 119984 65898
rect 517940 66454 518260 66496
rect 517940 66218 517982 66454
rect 518218 66218 518260 66454
rect 517940 66134 518260 66218
rect 517940 65898 517982 66134
rect 518218 65898 518260 66134
rect 517940 65856 518260 65898
rect 1096 53454 1332 53496
rect 1096 53134 1332 53218
rect 1096 52856 1332 52898
rect 110616 53454 110936 53496
rect 110616 53218 110658 53454
rect 110894 53218 110936 53454
rect 110616 53134 110936 53218
rect 110616 52898 110658 53134
rect 110894 52898 110936 53134
rect 110616 52856 110936 52898
rect 119004 53454 119324 53496
rect 119004 53218 119046 53454
rect 119282 53218 119324 53454
rect 119004 53134 119324 53218
rect 119004 52898 119046 53134
rect 119282 52898 119324 53134
rect 119004 52856 119324 52898
rect 518600 53454 518920 53496
rect 518600 53218 518642 53454
rect 518878 53218 518920 53454
rect 518600 53134 518920 53218
rect 518600 52898 518642 53134
rect 518878 52898 518920 53134
rect 518600 52856 518920 52898
rect 1664 40454 1984 40496
rect 1664 40218 1706 40454
rect 1942 40218 1984 40454
rect 1664 40134 1984 40218
rect 1664 39898 1706 40134
rect 1942 39898 1984 40134
rect 1664 39856 1984 39898
rect 109956 40454 110276 40496
rect 109956 40218 109998 40454
rect 110234 40218 110276 40454
rect 109956 40134 110276 40218
rect 109956 39898 109998 40134
rect 110234 39898 110276 40134
rect 109956 39856 110276 39898
rect 119664 40454 119984 40496
rect 119664 40218 119706 40454
rect 119942 40218 119984 40454
rect 119664 40134 119984 40218
rect 119664 39898 119706 40134
rect 119942 39898 119984 40134
rect 119664 39856 119984 39898
rect 517940 40454 518260 40496
rect 517940 40218 517982 40454
rect 518218 40218 518260 40454
rect 517940 40134 518260 40218
rect 517940 39898 517982 40134
rect 518218 39898 518260 40134
rect 517940 39856 518260 39898
rect 1096 27454 1332 27496
rect 1096 27134 1332 27218
rect 1096 26856 1332 26898
rect 110616 27454 110936 27496
rect 110616 27218 110658 27454
rect 110894 27218 110936 27454
rect 110616 27134 110936 27218
rect 110616 26898 110658 27134
rect 110894 26898 110936 27134
rect 110616 26856 110936 26898
rect 119004 27454 119324 27496
rect 119004 27218 119046 27454
rect 119282 27218 119324 27454
rect 119004 27134 119324 27218
rect 119004 26898 119046 27134
rect 119282 26898 119324 27134
rect 119004 26856 119324 26898
rect 518600 27454 518920 27496
rect 518600 27218 518642 27454
rect 518878 27218 518920 27454
rect 518600 27134 518920 27218
rect 518600 26898 518642 27134
rect 518878 26898 518920 27134
rect 518600 26856 518920 26898
rect 1664 14454 1984 14496
rect 1664 14218 1706 14454
rect 1942 14218 1984 14454
rect 1664 14134 1984 14218
rect 1664 13898 1706 14134
rect 1942 13898 1984 14134
rect 1664 13856 1984 13898
rect 109956 14454 110276 14496
rect 109956 14218 109998 14454
rect 110234 14218 110276 14454
rect 109956 14134 110276 14218
rect 109956 13898 109998 14134
rect 110234 13898 110276 14134
rect 109956 13856 110276 13898
rect 119664 14454 119984 14496
rect 119664 14218 119706 14454
rect 119942 14218 119984 14454
rect 119664 14134 119984 14218
rect 119664 13898 119706 14134
rect 119942 13898 119984 14134
rect 119664 13856 119984 13898
rect 517940 14454 518260 14496
rect 517940 14218 517982 14454
rect 518218 14218 518260 14454
rect 517940 14134 518260 14218
rect 517940 13898 517982 14134
rect 518218 13898 518260 14134
rect 517940 13856 518260 13898
rect 116531 12748 116597 12749
rect 116531 12684 116532 12748
rect 116596 12684 116597 12748
rect 116531 12683 116597 12684
rect 116163 6356 116229 6357
rect 116163 6292 116164 6356
rect 116228 6292 116229 6356
rect 116163 6291 116229 6292
rect 116166 1461 116226 6291
rect 116534 1869 116594 12683
rect 116715 10164 116781 10165
rect 116715 10100 116716 10164
rect 116780 10100 116781 10164
rect 116715 10099 116781 10100
rect 116531 1868 116597 1869
rect 116531 1804 116532 1868
rect 116596 1804 116597 1868
rect 116531 1803 116597 1804
rect 116718 1733 116778 10099
rect 117267 8396 117333 8397
rect 117267 8332 117268 8396
rect 117332 8332 117333 8396
rect 117267 8331 117333 8332
rect 116715 1732 116781 1733
rect 116715 1668 116716 1732
rect 116780 1668 116781 1732
rect 116715 1667 116781 1668
rect 117270 1597 117330 8331
rect 117267 1596 117333 1597
rect 117267 1532 117268 1596
rect 117332 1532 117333 1596
rect 117267 1531 117333 1532
rect 116163 1460 116229 1461
rect 116163 1396 116164 1460
rect 116228 1396 116229 1460
rect 116163 1395 116229 1396
<< via4 >>
rect 1706 144218 1942 144454
rect 1706 143898 1942 144134
rect 109998 144218 110234 144454
rect 109998 143898 110234 144134
rect 119706 144218 119942 144454
rect 119706 143898 119942 144134
rect 517982 144218 518218 144454
rect 517982 143898 518218 144134
rect 1096 131218 1332 131454
rect 1096 130898 1332 131134
rect 110658 131218 110894 131454
rect 110658 130898 110894 131134
rect 119046 131218 119282 131454
rect 119046 130898 119282 131134
rect 518642 131218 518878 131454
rect 518642 130898 518878 131134
rect 1706 118218 1942 118454
rect 1706 117898 1942 118134
rect 109998 118218 110234 118454
rect 109998 117898 110234 118134
rect 119706 118218 119942 118454
rect 119706 117898 119942 118134
rect 517982 118218 518218 118454
rect 517982 117898 518218 118134
rect 1096 105218 1332 105454
rect 1096 104898 1332 105134
rect 110658 105218 110894 105454
rect 110658 104898 110894 105134
rect 119046 105218 119282 105454
rect 119046 104898 119282 105134
rect 518642 105218 518878 105454
rect 518642 104898 518878 105134
rect 1706 92218 1942 92454
rect 1706 91898 1942 92134
rect 109998 92218 110234 92454
rect 109998 91898 110234 92134
rect 119706 92218 119942 92454
rect 119706 91898 119942 92134
rect 517982 92218 518218 92454
rect 517982 91898 518218 92134
rect 1096 79218 1332 79454
rect 1096 78898 1332 79134
rect 110658 79218 110894 79454
rect 110658 78898 110894 79134
rect 119046 79218 119282 79454
rect 119046 78898 119282 79134
rect 518642 79218 518878 79454
rect 518642 78898 518878 79134
rect 1706 66218 1942 66454
rect 1706 65898 1942 66134
rect 109998 66218 110234 66454
rect 109998 65898 110234 66134
rect 119706 66218 119942 66454
rect 119706 65898 119942 66134
rect 517982 66218 518218 66454
rect 517982 65898 518218 66134
rect 1096 53218 1332 53454
rect 1096 52898 1332 53134
rect 110658 53218 110894 53454
rect 110658 52898 110894 53134
rect 119046 53218 119282 53454
rect 119046 52898 119282 53134
rect 518642 53218 518878 53454
rect 518642 52898 518878 53134
rect 1706 40218 1942 40454
rect 1706 39898 1942 40134
rect 109998 40218 110234 40454
rect 109998 39898 110234 40134
rect 119706 40218 119942 40454
rect 119706 39898 119942 40134
rect 517982 40218 518218 40454
rect 517982 39898 518218 40134
rect 1096 27218 1332 27454
rect 1096 26898 1332 27134
rect 110658 27218 110894 27454
rect 110658 26898 110894 27134
rect 119046 27218 119282 27454
rect 119046 26898 119282 27134
rect 518642 27218 518878 27454
rect 518642 26898 518878 27134
rect 1706 14218 1942 14454
rect 1706 13898 1942 14134
rect 109998 14218 110234 14454
rect 109998 13898 110234 14134
rect 119706 14218 119942 14454
rect 119706 13898 119942 14134
rect 517982 14218 518218 14454
rect 517982 13898 518218 14134
<< metal5 >>
rect 1104 156856 522836 157496
rect 1104 144454 2200 144496
rect 1104 144218 1706 144454
rect 1942 144218 2200 144454
rect 1104 144134 2200 144218
rect 1104 143898 1706 144134
rect 1942 143898 2200 144134
rect 1104 143856 2200 143898
rect 109800 144454 120200 144496
rect 109800 144218 109998 144454
rect 110234 144218 119706 144454
rect 119942 144218 120200 144454
rect 109800 144134 120200 144218
rect 109800 143898 109998 144134
rect 110234 143898 119706 144134
rect 119942 143898 120200 144134
rect 109800 143856 120200 143898
rect 517800 144454 522836 144496
rect 517800 144218 517982 144454
rect 518218 144218 522836 144454
rect 517800 144134 522836 144218
rect 517800 143898 517982 144134
rect 518218 143898 522836 144134
rect 517800 143856 522836 143898
rect 1072 131454 2200 131496
rect 1072 131218 1096 131454
rect 1332 131218 2200 131454
rect 1072 131134 2200 131218
rect 1072 130898 1096 131134
rect 1332 130898 2200 131134
rect 1072 130856 2200 130898
rect 109800 131454 120200 131496
rect 109800 131218 110658 131454
rect 110894 131218 119046 131454
rect 119282 131218 120200 131454
rect 109800 131134 120200 131218
rect 109800 130898 110658 131134
rect 110894 130898 119046 131134
rect 119282 130898 120200 131134
rect 109800 130856 120200 130898
rect 517800 131454 522836 131496
rect 517800 131218 518642 131454
rect 518878 131218 522836 131454
rect 517800 131134 522836 131218
rect 517800 130898 518642 131134
rect 518878 130898 522836 131134
rect 517800 130856 522836 130898
rect 1104 118454 2200 118496
rect 1104 118218 1706 118454
rect 1942 118218 2200 118454
rect 1104 118134 2200 118218
rect 1104 117898 1706 118134
rect 1942 117898 2200 118134
rect 1104 117856 2200 117898
rect 109800 118454 120200 118496
rect 109800 118218 109998 118454
rect 110234 118218 119706 118454
rect 119942 118218 120200 118454
rect 109800 118134 120200 118218
rect 109800 117898 109998 118134
rect 110234 117898 119706 118134
rect 119942 117898 120200 118134
rect 109800 117856 120200 117898
rect 517800 118454 522836 118496
rect 517800 118218 517982 118454
rect 518218 118218 522836 118454
rect 517800 118134 522836 118218
rect 517800 117898 517982 118134
rect 518218 117898 522836 118134
rect 517800 117856 522836 117898
rect 1072 105454 2200 105496
rect 1072 105218 1096 105454
rect 1332 105218 2200 105454
rect 1072 105134 2200 105218
rect 1072 104898 1096 105134
rect 1332 104898 2200 105134
rect 1072 104856 2200 104898
rect 109800 105454 120200 105496
rect 109800 105218 110658 105454
rect 110894 105218 119046 105454
rect 119282 105218 120200 105454
rect 109800 105134 120200 105218
rect 109800 104898 110658 105134
rect 110894 104898 119046 105134
rect 119282 104898 120200 105134
rect 109800 104856 120200 104898
rect 517800 105454 522836 105496
rect 517800 105218 518642 105454
rect 518878 105218 522836 105454
rect 517800 105134 522836 105218
rect 517800 104898 518642 105134
rect 518878 104898 522836 105134
rect 517800 104856 522836 104898
rect 1104 92454 2200 92496
rect 1104 92218 1706 92454
rect 1942 92218 2200 92454
rect 1104 92134 2200 92218
rect 1104 91898 1706 92134
rect 1942 91898 2200 92134
rect 1104 91856 2200 91898
rect 109800 92454 120200 92496
rect 109800 92218 109998 92454
rect 110234 92218 119706 92454
rect 119942 92218 120200 92454
rect 109800 92134 120200 92218
rect 109800 91898 109998 92134
rect 110234 91898 119706 92134
rect 119942 91898 120200 92134
rect 109800 91856 120200 91898
rect 517800 92454 522836 92496
rect 517800 92218 517982 92454
rect 518218 92218 522836 92454
rect 517800 92134 522836 92218
rect 517800 91898 517982 92134
rect 518218 91898 522836 92134
rect 517800 91856 522836 91898
rect 1072 79454 2200 79496
rect 1072 79218 1096 79454
rect 1332 79218 2200 79454
rect 1072 79134 2200 79218
rect 1072 78898 1096 79134
rect 1332 78898 2200 79134
rect 1072 78856 2200 78898
rect 109800 79454 120200 79496
rect 109800 79218 110658 79454
rect 110894 79218 119046 79454
rect 119282 79218 120200 79454
rect 109800 79134 120200 79218
rect 109800 78898 110658 79134
rect 110894 78898 119046 79134
rect 119282 78898 120200 79134
rect 109800 78856 120200 78898
rect 517800 79454 522836 79496
rect 517800 79218 518642 79454
rect 518878 79218 522836 79454
rect 517800 79134 522836 79218
rect 517800 78898 518642 79134
rect 518878 78898 522836 79134
rect 517800 78856 522836 78898
rect 1104 66454 2200 66496
rect 1104 66218 1706 66454
rect 1942 66218 2200 66454
rect 1104 66134 2200 66218
rect 1104 65898 1706 66134
rect 1942 65898 2200 66134
rect 1104 65856 2200 65898
rect 109800 66454 120200 66496
rect 109800 66218 109998 66454
rect 110234 66218 119706 66454
rect 119942 66218 120200 66454
rect 109800 66134 120200 66218
rect 109800 65898 109998 66134
rect 110234 65898 119706 66134
rect 119942 65898 120200 66134
rect 109800 65856 120200 65898
rect 517800 66454 522836 66496
rect 517800 66218 517982 66454
rect 518218 66218 522836 66454
rect 517800 66134 522836 66218
rect 517800 65898 517982 66134
rect 518218 65898 522836 66134
rect 517800 65856 522836 65898
rect 1072 53454 2200 53496
rect 1072 53218 1096 53454
rect 1332 53218 2200 53454
rect 1072 53134 2200 53218
rect 1072 52898 1096 53134
rect 1332 52898 2200 53134
rect 1072 52856 2200 52898
rect 109800 53454 120200 53496
rect 109800 53218 110658 53454
rect 110894 53218 119046 53454
rect 119282 53218 120200 53454
rect 109800 53134 120200 53218
rect 109800 52898 110658 53134
rect 110894 52898 119046 53134
rect 119282 52898 120200 53134
rect 109800 52856 120200 52898
rect 517800 53454 522836 53496
rect 517800 53218 518642 53454
rect 518878 53218 522836 53454
rect 517800 53134 522836 53218
rect 517800 52898 518642 53134
rect 518878 52898 522836 53134
rect 517800 52856 522836 52898
rect 1104 40454 2200 40496
rect 1104 40218 1706 40454
rect 1942 40218 2200 40454
rect 1104 40134 2200 40218
rect 1104 39898 1706 40134
rect 1942 39898 2200 40134
rect 1104 39856 2200 39898
rect 109800 40454 120200 40496
rect 109800 40218 109998 40454
rect 110234 40218 119706 40454
rect 119942 40218 120200 40454
rect 109800 40134 120200 40218
rect 109800 39898 109998 40134
rect 110234 39898 119706 40134
rect 119942 39898 120200 40134
rect 109800 39856 120200 39898
rect 517800 40454 522836 40496
rect 517800 40218 517982 40454
rect 518218 40218 522836 40454
rect 517800 40134 522836 40218
rect 517800 39898 517982 40134
rect 518218 39898 522836 40134
rect 517800 39856 522836 39898
rect 1072 27454 2200 27496
rect 1072 27218 1096 27454
rect 1332 27218 2200 27454
rect 1072 27134 2200 27218
rect 1072 26898 1096 27134
rect 1332 26898 2200 27134
rect 1072 26856 2200 26898
rect 109800 27454 120200 27496
rect 109800 27218 110658 27454
rect 110894 27218 119046 27454
rect 119282 27218 120200 27454
rect 109800 27134 120200 27218
rect 109800 26898 110658 27134
rect 110894 26898 119046 27134
rect 119282 26898 120200 27134
rect 109800 26856 120200 26898
rect 517800 27454 522836 27496
rect 517800 27218 518642 27454
rect 518878 27218 522836 27454
rect 517800 27134 522836 27218
rect 517800 26898 518642 27134
rect 518878 26898 522836 27134
rect 517800 26856 522836 26898
rect 1104 14454 2200 14496
rect 1104 14218 1706 14454
rect 1942 14218 2200 14454
rect 1104 14134 2200 14218
rect 1104 13898 1706 14134
rect 1942 13898 2200 14134
rect 1104 13856 2200 13898
rect 109800 14454 120200 14496
rect 109800 14218 109998 14454
rect 110234 14218 119706 14454
rect 119942 14218 120200 14454
rect 109800 14134 120200 14218
rect 109800 13898 109998 14134
rect 110234 13898 119706 14134
rect 119942 13898 120200 14134
rect 109800 13856 120200 13898
rect 517800 14454 522836 14496
rect 517800 14218 517982 14454
rect 518218 14218 522836 14454
rect 517800 14134 522836 14218
rect 517800 13898 517982 14134
rect 518218 13898 522836 14134
rect 517800 13856 522836 13898
use mgmt_core  core
timestamp 1640295518
transform 1 0 119000 0 1 2000
box 0 0 400000 148000
use DFFRAM  DFFRAM
timestamp 1640295518
transform 1 0 1000 0 1 2000
box 4 0 110000 148000
<< labels >>
rlabel metal5 s 1104 26856 2200 27496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 26856 120200 27496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 26856 522836 27496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 52856 2200 53496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 52856 120200 53496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 52856 522836 53496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 78856 2200 79496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 78856 120200 79496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 78856 522836 79496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 104856 2200 105496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 104856 120200 105496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 104856 522836 105496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 130856 2200 131496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 130856 120200 131496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 130856 522836 131496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 156856 522836 157496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 13856 2200 14496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 13856 120200 14496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 13856 522836 14496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 39856 2200 40496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 39856 120200 40496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 39856 522836 40496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 65856 2200 66496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 65856 120200 66496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 65856 522836 66496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 91856 2200 92496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 91856 120200 92496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 91856 522836 92496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 117856 2200 118496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 117856 120200 118496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 117856 522836 118496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 143856 2200 144496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 143856 120200 144496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 143856 522836 144496 6 VPWR
port 1 nsew power input
rlabel metal2 s 294786 -400 294842 800 6 core_clk
port 2 nsew signal input
rlabel metal2 s 98274 -400 98330 800 6 core_rstn
port 3 nsew signal input
rlabel metal3 s 523200 63792 524400 63912 6 debug_in
port 4 nsew signal input
rlabel metal3 s 523200 65288 524400 65408 6 debug_mode
port 5 nsew signal tristate
rlabel metal3 s 523200 66784 524400 66904 6 debug_oeb
port 6 nsew signal tristate
rlabel metal3 s 523200 68280 524400 68400 6 debug_out
port 7 nsew signal tristate
rlabel metal3 s 523200 145120 524400 145240 6 flash_clk
port 8 nsew signal tristate
rlabel metal3 s 523200 143624 524400 143744 6 flash_csb
port 9 nsew signal tristate
rlabel metal3 s 523200 146616 524400 146736 6 flash_io0_di
port 10 nsew signal input
rlabel metal3 s 523200 148112 524400 148232 6 flash_io0_do
port 11 nsew signal tristate
rlabel metal3 s 523200 149608 524400 149728 6 flash_io0_oeb
port 12 nsew signal tristate
rlabel metal3 s 523200 151104 524400 151224 6 flash_io1_di
port 13 nsew signal input
rlabel metal3 s 523200 152600 524400 152720 6 flash_io1_do
port 14 nsew signal tristate
rlabel metal3 s 523200 154096 524400 154216 6 flash_io1_oeb
port 15 nsew signal tristate
rlabel metal3 s 523200 155592 524400 155712 6 flash_io2_di
port 16 nsew signal input
rlabel metal3 s 523200 157088 524400 157208 6 flash_io2_do
port 17 nsew signal tristate
rlabel metal3 s 523200 158584 524400 158704 6 flash_io2_oeb
port 18 nsew signal tristate
rlabel metal3 s 523200 160080 524400 160200 6 flash_io3_di
port 19 nsew signal input
rlabel metal3 s 523200 161576 524400 161696 6 flash_io3_do
port 20 nsew signal tristate
rlabel metal3 s 523200 163072 524400 163192 6 flash_io3_oeb
port 21 nsew signal tristate
rlabel metal2 s 32770 -400 32826 800 6 gpio_in_pad
port 22 nsew signal input
rlabel metal2 s 163778 -400 163834 800 6 gpio_inenb_pad
port 23 nsew signal tristate
rlabel metal2 s 229282 -400 229338 800 6 gpio_mode0_pad
port 24 nsew signal tristate
rlabel metal2 s 360290 -400 360346 800 6 gpio_mode1_pad
port 25 nsew signal tristate
rlabel metal2 s 425794 -400 425850 800 6 gpio_out_pad
port 26 nsew signal tristate
rlabel metal2 s 491298 -400 491354 800 6 gpio_outenb_pad
port 27 nsew signal tristate
rlabel metal3 s 523200 90856 524400 90976 6 hk_ack_i
port 28 nsew signal input
rlabel metal3 s 523200 93848 524400 93968 6 hk_cyc_o
port 29 nsew signal tristate
rlabel metal3 s 523200 95480 524400 95600 6 hk_dat_i[0]
port 30 nsew signal input
rlabel metal3 s 523200 110440 524400 110560 6 hk_dat_i[10]
port 31 nsew signal input
rlabel metal3 s 523200 111936 524400 112056 6 hk_dat_i[11]
port 32 nsew signal input
rlabel metal3 s 523200 113432 524400 113552 6 hk_dat_i[12]
port 33 nsew signal input
rlabel metal3 s 523200 114928 524400 115048 6 hk_dat_i[13]
port 34 nsew signal input
rlabel metal3 s 523200 116424 524400 116544 6 hk_dat_i[14]
port 35 nsew signal input
rlabel metal3 s 523200 118056 524400 118176 6 hk_dat_i[15]
port 36 nsew signal input
rlabel metal3 s 523200 119552 524400 119672 6 hk_dat_i[16]
port 37 nsew signal input
rlabel metal3 s 523200 121048 524400 121168 6 hk_dat_i[17]
port 38 nsew signal input
rlabel metal3 s 523200 122544 524400 122664 6 hk_dat_i[18]
port 39 nsew signal input
rlabel metal3 s 523200 124040 524400 124160 6 hk_dat_i[19]
port 40 nsew signal input
rlabel metal3 s 523200 96976 524400 97096 6 hk_dat_i[1]
port 41 nsew signal input
rlabel metal3 s 523200 125536 524400 125656 6 hk_dat_i[20]
port 42 nsew signal input
rlabel metal3 s 523200 127032 524400 127152 6 hk_dat_i[21]
port 43 nsew signal input
rlabel metal3 s 523200 128528 524400 128648 6 hk_dat_i[22]
port 44 nsew signal input
rlabel metal3 s 523200 130024 524400 130144 6 hk_dat_i[23]
port 45 nsew signal input
rlabel metal3 s 523200 131520 524400 131640 6 hk_dat_i[24]
port 46 nsew signal input
rlabel metal3 s 523200 133016 524400 133136 6 hk_dat_i[25]
port 47 nsew signal input
rlabel metal3 s 523200 134512 524400 134632 6 hk_dat_i[26]
port 48 nsew signal input
rlabel metal3 s 523200 136008 524400 136128 6 hk_dat_i[27]
port 49 nsew signal input
rlabel metal3 s 523200 137504 524400 137624 6 hk_dat_i[28]
port 50 nsew signal input
rlabel metal3 s 523200 139000 524400 139120 6 hk_dat_i[29]
port 51 nsew signal input
rlabel metal3 s 523200 98472 524400 98592 6 hk_dat_i[2]
port 52 nsew signal input
rlabel metal3 s 523200 140496 524400 140616 6 hk_dat_i[30]
port 53 nsew signal input
rlabel metal3 s 523200 142128 524400 142248 6 hk_dat_i[31]
port 54 nsew signal input
rlabel metal3 s 523200 99968 524400 100088 6 hk_dat_i[3]
port 55 nsew signal input
rlabel metal3 s 523200 101464 524400 101584 6 hk_dat_i[4]
port 56 nsew signal input
rlabel metal3 s 523200 102960 524400 103080 6 hk_dat_i[5]
port 57 nsew signal input
rlabel metal3 s 523200 104456 524400 104576 6 hk_dat_i[6]
port 58 nsew signal input
rlabel metal3 s 523200 105952 524400 106072 6 hk_dat_i[7]
port 59 nsew signal input
rlabel metal3 s 523200 107448 524400 107568 6 hk_dat_i[8]
port 60 nsew signal input
rlabel metal3 s 523200 108944 524400 109064 6 hk_dat_i[9]
port 61 nsew signal input
rlabel metal3 s 523200 92352 524400 92472 6 hk_stb_o
port 62 nsew signal tristate
rlabel metal2 s 521842 163200 521898 164400 6 irq[0]
port 63 nsew signal input
rlabel metal2 s 522670 163200 522726 164400 6 irq[1]
port 64 nsew signal input
rlabel metal2 s 523498 163200 523554 164400 6 irq[2]
port 65 nsew signal input
rlabel metal3 s 523200 74400 524400 74520 6 irq[3]
port 66 nsew signal input
rlabel metal3 s 523200 72904 524400 73024 6 irq[4]
port 67 nsew signal input
rlabel metal3 s 523200 71408 524400 71528 6 irq[5]
port 68 nsew signal input
rlabel metal2 s 386 163200 442 164400 6 la_iena[0]
port 69 nsew signal tristate
rlabel metal2 s 336830 163200 336886 164400 6 la_iena[100]
port 70 nsew signal tristate
rlabel metal2 s 340142 163200 340198 164400 6 la_iena[101]
port 71 nsew signal tristate
rlabel metal2 s 343546 163200 343602 164400 6 la_iena[102]
port 72 nsew signal tristate
rlabel metal2 s 346858 163200 346914 164400 6 la_iena[103]
port 73 nsew signal tristate
rlabel metal2 s 350262 163200 350318 164400 6 la_iena[104]
port 74 nsew signal tristate
rlabel metal2 s 353666 163200 353722 164400 6 la_iena[105]
port 75 nsew signal tristate
rlabel metal2 s 356978 163200 357034 164400 6 la_iena[106]
port 76 nsew signal tristate
rlabel metal2 s 360382 163200 360438 164400 6 la_iena[107]
port 77 nsew signal tristate
rlabel metal2 s 363694 163200 363750 164400 6 la_iena[108]
port 78 nsew signal tristate
rlabel metal2 s 367098 163200 367154 164400 6 la_iena[109]
port 79 nsew signal tristate
rlabel metal2 s 33966 163200 34022 164400 6 la_iena[10]
port 80 nsew signal tristate
rlabel metal2 s 370410 163200 370466 164400 6 la_iena[110]
port 81 nsew signal tristate
rlabel metal2 s 373814 163200 373870 164400 6 la_iena[111]
port 82 nsew signal tristate
rlabel metal2 s 377218 163200 377274 164400 6 la_iena[112]
port 83 nsew signal tristate
rlabel metal2 s 380530 163200 380586 164400 6 la_iena[113]
port 84 nsew signal tristate
rlabel metal2 s 383934 163200 383990 164400 6 la_iena[114]
port 85 nsew signal tristate
rlabel metal2 s 387246 163200 387302 164400 6 la_iena[115]
port 86 nsew signal tristate
rlabel metal2 s 390650 163200 390706 164400 6 la_iena[116]
port 87 nsew signal tristate
rlabel metal2 s 393962 163200 394018 164400 6 la_iena[117]
port 88 nsew signal tristate
rlabel metal2 s 397366 163200 397422 164400 6 la_iena[118]
port 89 nsew signal tristate
rlabel metal2 s 400770 163200 400826 164400 6 la_iena[119]
port 90 nsew signal tristate
rlabel metal2 s 37370 163200 37426 164400 6 la_iena[11]
port 91 nsew signal tristate
rlabel metal2 s 404082 163200 404138 164400 6 la_iena[120]
port 92 nsew signal tristate
rlabel metal2 s 407486 163200 407542 164400 6 la_iena[121]
port 93 nsew signal tristate
rlabel metal2 s 410798 163200 410854 164400 6 la_iena[122]
port 94 nsew signal tristate
rlabel metal2 s 414202 163200 414258 164400 6 la_iena[123]
port 95 nsew signal tristate
rlabel metal2 s 417514 163200 417570 164400 6 la_iena[124]
port 96 nsew signal tristate
rlabel metal2 s 420918 163200 420974 164400 6 la_iena[125]
port 97 nsew signal tristate
rlabel metal2 s 424322 163200 424378 164400 6 la_iena[126]
port 98 nsew signal tristate
rlabel metal2 s 427634 163200 427690 164400 6 la_iena[127]
port 99 nsew signal tristate
rlabel metal2 s 40682 163200 40738 164400 6 la_iena[12]
port 100 nsew signal tristate
rlabel metal2 s 44086 163200 44142 164400 6 la_iena[13]
port 101 nsew signal tristate
rlabel metal2 s 47490 163200 47546 164400 6 la_iena[14]
port 102 nsew signal tristate
rlabel metal2 s 50802 163200 50858 164400 6 la_iena[15]
port 103 nsew signal tristate
rlabel metal2 s 54206 163200 54262 164400 6 la_iena[16]
port 104 nsew signal tristate
rlabel metal2 s 57518 163200 57574 164400 6 la_iena[17]
port 105 nsew signal tristate
rlabel metal2 s 60922 163200 60978 164400 6 la_iena[18]
port 106 nsew signal tristate
rlabel metal2 s 64234 163200 64290 164400 6 la_iena[19]
port 107 nsew signal tristate
rlabel metal2 s 3698 163200 3754 164400 6 la_iena[1]
port 108 nsew signal tristate
rlabel metal2 s 67638 163200 67694 164400 6 la_iena[20]
port 109 nsew signal tristate
rlabel metal2 s 71042 163200 71098 164400 6 la_iena[21]
port 110 nsew signal tristate
rlabel metal2 s 74354 163200 74410 164400 6 la_iena[22]
port 111 nsew signal tristate
rlabel metal2 s 77758 163200 77814 164400 6 la_iena[23]
port 112 nsew signal tristate
rlabel metal2 s 81070 163200 81126 164400 6 la_iena[24]
port 113 nsew signal tristate
rlabel metal2 s 84474 163200 84530 164400 6 la_iena[25]
port 114 nsew signal tristate
rlabel metal2 s 87786 163200 87842 164400 6 la_iena[26]
port 115 nsew signal tristate
rlabel metal2 s 91190 163200 91246 164400 6 la_iena[27]
port 116 nsew signal tristate
rlabel metal2 s 94594 163200 94650 164400 6 la_iena[28]
port 117 nsew signal tristate
rlabel metal2 s 97906 163200 97962 164400 6 la_iena[29]
port 118 nsew signal tristate
rlabel metal2 s 7102 163200 7158 164400 6 la_iena[2]
port 119 nsew signal tristate
rlabel metal2 s 101310 163200 101366 164400 6 la_iena[30]
port 120 nsew signal tristate
rlabel metal2 s 104622 163200 104678 164400 6 la_iena[31]
port 121 nsew signal tristate
rlabel metal2 s 108026 163200 108082 164400 6 la_iena[32]
port 122 nsew signal tristate
rlabel metal2 s 111338 163200 111394 164400 6 la_iena[33]
port 123 nsew signal tristate
rlabel metal2 s 114742 163200 114798 164400 6 la_iena[34]
port 124 nsew signal tristate
rlabel metal2 s 118146 163200 118202 164400 6 la_iena[35]
port 125 nsew signal tristate
rlabel metal2 s 121458 163200 121514 164400 6 la_iena[36]
port 126 nsew signal tristate
rlabel metal2 s 124862 163200 124918 164400 6 la_iena[37]
port 127 nsew signal tristate
rlabel metal2 s 128174 163200 128230 164400 6 la_iena[38]
port 128 nsew signal tristate
rlabel metal2 s 131578 163200 131634 164400 6 la_iena[39]
port 129 nsew signal tristate
rlabel metal2 s 10414 163200 10470 164400 6 la_iena[3]
port 130 nsew signal tristate
rlabel metal2 s 134890 163200 134946 164400 6 la_iena[40]
port 131 nsew signal tristate
rlabel metal2 s 138294 163200 138350 164400 6 la_iena[41]
port 132 nsew signal tristate
rlabel metal2 s 141698 163200 141754 164400 6 la_iena[42]
port 133 nsew signal tristate
rlabel metal2 s 145010 163200 145066 164400 6 la_iena[43]
port 134 nsew signal tristate
rlabel metal2 s 148414 163200 148470 164400 6 la_iena[44]
port 135 nsew signal tristate
rlabel metal2 s 151726 163200 151782 164400 6 la_iena[45]
port 136 nsew signal tristate
rlabel metal2 s 155130 163200 155186 164400 6 la_iena[46]
port 137 nsew signal tristate
rlabel metal2 s 158442 163200 158498 164400 6 la_iena[47]
port 138 nsew signal tristate
rlabel metal2 s 161846 163200 161902 164400 6 la_iena[48]
port 139 nsew signal tristate
rlabel metal2 s 165250 163200 165306 164400 6 la_iena[49]
port 140 nsew signal tristate
rlabel metal2 s 13818 163200 13874 164400 6 la_iena[4]
port 141 nsew signal tristate
rlabel metal2 s 168562 163200 168618 164400 6 la_iena[50]
port 142 nsew signal tristate
rlabel metal2 s 171966 163200 172022 164400 6 la_iena[51]
port 143 nsew signal tristate
rlabel metal2 s 175278 163200 175334 164400 6 la_iena[52]
port 144 nsew signal tristate
rlabel metal2 s 178682 163200 178738 164400 6 la_iena[53]
port 145 nsew signal tristate
rlabel metal2 s 181994 163200 182050 164400 6 la_iena[54]
port 146 nsew signal tristate
rlabel metal2 s 185398 163200 185454 164400 6 la_iena[55]
port 147 nsew signal tristate
rlabel metal2 s 188802 163200 188858 164400 6 la_iena[56]
port 148 nsew signal tristate
rlabel metal2 s 192114 163200 192170 164400 6 la_iena[57]
port 149 nsew signal tristate
rlabel metal2 s 195518 163200 195574 164400 6 la_iena[58]
port 150 nsew signal tristate
rlabel metal2 s 198830 163200 198886 164400 6 la_iena[59]
port 151 nsew signal tristate
rlabel metal2 s 17130 163200 17186 164400 6 la_iena[5]
port 152 nsew signal tristate
rlabel metal2 s 202234 163200 202290 164400 6 la_iena[60]
port 153 nsew signal tristate
rlabel metal2 s 205546 163200 205602 164400 6 la_iena[61]
port 154 nsew signal tristate
rlabel metal2 s 208950 163200 209006 164400 6 la_iena[62]
port 155 nsew signal tristate
rlabel metal2 s 212354 163200 212410 164400 6 la_iena[63]
port 156 nsew signal tristate
rlabel metal2 s 215666 163200 215722 164400 6 la_iena[64]
port 157 nsew signal tristate
rlabel metal2 s 219070 163200 219126 164400 6 la_iena[65]
port 158 nsew signal tristate
rlabel metal2 s 222382 163200 222438 164400 6 la_iena[66]
port 159 nsew signal tristate
rlabel metal2 s 225786 163200 225842 164400 6 la_iena[67]
port 160 nsew signal tristate
rlabel metal2 s 229098 163200 229154 164400 6 la_iena[68]
port 161 nsew signal tristate
rlabel metal2 s 232502 163200 232558 164400 6 la_iena[69]
port 162 nsew signal tristate
rlabel metal2 s 20534 163200 20590 164400 6 la_iena[6]
port 163 nsew signal tristate
rlabel metal2 s 235906 163200 235962 164400 6 la_iena[70]
port 164 nsew signal tristate
rlabel metal2 s 239218 163200 239274 164400 6 la_iena[71]
port 165 nsew signal tristate
rlabel metal2 s 242622 163200 242678 164400 6 la_iena[72]
port 166 nsew signal tristate
rlabel metal2 s 245934 163200 245990 164400 6 la_iena[73]
port 167 nsew signal tristate
rlabel metal2 s 249338 163200 249394 164400 6 la_iena[74]
port 168 nsew signal tristate
rlabel metal2 s 252650 163200 252706 164400 6 la_iena[75]
port 169 nsew signal tristate
rlabel metal2 s 256054 163200 256110 164400 6 la_iena[76]
port 170 nsew signal tristate
rlabel metal2 s 259458 163200 259514 164400 6 la_iena[77]
port 171 nsew signal tristate
rlabel metal2 s 262770 163200 262826 164400 6 la_iena[78]
port 172 nsew signal tristate
rlabel metal2 s 266174 163200 266230 164400 6 la_iena[79]
port 173 nsew signal tristate
rlabel metal2 s 23938 163200 23994 164400 6 la_iena[7]
port 174 nsew signal tristate
rlabel metal2 s 269486 163200 269542 164400 6 la_iena[80]
port 175 nsew signal tristate
rlabel metal2 s 272890 163200 272946 164400 6 la_iena[81]
port 176 nsew signal tristate
rlabel metal2 s 276202 163200 276258 164400 6 la_iena[82]
port 177 nsew signal tristate
rlabel metal2 s 279606 163200 279662 164400 6 la_iena[83]
port 178 nsew signal tristate
rlabel metal2 s 283010 163200 283066 164400 6 la_iena[84]
port 179 nsew signal tristate
rlabel metal2 s 286322 163200 286378 164400 6 la_iena[85]
port 180 nsew signal tristate
rlabel metal2 s 289726 163200 289782 164400 6 la_iena[86]
port 181 nsew signal tristate
rlabel metal2 s 293038 163200 293094 164400 6 la_iena[87]
port 182 nsew signal tristate
rlabel metal2 s 296442 163200 296498 164400 6 la_iena[88]
port 183 nsew signal tristate
rlabel metal2 s 299754 163200 299810 164400 6 la_iena[89]
port 184 nsew signal tristate
rlabel metal2 s 27250 163200 27306 164400 6 la_iena[8]
port 185 nsew signal tristate
rlabel metal2 s 303158 163200 303214 164400 6 la_iena[90]
port 186 nsew signal tristate
rlabel metal2 s 306562 163200 306618 164400 6 la_iena[91]
port 187 nsew signal tristate
rlabel metal2 s 309874 163200 309930 164400 6 la_iena[92]
port 188 nsew signal tristate
rlabel metal2 s 313278 163200 313334 164400 6 la_iena[93]
port 189 nsew signal tristate
rlabel metal2 s 316590 163200 316646 164400 6 la_iena[94]
port 190 nsew signal tristate
rlabel metal2 s 319994 163200 320050 164400 6 la_iena[95]
port 191 nsew signal tristate
rlabel metal2 s 323306 163200 323362 164400 6 la_iena[96]
port 192 nsew signal tristate
rlabel metal2 s 326710 163200 326766 164400 6 la_iena[97]
port 193 nsew signal tristate
rlabel metal2 s 330114 163200 330170 164400 6 la_iena[98]
port 194 nsew signal tristate
rlabel metal2 s 333426 163200 333482 164400 6 la_iena[99]
port 195 nsew signal tristate
rlabel metal2 s 30654 163200 30710 164400 6 la_iena[9]
port 196 nsew signal tristate
rlabel metal2 s 1214 163200 1270 164400 6 la_input[0]
port 197 nsew signal input
rlabel metal2 s 337658 163200 337714 164400 6 la_input[100]
port 198 nsew signal input
rlabel metal2 s 340970 163200 341026 164400 6 la_input[101]
port 199 nsew signal input
rlabel metal2 s 344374 163200 344430 164400 6 la_input[102]
port 200 nsew signal input
rlabel metal2 s 347778 163200 347834 164400 6 la_input[103]
port 201 nsew signal input
rlabel metal2 s 351090 163200 351146 164400 6 la_input[104]
port 202 nsew signal input
rlabel metal2 s 354494 163200 354550 164400 6 la_input[105]
port 203 nsew signal input
rlabel metal2 s 357806 163200 357862 164400 6 la_input[106]
port 204 nsew signal input
rlabel metal2 s 361210 163200 361266 164400 6 la_input[107]
port 205 nsew signal input
rlabel metal2 s 364522 163200 364578 164400 6 la_input[108]
port 206 nsew signal input
rlabel metal2 s 367926 163200 367982 164400 6 la_input[109]
port 207 nsew signal input
rlabel metal2 s 34794 163200 34850 164400 6 la_input[10]
port 208 nsew signal input
rlabel metal2 s 371330 163200 371386 164400 6 la_input[110]
port 209 nsew signal input
rlabel metal2 s 374642 163200 374698 164400 6 la_input[111]
port 210 nsew signal input
rlabel metal2 s 378046 163200 378102 164400 6 la_input[112]
port 211 nsew signal input
rlabel metal2 s 381358 163200 381414 164400 6 la_input[113]
port 212 nsew signal input
rlabel metal2 s 384762 163200 384818 164400 6 la_input[114]
port 213 nsew signal input
rlabel metal2 s 388074 163200 388130 164400 6 la_input[115]
port 214 nsew signal input
rlabel metal2 s 391478 163200 391534 164400 6 la_input[116]
port 215 nsew signal input
rlabel metal2 s 394882 163200 394938 164400 6 la_input[117]
port 216 nsew signal input
rlabel metal2 s 398194 163200 398250 164400 6 la_input[118]
port 217 nsew signal input
rlabel metal2 s 401598 163200 401654 164400 6 la_input[119]
port 218 nsew signal input
rlabel metal2 s 38198 163200 38254 164400 6 la_input[11]
port 219 nsew signal input
rlabel metal2 s 404910 163200 404966 164400 6 la_input[120]
port 220 nsew signal input
rlabel metal2 s 408314 163200 408370 164400 6 la_input[121]
port 221 nsew signal input
rlabel metal2 s 411626 163200 411682 164400 6 la_input[122]
port 222 nsew signal input
rlabel metal2 s 415030 163200 415086 164400 6 la_input[123]
port 223 nsew signal input
rlabel metal2 s 418434 163200 418490 164400 6 la_input[124]
port 224 nsew signal input
rlabel metal2 s 421746 163200 421802 164400 6 la_input[125]
port 225 nsew signal input
rlabel metal2 s 425150 163200 425206 164400 6 la_input[126]
port 226 nsew signal input
rlabel metal2 s 428462 163200 428518 164400 6 la_input[127]
port 227 nsew signal input
rlabel metal2 s 41602 163200 41658 164400 6 la_input[12]
port 228 nsew signal input
rlabel metal2 s 44914 163200 44970 164400 6 la_input[13]
port 229 nsew signal input
rlabel metal2 s 48318 163200 48374 164400 6 la_input[14]
port 230 nsew signal input
rlabel metal2 s 51630 163200 51686 164400 6 la_input[15]
port 231 nsew signal input
rlabel metal2 s 55034 163200 55090 164400 6 la_input[16]
port 232 nsew signal input
rlabel metal2 s 58346 163200 58402 164400 6 la_input[17]
port 233 nsew signal input
rlabel metal2 s 61750 163200 61806 164400 6 la_input[18]
port 234 nsew signal input
rlabel metal2 s 65154 163200 65210 164400 6 la_input[19]
port 235 nsew signal input
rlabel metal2 s 4526 163200 4582 164400 6 la_input[1]
port 236 nsew signal input
rlabel metal2 s 68466 163200 68522 164400 6 la_input[20]
port 237 nsew signal input
rlabel metal2 s 71870 163200 71926 164400 6 la_input[21]
port 238 nsew signal input
rlabel metal2 s 75182 163200 75238 164400 6 la_input[22]
port 239 nsew signal input
rlabel metal2 s 78586 163200 78642 164400 6 la_input[23]
port 240 nsew signal input
rlabel metal2 s 81898 163200 81954 164400 6 la_input[24]
port 241 nsew signal input
rlabel metal2 s 85302 163200 85358 164400 6 la_input[25]
port 242 nsew signal input
rlabel metal2 s 88706 163200 88762 164400 6 la_input[26]
port 243 nsew signal input
rlabel metal2 s 92018 163200 92074 164400 6 la_input[27]
port 244 nsew signal input
rlabel metal2 s 95422 163200 95478 164400 6 la_input[28]
port 245 nsew signal input
rlabel metal2 s 98734 163200 98790 164400 6 la_input[29]
port 246 nsew signal input
rlabel metal2 s 7930 163200 7986 164400 6 la_input[2]
port 247 nsew signal input
rlabel metal2 s 102138 163200 102194 164400 6 la_input[30]
port 248 nsew signal input
rlabel metal2 s 105450 163200 105506 164400 6 la_input[31]
port 249 nsew signal input
rlabel metal2 s 108854 163200 108910 164400 6 la_input[32]
port 250 nsew signal input
rlabel metal2 s 112258 163200 112314 164400 6 la_input[33]
port 251 nsew signal input
rlabel metal2 s 115570 163200 115626 164400 6 la_input[34]
port 252 nsew signal input
rlabel metal2 s 118974 163200 119030 164400 6 la_input[35]
port 253 nsew signal input
rlabel metal2 s 122286 163200 122342 164400 6 la_input[36]
port 254 nsew signal input
rlabel metal2 s 125690 163200 125746 164400 6 la_input[37]
port 255 nsew signal input
rlabel metal2 s 129002 163200 129058 164400 6 la_input[38]
port 256 nsew signal input
rlabel metal2 s 132406 163200 132462 164400 6 la_input[39]
port 257 nsew signal input
rlabel metal2 s 11242 163200 11298 164400 6 la_input[3]
port 258 nsew signal input
rlabel metal2 s 135810 163200 135866 164400 6 la_input[40]
port 259 nsew signal input
rlabel metal2 s 139122 163200 139178 164400 6 la_input[41]
port 260 nsew signal input
rlabel metal2 s 142526 163200 142582 164400 6 la_input[42]
port 261 nsew signal input
rlabel metal2 s 145838 163200 145894 164400 6 la_input[43]
port 262 nsew signal input
rlabel metal2 s 149242 163200 149298 164400 6 la_input[44]
port 263 nsew signal input
rlabel metal2 s 152554 163200 152610 164400 6 la_input[45]
port 264 nsew signal input
rlabel metal2 s 155958 163200 156014 164400 6 la_input[46]
port 265 nsew signal input
rlabel metal2 s 159362 163200 159418 164400 6 la_input[47]
port 266 nsew signal input
rlabel metal2 s 162674 163200 162730 164400 6 la_input[48]
port 267 nsew signal input
rlabel metal2 s 166078 163200 166134 164400 6 la_input[49]
port 268 nsew signal input
rlabel metal2 s 14646 163200 14702 164400 6 la_input[4]
port 269 nsew signal input
rlabel metal2 s 169390 163200 169446 164400 6 la_input[50]
port 270 nsew signal input
rlabel metal2 s 172794 163200 172850 164400 6 la_input[51]
port 271 nsew signal input
rlabel metal2 s 176106 163200 176162 164400 6 la_input[52]
port 272 nsew signal input
rlabel metal2 s 179510 163200 179566 164400 6 la_input[53]
port 273 nsew signal input
rlabel metal2 s 182914 163200 182970 164400 6 la_input[54]
port 274 nsew signal input
rlabel metal2 s 186226 163200 186282 164400 6 la_input[55]
port 275 nsew signal input
rlabel metal2 s 189630 163200 189686 164400 6 la_input[56]
port 276 nsew signal input
rlabel metal2 s 192942 163200 192998 164400 6 la_input[57]
port 277 nsew signal input
rlabel metal2 s 196346 163200 196402 164400 6 la_input[58]
port 278 nsew signal input
rlabel metal2 s 199658 163200 199714 164400 6 la_input[59]
port 279 nsew signal input
rlabel metal2 s 18050 163200 18106 164400 6 la_input[5]
port 280 nsew signal input
rlabel metal2 s 203062 163200 203118 164400 6 la_input[60]
port 281 nsew signal input
rlabel metal2 s 206466 163200 206522 164400 6 la_input[61]
port 282 nsew signal input
rlabel metal2 s 209778 163200 209834 164400 6 la_input[62]
port 283 nsew signal input
rlabel metal2 s 213182 163200 213238 164400 6 la_input[63]
port 284 nsew signal input
rlabel metal2 s 216494 163200 216550 164400 6 la_input[64]
port 285 nsew signal input
rlabel metal2 s 219898 163200 219954 164400 6 la_input[65]
port 286 nsew signal input
rlabel metal2 s 223210 163200 223266 164400 6 la_input[66]
port 287 nsew signal input
rlabel metal2 s 226614 163200 226670 164400 6 la_input[67]
port 288 nsew signal input
rlabel metal2 s 230018 163200 230074 164400 6 la_input[68]
port 289 nsew signal input
rlabel metal2 s 233330 163200 233386 164400 6 la_input[69]
port 290 nsew signal input
rlabel metal2 s 21362 163200 21418 164400 6 la_input[6]
port 291 nsew signal input
rlabel metal2 s 236734 163200 236790 164400 6 la_input[70]
port 292 nsew signal input
rlabel metal2 s 240046 163200 240102 164400 6 la_input[71]
port 293 nsew signal input
rlabel metal2 s 243450 163200 243506 164400 6 la_input[72]
port 294 nsew signal input
rlabel metal2 s 246762 163200 246818 164400 6 la_input[73]
port 295 nsew signal input
rlabel metal2 s 250166 163200 250222 164400 6 la_input[74]
port 296 nsew signal input
rlabel metal2 s 253570 163200 253626 164400 6 la_input[75]
port 297 nsew signal input
rlabel metal2 s 256882 163200 256938 164400 6 la_input[76]
port 298 nsew signal input
rlabel metal2 s 260286 163200 260342 164400 6 la_input[77]
port 299 nsew signal input
rlabel metal2 s 263598 163200 263654 164400 6 la_input[78]
port 300 nsew signal input
rlabel metal2 s 267002 163200 267058 164400 6 la_input[79]
port 301 nsew signal input
rlabel metal2 s 24766 163200 24822 164400 6 la_input[7]
port 302 nsew signal input
rlabel metal2 s 270314 163200 270370 164400 6 la_input[80]
port 303 nsew signal input
rlabel metal2 s 273718 163200 273774 164400 6 la_input[81]
port 304 nsew signal input
rlabel metal2 s 277122 163200 277178 164400 6 la_input[82]
port 305 nsew signal input
rlabel metal2 s 280434 163200 280490 164400 6 la_input[83]
port 306 nsew signal input
rlabel metal2 s 283838 163200 283894 164400 6 la_input[84]
port 307 nsew signal input
rlabel metal2 s 287150 163200 287206 164400 6 la_input[85]
port 308 nsew signal input
rlabel metal2 s 290554 163200 290610 164400 6 la_input[86]
port 309 nsew signal input
rlabel metal2 s 293866 163200 293922 164400 6 la_input[87]
port 310 nsew signal input
rlabel metal2 s 297270 163200 297326 164400 6 la_input[88]
port 311 nsew signal input
rlabel metal2 s 300674 163200 300730 164400 6 la_input[89]
port 312 nsew signal input
rlabel metal2 s 28078 163200 28134 164400 6 la_input[8]
port 313 nsew signal input
rlabel metal2 s 303986 163200 304042 164400 6 la_input[90]
port 314 nsew signal input
rlabel metal2 s 307390 163200 307446 164400 6 la_input[91]
port 315 nsew signal input
rlabel metal2 s 310702 163200 310758 164400 6 la_input[92]
port 316 nsew signal input
rlabel metal2 s 314106 163200 314162 164400 6 la_input[93]
port 317 nsew signal input
rlabel metal2 s 317418 163200 317474 164400 6 la_input[94]
port 318 nsew signal input
rlabel metal2 s 320822 163200 320878 164400 6 la_input[95]
port 319 nsew signal input
rlabel metal2 s 324226 163200 324282 164400 6 la_input[96]
port 320 nsew signal input
rlabel metal2 s 327538 163200 327594 164400 6 la_input[97]
port 321 nsew signal input
rlabel metal2 s 330942 163200 330998 164400 6 la_input[98]
port 322 nsew signal input
rlabel metal2 s 334254 163200 334310 164400 6 la_input[99]
port 323 nsew signal input
rlabel metal2 s 31482 163200 31538 164400 6 la_input[9]
port 324 nsew signal input
rlabel metal2 s 2042 163200 2098 164400 6 la_oenb[0]
port 325 nsew signal tristate
rlabel metal2 s 338486 163200 338542 164400 6 la_oenb[100]
port 326 nsew signal tristate
rlabel metal2 s 341890 163200 341946 164400 6 la_oenb[101]
port 327 nsew signal tristate
rlabel metal2 s 345202 163200 345258 164400 6 la_oenb[102]
port 328 nsew signal tristate
rlabel metal2 s 348606 163200 348662 164400 6 la_oenb[103]
port 329 nsew signal tristate
rlabel metal2 s 351918 163200 351974 164400 6 la_oenb[104]
port 330 nsew signal tristate
rlabel metal2 s 355322 163200 355378 164400 6 la_oenb[105]
port 331 nsew signal tristate
rlabel metal2 s 358634 163200 358690 164400 6 la_oenb[106]
port 332 nsew signal tristate
rlabel metal2 s 362038 163200 362094 164400 6 la_oenb[107]
port 333 nsew signal tristate
rlabel metal2 s 365442 163200 365498 164400 6 la_oenb[108]
port 334 nsew signal tristate
rlabel metal2 s 368754 163200 368810 164400 6 la_oenb[109]
port 335 nsew signal tristate
rlabel metal2 s 35714 163200 35770 164400 6 la_oenb[10]
port 336 nsew signal tristate
rlabel metal2 s 372158 163200 372214 164400 6 la_oenb[110]
port 337 nsew signal tristate
rlabel metal2 s 375470 163200 375526 164400 6 la_oenb[111]
port 338 nsew signal tristate
rlabel metal2 s 378874 163200 378930 164400 6 la_oenb[112]
port 339 nsew signal tristate
rlabel metal2 s 382186 163200 382242 164400 6 la_oenb[113]
port 340 nsew signal tristate
rlabel metal2 s 385590 163200 385646 164400 6 la_oenb[114]
port 341 nsew signal tristate
rlabel metal2 s 388994 163200 389050 164400 6 la_oenb[115]
port 342 nsew signal tristate
rlabel metal2 s 392306 163200 392362 164400 6 la_oenb[116]
port 343 nsew signal tristate
rlabel metal2 s 395710 163200 395766 164400 6 la_oenb[117]
port 344 nsew signal tristate
rlabel metal2 s 399022 163200 399078 164400 6 la_oenb[118]
port 345 nsew signal tristate
rlabel metal2 s 402426 163200 402482 164400 6 la_oenb[119]
port 346 nsew signal tristate
rlabel metal2 s 39026 163200 39082 164400 6 la_oenb[11]
port 347 nsew signal tristate
rlabel metal2 s 405738 163200 405794 164400 6 la_oenb[120]
port 348 nsew signal tristate
rlabel metal2 s 409142 163200 409198 164400 6 la_oenb[121]
port 349 nsew signal tristate
rlabel metal2 s 412546 163200 412602 164400 6 la_oenb[122]
port 350 nsew signal tristate
rlabel metal2 s 415858 163200 415914 164400 6 la_oenb[123]
port 351 nsew signal tristate
rlabel metal2 s 419262 163200 419318 164400 6 la_oenb[124]
port 352 nsew signal tristate
rlabel metal2 s 422574 163200 422630 164400 6 la_oenb[125]
port 353 nsew signal tristate
rlabel metal2 s 425978 163200 426034 164400 6 la_oenb[126]
port 354 nsew signal tristate
rlabel metal2 s 429290 163200 429346 164400 6 la_oenb[127]
port 355 nsew signal tristate
rlabel metal2 s 42430 163200 42486 164400 6 la_oenb[12]
port 356 nsew signal tristate
rlabel metal2 s 45742 163200 45798 164400 6 la_oenb[13]
port 357 nsew signal tristate
rlabel metal2 s 49146 163200 49202 164400 6 la_oenb[14]
port 358 nsew signal tristate
rlabel metal2 s 52458 163200 52514 164400 6 la_oenb[15]
port 359 nsew signal tristate
rlabel metal2 s 55862 163200 55918 164400 6 la_oenb[16]
port 360 nsew signal tristate
rlabel metal2 s 59266 163200 59322 164400 6 la_oenb[17]
port 361 nsew signal tristate
rlabel metal2 s 62578 163200 62634 164400 6 la_oenb[18]
port 362 nsew signal tristate
rlabel metal2 s 65982 163200 66038 164400 6 la_oenb[19]
port 363 nsew signal tristate
rlabel metal2 s 5354 163200 5410 164400 6 la_oenb[1]
port 364 nsew signal tristate
rlabel metal2 s 69294 163200 69350 164400 6 la_oenb[20]
port 365 nsew signal tristate
rlabel metal2 s 72698 163200 72754 164400 6 la_oenb[21]
port 366 nsew signal tristate
rlabel metal2 s 76010 163200 76066 164400 6 la_oenb[22]
port 367 nsew signal tristate
rlabel metal2 s 79414 163200 79470 164400 6 la_oenb[23]
port 368 nsew signal tristate
rlabel metal2 s 82818 163200 82874 164400 6 la_oenb[24]
port 369 nsew signal tristate
rlabel metal2 s 86130 163200 86186 164400 6 la_oenb[25]
port 370 nsew signal tristate
rlabel metal2 s 89534 163200 89590 164400 6 la_oenb[26]
port 371 nsew signal tristate
rlabel metal2 s 92846 163200 92902 164400 6 la_oenb[27]
port 372 nsew signal tristate
rlabel metal2 s 96250 163200 96306 164400 6 la_oenb[28]
port 373 nsew signal tristate
rlabel metal2 s 99562 163200 99618 164400 6 la_oenb[29]
port 374 nsew signal tristate
rlabel metal2 s 8758 163200 8814 164400 6 la_oenb[2]
port 375 nsew signal tristate
rlabel metal2 s 102966 163200 103022 164400 6 la_oenb[30]
port 376 nsew signal tristate
rlabel metal2 s 106370 163200 106426 164400 6 la_oenb[31]
port 377 nsew signal tristate
rlabel metal2 s 109682 163200 109738 164400 6 la_oenb[32]
port 378 nsew signal tristate
rlabel metal2 s 113086 163200 113142 164400 6 la_oenb[33]
port 379 nsew signal tristate
rlabel metal2 s 116398 163200 116454 164400 6 la_oenb[34]
port 380 nsew signal tristate
rlabel metal2 s 119802 163200 119858 164400 6 la_oenb[35]
port 381 nsew signal tristate
rlabel metal2 s 123114 163200 123170 164400 6 la_oenb[36]
port 382 nsew signal tristate
rlabel metal2 s 126518 163200 126574 164400 6 la_oenb[37]
port 383 nsew signal tristate
rlabel metal2 s 129922 163200 129978 164400 6 la_oenb[38]
port 384 nsew signal tristate
rlabel metal2 s 133234 163200 133290 164400 6 la_oenb[39]
port 385 nsew signal tristate
rlabel metal2 s 12162 163200 12218 164400 6 la_oenb[3]
port 386 nsew signal tristate
rlabel metal2 s 136638 163200 136694 164400 6 la_oenb[40]
port 387 nsew signal tristate
rlabel metal2 s 139950 163200 140006 164400 6 la_oenb[41]
port 388 nsew signal tristate
rlabel metal2 s 143354 163200 143410 164400 6 la_oenb[42]
port 389 nsew signal tristate
rlabel metal2 s 146666 163200 146722 164400 6 la_oenb[43]
port 390 nsew signal tristate
rlabel metal2 s 150070 163200 150126 164400 6 la_oenb[44]
port 391 nsew signal tristate
rlabel metal2 s 153474 163200 153530 164400 6 la_oenb[45]
port 392 nsew signal tristate
rlabel metal2 s 156786 163200 156842 164400 6 la_oenb[46]
port 393 nsew signal tristate
rlabel metal2 s 160190 163200 160246 164400 6 la_oenb[47]
port 394 nsew signal tristate
rlabel metal2 s 163502 163200 163558 164400 6 la_oenb[48]
port 395 nsew signal tristate
rlabel metal2 s 166906 163200 166962 164400 6 la_oenb[49]
port 396 nsew signal tristate
rlabel metal2 s 15474 163200 15530 164400 6 la_oenb[4]
port 397 nsew signal tristate
rlabel metal2 s 170218 163200 170274 164400 6 la_oenb[50]
port 398 nsew signal tristate
rlabel metal2 s 173622 163200 173678 164400 6 la_oenb[51]
port 399 nsew signal tristate
rlabel metal2 s 177026 163200 177082 164400 6 la_oenb[52]
port 400 nsew signal tristate
rlabel metal2 s 180338 163200 180394 164400 6 la_oenb[53]
port 401 nsew signal tristate
rlabel metal2 s 183742 163200 183798 164400 6 la_oenb[54]
port 402 nsew signal tristate
rlabel metal2 s 187054 163200 187110 164400 6 la_oenb[55]
port 403 nsew signal tristate
rlabel metal2 s 190458 163200 190514 164400 6 la_oenb[56]
port 404 nsew signal tristate
rlabel metal2 s 193770 163200 193826 164400 6 la_oenb[57]
port 405 nsew signal tristate
rlabel metal2 s 197174 163200 197230 164400 6 la_oenb[58]
port 406 nsew signal tristate
rlabel metal2 s 200578 163200 200634 164400 6 la_oenb[59]
port 407 nsew signal tristate
rlabel metal2 s 18878 163200 18934 164400 6 la_oenb[5]
port 408 nsew signal tristate
rlabel metal2 s 203890 163200 203946 164400 6 la_oenb[60]
port 409 nsew signal tristate
rlabel metal2 s 207294 163200 207350 164400 6 la_oenb[61]
port 410 nsew signal tristate
rlabel metal2 s 210606 163200 210662 164400 6 la_oenb[62]
port 411 nsew signal tristate
rlabel metal2 s 214010 163200 214066 164400 6 la_oenb[63]
port 412 nsew signal tristate
rlabel metal2 s 217322 163200 217378 164400 6 la_oenb[64]
port 413 nsew signal tristate
rlabel metal2 s 220726 163200 220782 164400 6 la_oenb[65]
port 414 nsew signal tristate
rlabel metal2 s 224130 163200 224186 164400 6 la_oenb[66]
port 415 nsew signal tristate
rlabel metal2 s 227442 163200 227498 164400 6 la_oenb[67]
port 416 nsew signal tristate
rlabel metal2 s 230846 163200 230902 164400 6 la_oenb[68]
port 417 nsew signal tristate
rlabel metal2 s 234158 163200 234214 164400 6 la_oenb[69]
port 418 nsew signal tristate
rlabel metal2 s 22190 163200 22246 164400 6 la_oenb[6]
port 419 nsew signal tristate
rlabel metal2 s 237562 163200 237618 164400 6 la_oenb[70]
port 420 nsew signal tristate
rlabel metal2 s 240874 163200 240930 164400 6 la_oenb[71]
port 421 nsew signal tristate
rlabel metal2 s 244278 163200 244334 164400 6 la_oenb[72]
port 422 nsew signal tristate
rlabel metal2 s 247682 163200 247738 164400 6 la_oenb[73]
port 423 nsew signal tristate
rlabel metal2 s 250994 163200 251050 164400 6 la_oenb[74]
port 424 nsew signal tristate
rlabel metal2 s 254398 163200 254454 164400 6 la_oenb[75]
port 425 nsew signal tristate
rlabel metal2 s 257710 163200 257766 164400 6 la_oenb[76]
port 426 nsew signal tristate
rlabel metal2 s 261114 163200 261170 164400 6 la_oenb[77]
port 427 nsew signal tristate
rlabel metal2 s 264426 163200 264482 164400 6 la_oenb[78]
port 428 nsew signal tristate
rlabel metal2 s 267830 163200 267886 164400 6 la_oenb[79]
port 429 nsew signal tristate
rlabel metal2 s 25594 163200 25650 164400 6 la_oenb[7]
port 430 nsew signal tristate
rlabel metal2 s 271234 163200 271290 164400 6 la_oenb[80]
port 431 nsew signal tristate
rlabel metal2 s 274546 163200 274602 164400 6 la_oenb[81]
port 432 nsew signal tristate
rlabel metal2 s 277950 163200 278006 164400 6 la_oenb[82]
port 433 nsew signal tristate
rlabel metal2 s 281262 163200 281318 164400 6 la_oenb[83]
port 434 nsew signal tristate
rlabel metal2 s 284666 163200 284722 164400 6 la_oenb[84]
port 435 nsew signal tristate
rlabel metal2 s 287978 163200 288034 164400 6 la_oenb[85]
port 436 nsew signal tristate
rlabel metal2 s 291382 163200 291438 164400 6 la_oenb[86]
port 437 nsew signal tristate
rlabel metal2 s 294786 163200 294842 164400 6 la_oenb[87]
port 438 nsew signal tristate
rlabel metal2 s 298098 163200 298154 164400 6 la_oenb[88]
port 439 nsew signal tristate
rlabel metal2 s 301502 163200 301558 164400 6 la_oenb[89]
port 440 nsew signal tristate
rlabel metal2 s 28906 163200 28962 164400 6 la_oenb[8]
port 441 nsew signal tristate
rlabel metal2 s 304814 163200 304870 164400 6 la_oenb[90]
port 442 nsew signal tristate
rlabel metal2 s 308218 163200 308274 164400 6 la_oenb[91]
port 443 nsew signal tristate
rlabel metal2 s 311530 163200 311586 164400 6 la_oenb[92]
port 444 nsew signal tristate
rlabel metal2 s 314934 163200 314990 164400 6 la_oenb[93]
port 445 nsew signal tristate
rlabel metal2 s 318338 163200 318394 164400 6 la_oenb[94]
port 446 nsew signal tristate
rlabel metal2 s 321650 163200 321706 164400 6 la_oenb[95]
port 447 nsew signal tristate
rlabel metal2 s 325054 163200 325110 164400 6 la_oenb[96]
port 448 nsew signal tristate
rlabel metal2 s 328366 163200 328422 164400 6 la_oenb[97]
port 449 nsew signal tristate
rlabel metal2 s 331770 163200 331826 164400 6 la_oenb[98]
port 450 nsew signal tristate
rlabel metal2 s 335082 163200 335138 164400 6 la_oenb[99]
port 451 nsew signal tristate
rlabel metal2 s 32310 163200 32366 164400 6 la_oenb[9]
port 452 nsew signal tristate
rlabel metal2 s 2870 163200 2926 164400 6 la_output[0]
port 453 nsew signal tristate
rlabel metal2 s 339314 163200 339370 164400 6 la_output[100]
port 454 nsew signal tristate
rlabel metal2 s 342718 163200 342774 164400 6 la_output[101]
port 455 nsew signal tristate
rlabel metal2 s 346030 163200 346086 164400 6 la_output[102]
port 456 nsew signal tristate
rlabel metal2 s 349434 163200 349490 164400 6 la_output[103]
port 457 nsew signal tristate
rlabel metal2 s 352746 163200 352802 164400 6 la_output[104]
port 458 nsew signal tristate
rlabel metal2 s 356150 163200 356206 164400 6 la_output[105]
port 459 nsew signal tristate
rlabel metal2 s 359554 163200 359610 164400 6 la_output[106]
port 460 nsew signal tristate
rlabel metal2 s 362866 163200 362922 164400 6 la_output[107]
port 461 nsew signal tristate
rlabel metal2 s 366270 163200 366326 164400 6 la_output[108]
port 462 nsew signal tristate
rlabel metal2 s 369582 163200 369638 164400 6 la_output[109]
port 463 nsew signal tristate
rlabel metal2 s 36542 163200 36598 164400 6 la_output[10]
port 464 nsew signal tristate
rlabel metal2 s 372986 163200 373042 164400 6 la_output[110]
port 465 nsew signal tristate
rlabel metal2 s 376298 163200 376354 164400 6 la_output[111]
port 466 nsew signal tristate
rlabel metal2 s 379702 163200 379758 164400 6 la_output[112]
port 467 nsew signal tristate
rlabel metal2 s 383106 163200 383162 164400 6 la_output[113]
port 468 nsew signal tristate
rlabel metal2 s 386418 163200 386474 164400 6 la_output[114]
port 469 nsew signal tristate
rlabel metal2 s 389822 163200 389878 164400 6 la_output[115]
port 470 nsew signal tristate
rlabel metal2 s 393134 163200 393190 164400 6 la_output[116]
port 471 nsew signal tristate
rlabel metal2 s 396538 163200 396594 164400 6 la_output[117]
port 472 nsew signal tristate
rlabel metal2 s 399850 163200 399906 164400 6 la_output[118]
port 473 nsew signal tristate
rlabel metal2 s 403254 163200 403310 164400 6 la_output[119]
port 474 nsew signal tristate
rlabel metal2 s 39854 163200 39910 164400 6 la_output[11]
port 475 nsew signal tristate
rlabel metal2 s 406658 163200 406714 164400 6 la_output[120]
port 476 nsew signal tristate
rlabel metal2 s 409970 163200 410026 164400 6 la_output[121]
port 477 nsew signal tristate
rlabel metal2 s 413374 163200 413430 164400 6 la_output[122]
port 478 nsew signal tristate
rlabel metal2 s 416686 163200 416742 164400 6 la_output[123]
port 479 nsew signal tristate
rlabel metal2 s 420090 163200 420146 164400 6 la_output[124]
port 480 nsew signal tristate
rlabel metal2 s 423402 163200 423458 164400 6 la_output[125]
port 481 nsew signal tristate
rlabel metal2 s 426806 163200 426862 164400 6 la_output[126]
port 482 nsew signal tristate
rlabel metal2 s 430210 163200 430266 164400 6 la_output[127]
port 483 nsew signal tristate
rlabel metal2 s 43258 163200 43314 164400 6 la_output[12]
port 484 nsew signal tristate
rlabel metal2 s 46570 163200 46626 164400 6 la_output[13]
port 485 nsew signal tristate
rlabel metal2 s 49974 163200 50030 164400 6 la_output[14]
port 486 nsew signal tristate
rlabel metal2 s 53378 163200 53434 164400 6 la_output[15]
port 487 nsew signal tristate
rlabel metal2 s 56690 163200 56746 164400 6 la_output[16]
port 488 nsew signal tristate
rlabel metal2 s 60094 163200 60150 164400 6 la_output[17]
port 489 nsew signal tristate
rlabel metal2 s 63406 163200 63462 164400 6 la_output[18]
port 490 nsew signal tristate
rlabel metal2 s 66810 163200 66866 164400 6 la_output[19]
port 491 nsew signal tristate
rlabel metal2 s 6274 163200 6330 164400 6 la_output[1]
port 492 nsew signal tristate
rlabel metal2 s 70122 163200 70178 164400 6 la_output[20]
port 493 nsew signal tristate
rlabel metal2 s 73526 163200 73582 164400 6 la_output[21]
port 494 nsew signal tristate
rlabel metal2 s 76930 163200 76986 164400 6 la_output[22]
port 495 nsew signal tristate
rlabel metal2 s 80242 163200 80298 164400 6 la_output[23]
port 496 nsew signal tristate
rlabel metal2 s 83646 163200 83702 164400 6 la_output[24]
port 497 nsew signal tristate
rlabel metal2 s 86958 163200 87014 164400 6 la_output[25]
port 498 nsew signal tristate
rlabel metal2 s 90362 163200 90418 164400 6 la_output[26]
port 499 nsew signal tristate
rlabel metal2 s 93674 163200 93730 164400 6 la_output[27]
port 500 nsew signal tristate
rlabel metal2 s 97078 163200 97134 164400 6 la_output[28]
port 501 nsew signal tristate
rlabel metal2 s 100482 163200 100538 164400 6 la_output[29]
port 502 nsew signal tristate
rlabel metal2 s 9586 163200 9642 164400 6 la_output[2]
port 503 nsew signal tristate
rlabel metal2 s 103794 163200 103850 164400 6 la_output[30]
port 504 nsew signal tristate
rlabel metal2 s 107198 163200 107254 164400 6 la_output[31]
port 505 nsew signal tristate
rlabel metal2 s 110510 163200 110566 164400 6 la_output[32]
port 506 nsew signal tristate
rlabel metal2 s 113914 163200 113970 164400 6 la_output[33]
port 507 nsew signal tristate
rlabel metal2 s 117226 163200 117282 164400 6 la_output[34]
port 508 nsew signal tristate
rlabel metal2 s 120630 163200 120686 164400 6 la_output[35]
port 509 nsew signal tristate
rlabel metal2 s 124034 163200 124090 164400 6 la_output[36]
port 510 nsew signal tristate
rlabel metal2 s 127346 163200 127402 164400 6 la_output[37]
port 511 nsew signal tristate
rlabel metal2 s 130750 163200 130806 164400 6 la_output[38]
port 512 nsew signal tristate
rlabel metal2 s 134062 163200 134118 164400 6 la_output[39]
port 513 nsew signal tristate
rlabel metal2 s 12990 163200 13046 164400 6 la_output[3]
port 514 nsew signal tristate
rlabel metal2 s 137466 163200 137522 164400 6 la_output[40]
port 515 nsew signal tristate
rlabel metal2 s 140778 163200 140834 164400 6 la_output[41]
port 516 nsew signal tristate
rlabel metal2 s 144182 163200 144238 164400 6 la_output[42]
port 517 nsew signal tristate
rlabel metal2 s 147586 163200 147642 164400 6 la_output[43]
port 518 nsew signal tristate
rlabel metal2 s 150898 163200 150954 164400 6 la_output[44]
port 519 nsew signal tristate
rlabel metal2 s 154302 163200 154358 164400 6 la_output[45]
port 520 nsew signal tristate
rlabel metal2 s 157614 163200 157670 164400 6 la_output[46]
port 521 nsew signal tristate
rlabel metal2 s 161018 163200 161074 164400 6 la_output[47]
port 522 nsew signal tristate
rlabel metal2 s 164330 163200 164386 164400 6 la_output[48]
port 523 nsew signal tristate
rlabel metal2 s 167734 163200 167790 164400 6 la_output[49]
port 524 nsew signal tristate
rlabel metal2 s 16302 163200 16358 164400 6 la_output[4]
port 525 nsew signal tristate
rlabel metal2 s 171138 163200 171194 164400 6 la_output[50]
port 526 nsew signal tristate
rlabel metal2 s 174450 163200 174506 164400 6 la_output[51]
port 527 nsew signal tristate
rlabel metal2 s 177854 163200 177910 164400 6 la_output[52]
port 528 nsew signal tristate
rlabel metal2 s 181166 163200 181222 164400 6 la_output[53]
port 529 nsew signal tristate
rlabel metal2 s 184570 163200 184626 164400 6 la_output[54]
port 530 nsew signal tristate
rlabel metal2 s 187882 163200 187938 164400 6 la_output[55]
port 531 nsew signal tristate
rlabel metal2 s 191286 163200 191342 164400 6 la_output[56]
port 532 nsew signal tristate
rlabel metal2 s 194690 163200 194746 164400 6 la_output[57]
port 533 nsew signal tristate
rlabel metal2 s 198002 163200 198058 164400 6 la_output[58]
port 534 nsew signal tristate
rlabel metal2 s 201406 163200 201462 164400 6 la_output[59]
port 535 nsew signal tristate
rlabel metal2 s 19706 163200 19762 164400 6 la_output[5]
port 536 nsew signal tristate
rlabel metal2 s 204718 163200 204774 164400 6 la_output[60]
port 537 nsew signal tristate
rlabel metal2 s 208122 163200 208178 164400 6 la_output[61]
port 538 nsew signal tristate
rlabel metal2 s 211434 163200 211490 164400 6 la_output[62]
port 539 nsew signal tristate
rlabel metal2 s 214838 163200 214894 164400 6 la_output[63]
port 540 nsew signal tristate
rlabel metal2 s 218242 163200 218298 164400 6 la_output[64]
port 541 nsew signal tristate
rlabel metal2 s 221554 163200 221610 164400 6 la_output[65]
port 542 nsew signal tristate
rlabel metal2 s 224958 163200 225014 164400 6 la_output[66]
port 543 nsew signal tristate
rlabel metal2 s 228270 163200 228326 164400 6 la_output[67]
port 544 nsew signal tristate
rlabel metal2 s 231674 163200 231730 164400 6 la_output[68]
port 545 nsew signal tristate
rlabel metal2 s 234986 163200 235042 164400 6 la_output[69]
port 546 nsew signal tristate
rlabel metal2 s 23018 163200 23074 164400 6 la_output[6]
port 547 nsew signal tristate
rlabel metal2 s 238390 163200 238446 164400 6 la_output[70]
port 548 nsew signal tristate
rlabel metal2 s 241794 163200 241850 164400 6 la_output[71]
port 549 nsew signal tristate
rlabel metal2 s 245106 163200 245162 164400 6 la_output[72]
port 550 nsew signal tristate
rlabel metal2 s 248510 163200 248566 164400 6 la_output[73]
port 551 nsew signal tristate
rlabel metal2 s 251822 163200 251878 164400 6 la_output[74]
port 552 nsew signal tristate
rlabel metal2 s 255226 163200 255282 164400 6 la_output[75]
port 553 nsew signal tristate
rlabel metal2 s 258538 163200 258594 164400 6 la_output[76]
port 554 nsew signal tristate
rlabel metal2 s 261942 163200 261998 164400 6 la_output[77]
port 555 nsew signal tristate
rlabel metal2 s 265346 163200 265402 164400 6 la_output[78]
port 556 nsew signal tristate
rlabel metal2 s 268658 163200 268714 164400 6 la_output[79]
port 557 nsew signal tristate
rlabel metal2 s 26422 163200 26478 164400 6 la_output[7]
port 558 nsew signal tristate
rlabel metal2 s 272062 163200 272118 164400 6 la_output[80]
port 559 nsew signal tristate
rlabel metal2 s 275374 163200 275430 164400 6 la_output[81]
port 560 nsew signal tristate
rlabel metal2 s 278778 163200 278834 164400 6 la_output[82]
port 561 nsew signal tristate
rlabel metal2 s 282090 163200 282146 164400 6 la_output[83]
port 562 nsew signal tristate
rlabel metal2 s 285494 163200 285550 164400 6 la_output[84]
port 563 nsew signal tristate
rlabel metal2 s 288898 163200 288954 164400 6 la_output[85]
port 564 nsew signal tristate
rlabel metal2 s 292210 163200 292266 164400 6 la_output[86]
port 565 nsew signal tristate
rlabel metal2 s 295614 163200 295670 164400 6 la_output[87]
port 566 nsew signal tristate
rlabel metal2 s 298926 163200 298982 164400 6 la_output[88]
port 567 nsew signal tristate
rlabel metal2 s 302330 163200 302386 164400 6 la_output[89]
port 568 nsew signal tristate
rlabel metal2 s 29826 163200 29882 164400 6 la_output[8]
port 569 nsew signal tristate
rlabel metal2 s 305642 163200 305698 164400 6 la_output[90]
port 570 nsew signal tristate
rlabel metal2 s 309046 163200 309102 164400 6 la_output[91]
port 571 nsew signal tristate
rlabel metal2 s 312450 163200 312506 164400 6 la_output[92]
port 572 nsew signal tristate
rlabel metal2 s 315762 163200 315818 164400 6 la_output[93]
port 573 nsew signal tristate
rlabel metal2 s 319166 163200 319222 164400 6 la_output[94]
port 574 nsew signal tristate
rlabel metal2 s 322478 163200 322534 164400 6 la_output[95]
port 575 nsew signal tristate
rlabel metal2 s 325882 163200 325938 164400 6 la_output[96]
port 576 nsew signal tristate
rlabel metal2 s 329194 163200 329250 164400 6 la_output[97]
port 577 nsew signal tristate
rlabel metal2 s 332598 163200 332654 164400 6 la_output[98]
port 578 nsew signal tristate
rlabel metal2 s 336002 163200 336058 164400 6 la_output[99]
port 579 nsew signal tristate
rlabel metal2 s 33138 163200 33194 164400 6 la_output[9]
port 580 nsew signal tristate
rlabel metal2 s 431038 163200 431094 164400 6 mprj_ack_i
port 581 nsew signal input
rlabel metal2 s 435178 163200 435234 164400 6 mprj_adr_o[0]
port 582 nsew signal tristate
rlabel metal2 s 463790 163200 463846 164400 6 mprj_adr_o[10]
port 583 nsew signal tristate
rlabel metal2 s 466366 163200 466422 164400 6 mprj_adr_o[11]
port 584 nsew signal tristate
rlabel metal2 s 468850 163200 468906 164400 6 mprj_adr_o[12]
port 585 nsew signal tristate
rlabel metal2 s 471426 163200 471482 164400 6 mprj_adr_o[13]
port 586 nsew signal tristate
rlabel metal2 s 473910 163200 473966 164400 6 mprj_adr_o[14]
port 587 nsew signal tristate
rlabel metal2 s 476394 163200 476450 164400 6 mprj_adr_o[15]
port 588 nsew signal tristate
rlabel metal2 s 478970 163200 479026 164400 6 mprj_adr_o[16]
port 589 nsew signal tristate
rlabel metal2 s 481454 163200 481510 164400 6 mprj_adr_o[17]
port 590 nsew signal tristate
rlabel metal2 s 484030 163200 484086 164400 6 mprj_adr_o[18]
port 591 nsew signal tristate
rlabel metal2 s 486514 163200 486570 164400 6 mprj_adr_o[19]
port 592 nsew signal tristate
rlabel metal2 s 438582 163200 438638 164400 6 mprj_adr_o[1]
port 593 nsew signal tristate
rlabel metal2 s 489090 163200 489146 164400 6 mprj_adr_o[20]
port 594 nsew signal tristate
rlabel metal2 s 491574 163200 491630 164400 6 mprj_adr_o[21]
port 595 nsew signal tristate
rlabel metal2 s 494058 163200 494114 164400 6 mprj_adr_o[22]
port 596 nsew signal tristate
rlabel metal2 s 496634 163200 496690 164400 6 mprj_adr_o[23]
port 597 nsew signal tristate
rlabel metal2 s 499118 163200 499174 164400 6 mprj_adr_o[24]
port 598 nsew signal tristate
rlabel metal2 s 501694 163200 501750 164400 6 mprj_adr_o[25]
port 599 nsew signal tristate
rlabel metal2 s 504178 163200 504234 164400 6 mprj_adr_o[26]
port 600 nsew signal tristate
rlabel metal2 s 506754 163200 506810 164400 6 mprj_adr_o[27]
port 601 nsew signal tristate
rlabel metal2 s 509238 163200 509294 164400 6 mprj_adr_o[28]
port 602 nsew signal tristate
rlabel metal2 s 511722 163200 511778 164400 6 mprj_adr_o[29]
port 603 nsew signal tristate
rlabel metal2 s 441986 163200 442042 164400 6 mprj_adr_o[2]
port 604 nsew signal tristate
rlabel metal2 s 514298 163200 514354 164400 6 mprj_adr_o[30]
port 605 nsew signal tristate
rlabel metal2 s 516782 163200 516838 164400 6 mprj_adr_o[31]
port 606 nsew signal tristate
rlabel metal2 s 445298 163200 445354 164400 6 mprj_adr_o[3]
port 607 nsew signal tristate
rlabel metal2 s 448702 163200 448758 164400 6 mprj_adr_o[4]
port 608 nsew signal tristate
rlabel metal2 s 451186 163200 451242 164400 6 mprj_adr_o[5]
port 609 nsew signal tristate
rlabel metal2 s 453762 163200 453818 164400 6 mprj_adr_o[6]
port 610 nsew signal tristate
rlabel metal2 s 456246 163200 456302 164400 6 mprj_adr_o[7]
port 611 nsew signal tristate
rlabel metal2 s 458730 163200 458786 164400 6 mprj_adr_o[8]
port 612 nsew signal tristate
rlabel metal2 s 461306 163200 461362 164400 6 mprj_adr_o[9]
port 613 nsew signal tristate
rlabel metal2 s 431866 163200 431922 164400 6 mprj_cyc_o
port 614 nsew signal tristate
rlabel metal2 s 436098 163200 436154 164400 6 mprj_dat_i[0]
port 615 nsew signal input
rlabel metal2 s 464618 163200 464674 164400 6 mprj_dat_i[10]
port 616 nsew signal input
rlabel metal2 s 467194 163200 467250 164400 6 mprj_dat_i[11]
port 617 nsew signal input
rlabel metal2 s 469678 163200 469734 164400 6 mprj_dat_i[12]
port 618 nsew signal input
rlabel metal2 s 472254 163200 472310 164400 6 mprj_dat_i[13]
port 619 nsew signal input
rlabel metal2 s 474738 163200 474794 164400 6 mprj_dat_i[14]
port 620 nsew signal input
rlabel metal2 s 477314 163200 477370 164400 6 mprj_dat_i[15]
port 621 nsew signal input
rlabel metal2 s 479798 163200 479854 164400 6 mprj_dat_i[16]
port 622 nsew signal input
rlabel metal2 s 482282 163200 482338 164400 6 mprj_dat_i[17]
port 623 nsew signal input
rlabel metal2 s 484858 163200 484914 164400 6 mprj_dat_i[18]
port 624 nsew signal input
rlabel metal2 s 487342 163200 487398 164400 6 mprj_dat_i[19]
port 625 nsew signal input
rlabel metal2 s 439410 163200 439466 164400 6 mprj_dat_i[1]
port 626 nsew signal input
rlabel metal2 s 489918 163200 489974 164400 6 mprj_dat_i[20]
port 627 nsew signal input
rlabel metal2 s 492402 163200 492458 164400 6 mprj_dat_i[21]
port 628 nsew signal input
rlabel metal2 s 494978 163200 495034 164400 6 mprj_dat_i[22]
port 629 nsew signal input
rlabel metal2 s 497462 163200 497518 164400 6 mprj_dat_i[23]
port 630 nsew signal input
rlabel metal2 s 499946 163200 500002 164400 6 mprj_dat_i[24]
port 631 nsew signal input
rlabel metal2 s 502522 163200 502578 164400 6 mprj_dat_i[25]
port 632 nsew signal input
rlabel metal2 s 505006 163200 505062 164400 6 mprj_dat_i[26]
port 633 nsew signal input
rlabel metal2 s 507582 163200 507638 164400 6 mprj_dat_i[27]
port 634 nsew signal input
rlabel metal2 s 510066 163200 510122 164400 6 mprj_dat_i[28]
port 635 nsew signal input
rlabel metal2 s 512642 163200 512698 164400 6 mprj_dat_i[29]
port 636 nsew signal input
rlabel metal2 s 442814 163200 442870 164400 6 mprj_dat_i[2]
port 637 nsew signal input
rlabel metal2 s 515126 163200 515182 164400 6 mprj_dat_i[30]
port 638 nsew signal input
rlabel metal2 s 517610 163200 517666 164400 6 mprj_dat_i[31]
port 639 nsew signal input
rlabel metal2 s 446126 163200 446182 164400 6 mprj_dat_i[3]
port 640 nsew signal input
rlabel metal2 s 449530 163200 449586 164400 6 mprj_dat_i[4]
port 641 nsew signal input
rlabel metal2 s 452014 163200 452070 164400 6 mprj_dat_i[5]
port 642 nsew signal input
rlabel metal2 s 454590 163200 454646 164400 6 mprj_dat_i[6]
port 643 nsew signal input
rlabel metal2 s 457074 163200 457130 164400 6 mprj_dat_i[7]
port 644 nsew signal input
rlabel metal2 s 459650 163200 459706 164400 6 mprj_dat_i[8]
port 645 nsew signal input
rlabel metal2 s 462134 163200 462190 164400 6 mprj_dat_i[9]
port 646 nsew signal input
rlabel metal2 s 436926 163200 436982 164400 6 mprj_dat_o[0]
port 647 nsew signal tristate
rlabel metal2 s 465538 163200 465594 164400 6 mprj_dat_o[10]
port 648 nsew signal tristate
rlabel metal2 s 468022 163200 468078 164400 6 mprj_dat_o[11]
port 649 nsew signal tristate
rlabel metal2 s 470506 163200 470562 164400 6 mprj_dat_o[12]
port 650 nsew signal tristate
rlabel metal2 s 473082 163200 473138 164400 6 mprj_dat_o[13]
port 651 nsew signal tristate
rlabel metal2 s 475566 163200 475622 164400 6 mprj_dat_o[14]
port 652 nsew signal tristate
rlabel metal2 s 478142 163200 478198 164400 6 mprj_dat_o[15]
port 653 nsew signal tristate
rlabel metal2 s 480626 163200 480682 164400 6 mprj_dat_o[16]
port 654 nsew signal tristate
rlabel metal2 s 483202 163200 483258 164400 6 mprj_dat_o[17]
port 655 nsew signal tristate
rlabel metal2 s 485686 163200 485742 164400 6 mprj_dat_o[18]
port 656 nsew signal tristate
rlabel metal2 s 488170 163200 488226 164400 6 mprj_dat_o[19]
port 657 nsew signal tristate
rlabel metal2 s 440238 163200 440294 164400 6 mprj_dat_o[1]
port 658 nsew signal tristate
rlabel metal2 s 490746 163200 490802 164400 6 mprj_dat_o[20]
port 659 nsew signal tristate
rlabel metal2 s 493230 163200 493286 164400 6 mprj_dat_o[21]
port 660 nsew signal tristate
rlabel metal2 s 495806 163200 495862 164400 6 mprj_dat_o[22]
port 661 nsew signal tristate
rlabel metal2 s 498290 163200 498346 164400 6 mprj_dat_o[23]
port 662 nsew signal tristate
rlabel metal2 s 500866 163200 500922 164400 6 mprj_dat_o[24]
port 663 nsew signal tristate
rlabel metal2 s 503350 163200 503406 164400 6 mprj_dat_o[25]
port 664 nsew signal tristate
rlabel metal2 s 505834 163200 505890 164400 6 mprj_dat_o[26]
port 665 nsew signal tristate
rlabel metal2 s 508410 163200 508466 164400 6 mprj_dat_o[27]
port 666 nsew signal tristate
rlabel metal2 s 510894 163200 510950 164400 6 mprj_dat_o[28]
port 667 nsew signal tristate
rlabel metal2 s 513470 163200 513526 164400 6 mprj_dat_o[29]
port 668 nsew signal tristate
rlabel metal2 s 443642 163200 443698 164400 6 mprj_dat_o[2]
port 669 nsew signal tristate
rlabel metal2 s 515954 163200 516010 164400 6 mprj_dat_o[30]
port 670 nsew signal tristate
rlabel metal2 s 518530 163200 518586 164400 6 mprj_dat_o[31]
port 671 nsew signal tristate
rlabel metal2 s 446954 163200 447010 164400 6 mprj_dat_o[3]
port 672 nsew signal tristate
rlabel metal2 s 450358 163200 450414 164400 6 mprj_dat_o[4]
port 673 nsew signal tristate
rlabel metal2 s 452842 163200 452898 164400 6 mprj_dat_o[5]
port 674 nsew signal tristate
rlabel metal2 s 455418 163200 455474 164400 6 mprj_dat_o[6]
port 675 nsew signal tristate
rlabel metal2 s 457902 163200 457958 164400 6 mprj_dat_o[7]
port 676 nsew signal tristate
rlabel metal2 s 460478 163200 460534 164400 6 mprj_dat_o[8]
port 677 nsew signal tristate
rlabel metal2 s 462962 163200 463018 164400 6 mprj_dat_o[9]
port 678 nsew signal tristate
rlabel metal2 s 437754 163200 437810 164400 6 mprj_sel_o[0]
port 679 nsew signal tristate
rlabel metal2 s 441066 163200 441122 164400 6 mprj_sel_o[1]
port 680 nsew signal tristate
rlabel metal2 s 444470 163200 444526 164400 6 mprj_sel_o[2]
port 681 nsew signal tristate
rlabel metal2 s 447874 163200 447930 164400 6 mprj_sel_o[3]
port 682 nsew signal tristate
rlabel metal2 s 432694 163200 432750 164400 6 mprj_stb_o
port 683 nsew signal tristate
rlabel metal2 s 433522 163200 433578 164400 6 mprj_wb_iena
port 684 nsew signal tristate
rlabel metal2 s 434350 163200 434406 164400 6 mprj_we_o
port 685 nsew signal tristate
rlabel metal3 s 523200 89360 524400 89480 6 qspi_enabled
port 686 nsew signal tristate
rlabel metal3 s 523200 83376 524400 83496 6 ser_rx
port 687 nsew signal input
rlabel metal3 s 523200 84872 524400 84992 6 ser_tx
port 688 nsew signal tristate
rlabel metal3 s 523200 80384 524400 80504 6 spi_csb
port 689 nsew signal tristate
rlabel metal3 s 523200 86368 524400 86488 6 spi_enabled
port 690 nsew signal tristate
rlabel metal3 s 523200 78888 524400 79008 6 spi_sck
port 691 nsew signal tristate
rlabel metal3 s 523200 81880 524400 82000 6 spi_sdi
port 692 nsew signal input
rlabel metal3 s 523200 77392 524400 77512 6 spi_sdo
port 693 nsew signal tristate
rlabel metal3 s 523200 75896 524400 76016 6 spi_sdoenb
port 694 nsew signal tristate
rlabel metal3 s 523200 2184 524400 2304 6 sram_ro_addr[0]
port 695 nsew signal input
rlabel metal3 s 523200 3680 524400 3800 6 sram_ro_addr[1]
port 696 nsew signal input
rlabel metal3 s 523200 5176 524400 5296 6 sram_ro_addr[2]
port 697 nsew signal input
rlabel metal3 s 523200 6672 524400 6792 6 sram_ro_addr[3]
port 698 nsew signal input
rlabel metal3 s 523200 8168 524400 8288 6 sram_ro_addr[4]
port 699 nsew signal input
rlabel metal3 s 523200 9664 524400 9784 6 sram_ro_addr[5]
port 700 nsew signal input
rlabel metal3 s 523200 11160 524400 11280 6 sram_ro_addr[6]
port 701 nsew signal input
rlabel metal3 s 523200 12656 524400 12776 6 sram_ro_addr[7]
port 702 nsew signal input
rlabel metal3 s 523200 14152 524400 14272 6 sram_ro_clk
port 703 nsew signal input
rlabel metal3 s 523200 688 524400 808 6 sram_ro_csb
port 704 nsew signal input
rlabel metal3 s 523200 15648 524400 15768 6 sram_ro_data[0]
port 705 nsew signal tristate
rlabel metal3 s 523200 30744 524400 30864 6 sram_ro_data[10]
port 706 nsew signal tristate
rlabel metal3 s 523200 32240 524400 32360 6 sram_ro_data[11]
port 707 nsew signal tristate
rlabel metal3 s 523200 33736 524400 33856 6 sram_ro_data[12]
port 708 nsew signal tristate
rlabel metal3 s 523200 35232 524400 35352 6 sram_ro_data[13]
port 709 nsew signal tristate
rlabel metal3 s 523200 36728 524400 36848 6 sram_ro_data[14]
port 710 nsew signal tristate
rlabel metal3 s 523200 38224 524400 38344 6 sram_ro_data[15]
port 711 nsew signal tristate
rlabel metal3 s 523200 39720 524400 39840 6 sram_ro_data[16]
port 712 nsew signal tristate
rlabel metal3 s 523200 41216 524400 41336 6 sram_ro_data[17]
port 713 nsew signal tristate
rlabel metal3 s 523200 42712 524400 42832 6 sram_ro_data[18]
port 714 nsew signal tristate
rlabel metal3 s 523200 44208 524400 44328 6 sram_ro_data[19]
port 715 nsew signal tristate
rlabel metal3 s 523200 17144 524400 17264 6 sram_ro_data[1]
port 716 nsew signal tristate
rlabel metal3 s 523200 45704 524400 45824 6 sram_ro_data[20]
port 717 nsew signal tristate
rlabel metal3 s 523200 47200 524400 47320 6 sram_ro_data[21]
port 718 nsew signal tristate
rlabel metal3 s 523200 48832 524400 48952 6 sram_ro_data[22]
port 719 nsew signal tristate
rlabel metal3 s 523200 50328 524400 50448 6 sram_ro_data[23]
port 720 nsew signal tristate
rlabel metal3 s 523200 51824 524400 51944 6 sram_ro_data[24]
port 721 nsew signal tristate
rlabel metal3 s 523200 53320 524400 53440 6 sram_ro_data[25]
port 722 nsew signal tristate
rlabel metal3 s 523200 54816 524400 54936 6 sram_ro_data[26]
port 723 nsew signal tristate
rlabel metal3 s 523200 56312 524400 56432 6 sram_ro_data[27]
port 724 nsew signal tristate
rlabel metal3 s 523200 57808 524400 57928 6 sram_ro_data[28]
port 725 nsew signal tristate
rlabel metal3 s 523200 59304 524400 59424 6 sram_ro_data[29]
port 726 nsew signal tristate
rlabel metal3 s 523200 18640 524400 18760 6 sram_ro_data[2]
port 727 nsew signal tristate
rlabel metal3 s 523200 60800 524400 60920 6 sram_ro_data[30]
port 728 nsew signal tristate
rlabel metal3 s 523200 62296 524400 62416 6 sram_ro_data[31]
port 729 nsew signal tristate
rlabel metal3 s 523200 20136 524400 20256 6 sram_ro_data[3]
port 730 nsew signal tristate
rlabel metal3 s 523200 21632 524400 21752 6 sram_ro_data[4]
port 731 nsew signal tristate
rlabel metal3 s 523200 23128 524400 23248 6 sram_ro_data[5]
port 732 nsew signal tristate
rlabel metal3 s 523200 24760 524400 24880 6 sram_ro_data[6]
port 733 nsew signal tristate
rlabel metal3 s 523200 26256 524400 26376 6 sram_ro_data[7]
port 734 nsew signal tristate
rlabel metal3 s 523200 27752 524400 27872 6 sram_ro_data[8]
port 735 nsew signal tristate
rlabel metal3 s 523200 29248 524400 29368 6 sram_ro_data[9]
port 736 nsew signal tristate
rlabel metal3 s 523200 69776 524400 69896 6 trap
port 737 nsew signal tristate
rlabel metal3 s 523200 87864 524400 87984 6 uart_enabled
port 738 nsew signal tristate
rlabel metal2 s 519358 163200 519414 164400 6 user_irq_ena[0]
port 739 nsew signal tristate
rlabel metal2 s 520186 163200 520242 164400 6 user_irq_ena[1]
port 740 nsew signal tristate
rlabel metal2 s 521014 163200 521070 164400 6 user_irq_ena[2]
port 741 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 524000 164000
<< end >>
