VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mgmt_core_wrapper
  CLASS BLOCK ;
  FOREIGN mgmt_core_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2700.000 BY 820.000 ;
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 91.730 10.000 93.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 580.000 91.730 640.000 93.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 2660.000 91.730 2694.220 93.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 221.730 10.000 223.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 580.000 221.730 640.000 223.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 2660.000 221.730 2694.220 223.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 351.730 10.000 353.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 580.000 351.730 640.000 353.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 2660.000 351.730 2694.220 353.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 481.730 10.000 483.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 580.000 481.730 640.000 483.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 2660.000 481.730 2694.220 483.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 611.730 10.000 613.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 580.000 611.730 640.000 613.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 2660.000 611.730 2694.220 613.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 741.730 10.000 743.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 580.000 741.730 640.000 743.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 2660.000 741.730 2694.220 743.330 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.730 10.000 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 580.000 26.730 640.000 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 2660.000 26.730 2694.220 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 156.730 10.000 158.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 580.000 156.730 640.000 158.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 2660.000 156.730 2694.220 158.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 286.730 10.000 288.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 580.000 286.730 640.000 288.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 2660.000 286.730 2694.220 288.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 416.730 10.000 418.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 580.000 416.730 640.000 418.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 2660.000 416.730 2694.220 418.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 546.730 10.000 548.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 580.000 546.730 640.000 548.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 2660.000 546.730 2694.220 548.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 676.730 10.000 678.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 580.000 676.730 640.000 678.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 2660.000 676.730 2694.220 678.330 ;
    END
  END VPWR
  PIN core_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2531.010 0.000 2531.290 4.000 ;
    END
  END core_clk
  PIN core_rstn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END core_rstn
  PIN debug_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 322.360 2700.000 322.960 ;
    END
  END debug_in
  PIN debug_mode
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 329.840 2700.000 330.440 ;
    END
  END debug_mode
  PIN debug_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 337.320 2700.000 337.920 ;
    END
  END debug_oeb
  PIN debug_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 344.800 2700.000 345.400 ;
    END
  END debug_out
  PIN flash_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 724.240 2700.000 724.840 ;
    END
  END flash_clk
  PIN flash_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 716.760 2700.000 717.360 ;
    END
  END flash_csb
  PIN flash_io0_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 732.400 2700.000 733.000 ;
    END
  END flash_io0_di
  PIN flash_io0_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 739.880 2700.000 740.480 ;
    END
  END flash_io0_do
  PIN flash_io0_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 747.360 2700.000 747.960 ;
    END
  END flash_io0_oeb
  PIN flash_io1_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 754.840 2700.000 755.440 ;
    END
  END flash_io1_di
  PIN flash_io1_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 762.320 2700.000 762.920 ;
    END
  END flash_io1_do
  PIN flash_io1_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 769.800 2700.000 770.400 ;
    END
  END flash_io1_oeb
  PIN flash_io2_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 777.960 2700.000 778.560 ;
    END
  END flash_io2_di
  PIN flash_io2_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 785.440 2700.000 786.040 ;
    END
  END flash_io2_do
  PIN flash_io2_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 792.920 2700.000 793.520 ;
    END
  END flash_io2_oeb
  PIN flash_io3_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 800.400 2700.000 801.000 ;
    END
  END flash_io3_di
  PIN flash_io3_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 807.880 2700.000 808.480 ;
    END
  END flash_io3_do
  PIN flash_io3_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 815.360 2700.000 815.960 ;
    END
  END flash_io3_oeb
  PIN gpio_in_pad
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 0.000 505.910 4.000 ;
    END
  END gpio_in_pad
  PIN gpio_inenb_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.270 0.000 843.550 4.000 ;
    END
  END gpio_inenb_pad
  PIN gpio_mode0_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1180.910 0.000 1181.190 4.000 ;
    END
  END gpio_mode0_pad
  PIN gpio_mode1_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1518.550 0.000 1518.830 4.000 ;
    END
  END gpio_mode1_pad
  PIN gpio_out_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1855.730 0.000 1856.010 4.000 ;
    END
  END gpio_out_pad
  PIN gpio_outenb_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2193.370 0.000 2193.650 4.000 ;
    END
  END gpio_outenb_pad
  PIN hk_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 459.040 2700.000 459.640 ;
    END
  END hk_ack_i
  PIN hk_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 474.000 2700.000 474.600 ;
    END
  END hk_dat_i[0]
  PIN hk_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 550.160 2700.000 550.760 ;
    END
  END hk_dat_i[10]
  PIN hk_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 557.640 2700.000 558.240 ;
    END
  END hk_dat_i[11]
  PIN hk_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 565.120 2700.000 565.720 ;
    END
  END hk_dat_i[12]
  PIN hk_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 572.600 2700.000 573.200 ;
    END
  END hk_dat_i[13]
  PIN hk_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 580.080 2700.000 580.680 ;
    END
  END hk_dat_i[14]
  PIN hk_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 587.560 2700.000 588.160 ;
    END
  END hk_dat_i[15]
  PIN hk_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 595.720 2700.000 596.320 ;
    END
  END hk_dat_i[16]
  PIN hk_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 603.200 2700.000 603.800 ;
    END
  END hk_dat_i[17]
  PIN hk_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 610.680 2700.000 611.280 ;
    END
  END hk_dat_i[18]
  PIN hk_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 618.160 2700.000 618.760 ;
    END
  END hk_dat_i[19]
  PIN hk_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 481.480 2700.000 482.080 ;
    END
  END hk_dat_i[1]
  PIN hk_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 625.640 2700.000 626.240 ;
    END
  END hk_dat_i[20]
  PIN hk_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 633.120 2700.000 633.720 ;
    END
  END hk_dat_i[21]
  PIN hk_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 641.280 2700.000 641.880 ;
    END
  END hk_dat_i[22]
  PIN hk_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 648.760 2700.000 649.360 ;
    END
  END hk_dat_i[23]
  PIN hk_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 656.240 2700.000 656.840 ;
    END
  END hk_dat_i[24]
  PIN hk_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 663.720 2700.000 664.320 ;
    END
  END hk_dat_i[25]
  PIN hk_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 671.200 2700.000 671.800 ;
    END
  END hk_dat_i[26]
  PIN hk_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 678.680 2700.000 679.280 ;
    END
  END hk_dat_i[27]
  PIN hk_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 686.840 2700.000 687.440 ;
    END
  END hk_dat_i[28]
  PIN hk_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 694.320 2700.000 694.920 ;
    END
  END hk_dat_i[29]
  PIN hk_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 488.960 2700.000 489.560 ;
    END
  END hk_dat_i[2]
  PIN hk_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 701.800 2700.000 702.400 ;
    END
  END hk_dat_i[30]
  PIN hk_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 709.280 2700.000 709.880 ;
    END
  END hk_dat_i[31]
  PIN hk_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 496.440 2700.000 497.040 ;
    END
  END hk_dat_i[3]
  PIN hk_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 504.600 2700.000 505.200 ;
    END
  END hk_dat_i[4]
  PIN hk_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 512.080 2700.000 512.680 ;
    END
  END hk_dat_i[5]
  PIN hk_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 519.560 2700.000 520.160 ;
    END
  END hk_dat_i[6]
  PIN hk_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 527.040 2700.000 527.640 ;
    END
  END hk_dat_i[7]
  PIN hk_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 534.520 2700.000 535.120 ;
    END
  END hk_dat_i[8]
  PIN hk_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 542.000 2700.000 542.600 ;
    END
  END hk_dat_i[9]
  PIN hk_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 466.520 2700.000 467.120 ;
    END
  END hk_stb_o
  PIN irq[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2688.790 816.000 2689.070 820.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2693.390 816.000 2693.670 820.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2697.530 816.000 2697.810 820.000 ;
    END
  END irq[2]
  PIN irq[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 375.400 2700.000 376.000 ;
    END
  END irq[3]
  PIN irq[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 367.920 2700.000 368.520 ;
    END
  END irq[4]
  PIN irq[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 359.760 2700.000 360.360 ;
    END
  END irq[5]
  PIN la_iena[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 816.000 2.210 820.000 ;
    END
  END la_iena[0]
  PIN la_iena[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1735.210 816.000 1735.490 820.000 ;
    END
  END la_iena[100]
  PIN la_iena[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1752.690 816.000 1752.970 820.000 ;
    END
  END la_iena[101]
  PIN la_iena[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1770.170 816.000 1770.450 820.000 ;
    END
  END la_iena[102]
  PIN la_iena[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.190 816.000 1787.470 820.000 ;
    END
  END la_iena[103]
  PIN la_iena[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1804.670 816.000 1804.950 820.000 ;
    END
  END la_iena[104]
  PIN la_iena[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1822.150 816.000 1822.430 820.000 ;
    END
  END la_iena[105]
  PIN la_iena[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1839.170 816.000 1839.450 820.000 ;
    END
  END la_iena[106]
  PIN la_iena[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1856.650 816.000 1856.930 820.000 ;
    END
  END la_iena[107]
  PIN la_iena[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1874.130 816.000 1874.410 820.000 ;
    END
  END la_iena[108]
  PIN la_iena[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1891.610 816.000 1891.890 820.000 ;
    END
  END la_iena[109]
  PIN la_iena[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 816.000 175.170 820.000 ;
    END
  END la_iena[10]
  PIN la_iena[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1908.630 816.000 1908.910 820.000 ;
    END
  END la_iena[110]
  PIN la_iena[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1926.110 816.000 1926.390 820.000 ;
    END
  END la_iena[111]
  PIN la_iena[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1943.590 816.000 1943.870 820.000 ;
    END
  END la_iena[112]
  PIN la_iena[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1960.610 816.000 1960.890 820.000 ;
    END
  END la_iena[113]
  PIN la_iena[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1978.090 816.000 1978.370 820.000 ;
    END
  END la_iena[114]
  PIN la_iena[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1995.570 816.000 1995.850 820.000 ;
    END
  END la_iena[115]
  PIN la_iena[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2012.590 816.000 2012.870 820.000 ;
    END
  END la_iena[116]
  PIN la_iena[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2030.070 816.000 2030.350 820.000 ;
    END
  END la_iena[117]
  PIN la_iena[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2047.550 816.000 2047.830 820.000 ;
    END
  END la_iena[118]
  PIN la_iena[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2064.570 816.000 2064.850 820.000 ;
    END
  END la_iena[119]
  PIN la_iena[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 816.000 192.650 820.000 ;
    END
  END la_iena[11]
  PIN la_iena[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2082.050 816.000 2082.330 820.000 ;
    END
  END la_iena[120]
  PIN la_iena[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2099.530 816.000 2099.810 820.000 ;
    END
  END la_iena[121]
  PIN la_iena[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2117.010 816.000 2117.290 820.000 ;
    END
  END la_iena[122]
  PIN la_iena[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2134.030 816.000 2134.310 820.000 ;
    END
  END la_iena[123]
  PIN la_iena[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2151.510 816.000 2151.790 820.000 ;
    END
  END la_iena[124]
  PIN la_iena[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2168.990 816.000 2169.270 820.000 ;
    END
  END la_iena[125]
  PIN la_iena[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2186.010 816.000 2186.290 820.000 ;
    END
  END la_iena[126]
  PIN la_iena[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2203.490 816.000 2203.770 820.000 ;
    END
  END la_iena[127]
  PIN la_iena[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 816.000 210.130 820.000 ;
    END
  END la_iena[12]
  PIN la_iena[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.870 816.000 227.150 820.000 ;
    END
  END la_iena[13]
  PIN la_iena[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 816.000 244.630 820.000 ;
    END
  END la_iena[14]
  PIN la_iena[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 816.000 262.110 820.000 ;
    END
  END la_iena[15]
  PIN la_iena[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 816.000 279.590 820.000 ;
    END
  END la_iena[16]
  PIN la_iena[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 816.000 296.610 820.000 ;
    END
  END la_iena[17]
  PIN la_iena[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.810 816.000 314.090 820.000 ;
    END
  END la_iena[18]
  PIN la_iena[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 816.000 331.570 820.000 ;
    END
  END la_iena[19]
  PIN la_iena[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 816.000 19.230 820.000 ;
    END
  END la_iena[1]
  PIN la_iena[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.310 816.000 348.590 820.000 ;
    END
  END la_iena[20]
  PIN la_iena[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 816.000 366.070 820.000 ;
    END
  END la_iena[21]
  PIN la_iena[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 816.000 383.550 820.000 ;
    END
  END la_iena[22]
  PIN la_iena[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.290 816.000 400.570 820.000 ;
    END
  END la_iena[23]
  PIN la_iena[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.770 816.000 418.050 820.000 ;
    END
  END la_iena[24]
  PIN la_iena[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.250 816.000 435.530 820.000 ;
    END
  END la_iena[25]
  PIN la_iena[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.270 816.000 452.550 820.000 ;
    END
  END la_iena[26]
  PIN la_iena[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.750 816.000 470.030 820.000 ;
    END
  END la_iena[27]
  PIN la_iena[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.230 816.000 487.510 820.000 ;
    END
  END la_iena[28]
  PIN la_iena[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.250 816.000 504.530 820.000 ;
    END
  END la_iena[29]
  PIN la_iena[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 816.000 36.710 820.000 ;
    END
  END la_iena[2]
  PIN la_iena[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 816.000 522.010 820.000 ;
    END
  END la_iena[30]
  PIN la_iena[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.210 816.000 539.490 820.000 ;
    END
  END la_iena[31]
  PIN la_iena[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 816.000 556.970 820.000 ;
    END
  END la_iena[32]
  PIN la_iena[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.710 816.000 573.990 820.000 ;
    END
  END la_iena[33]
  PIN la_iena[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.190 816.000 591.470 820.000 ;
    END
  END la_iena[34]
  PIN la_iena[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 816.000 608.950 820.000 ;
    END
  END la_iena[35]
  PIN la_iena[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.690 816.000 625.970 820.000 ;
    END
  END la_iena[36]
  PIN la_iena[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.170 816.000 643.450 820.000 ;
    END
  END la_iena[37]
  PIN la_iena[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.650 816.000 660.930 820.000 ;
    END
  END la_iena[38]
  PIN la_iena[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.670 816.000 677.950 820.000 ;
    END
  END la_iena[39]
  PIN la_iena[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 816.000 54.190 820.000 ;
    END
  END la_iena[3]
  PIN la_iena[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.150 816.000 695.430 820.000 ;
    END
  END la_iena[40]
  PIN la_iena[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.630 816.000 712.910 820.000 ;
    END
  END la_iena[41]
  PIN la_iena[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.650 816.000 729.930 820.000 ;
    END
  END la_iena[42]
  PIN la_iena[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 816.000 747.410 820.000 ;
    END
  END la_iena[43]
  PIN la_iena[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.610 816.000 764.890 820.000 ;
    END
  END la_iena[44]
  PIN la_iena[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.630 816.000 781.910 820.000 ;
    END
  END la_iena[45]
  PIN la_iena[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.110 816.000 799.390 820.000 ;
    END
  END la_iena[46]
  PIN la_iena[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.590 816.000 816.870 820.000 ;
    END
  END la_iena[47]
  PIN la_iena[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.070 816.000 834.350 820.000 ;
    END
  END la_iena[48]
  PIN la_iena[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.090 816.000 851.370 820.000 ;
    END
  END la_iena[49]
  PIN la_iena[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 816.000 71.210 820.000 ;
    END
  END la_iena[4]
  PIN la_iena[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.570 816.000 868.850 820.000 ;
    END
  END la_iena[50]
  PIN la_iena[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.050 816.000 886.330 820.000 ;
    END
  END la_iena[51]
  PIN la_iena[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.070 816.000 903.350 820.000 ;
    END
  END la_iena[52]
  PIN la_iena[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.550 816.000 920.830 820.000 ;
    END
  END la_iena[53]
  PIN la_iena[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.030 816.000 938.310 820.000 ;
    END
  END la_iena[54]
  PIN la_iena[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.050 816.000 955.330 820.000 ;
    END
  END la_iena[55]
  PIN la_iena[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.530 816.000 972.810 820.000 ;
    END
  END la_iena[56]
  PIN la_iena[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.010 816.000 990.290 820.000 ;
    END
  END la_iena[57]
  PIN la_iena[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.030 816.000 1007.310 820.000 ;
    END
  END la_iena[58]
  PIN la_iena[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.510 816.000 1024.790 820.000 ;
    END
  END la_iena[59]
  PIN la_iena[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 816.000 88.690 820.000 ;
    END
  END la_iena[5]
  PIN la_iena[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1041.990 816.000 1042.270 820.000 ;
    END
  END la_iena[60]
  PIN la_iena[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.470 816.000 1059.750 820.000 ;
    END
  END la_iena[61]
  PIN la_iena[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.490 816.000 1076.770 820.000 ;
    END
  END la_iena[62]
  PIN la_iena[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1093.970 816.000 1094.250 820.000 ;
    END
  END la_iena[63]
  PIN la_iena[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1111.450 816.000 1111.730 820.000 ;
    END
  END la_iena[64]
  PIN la_iena[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.470 816.000 1128.750 820.000 ;
    END
  END la_iena[65]
  PIN la_iena[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.950 816.000 1146.230 820.000 ;
    END
  END la_iena[66]
  PIN la_iena[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1163.430 816.000 1163.710 820.000 ;
    END
  END la_iena[67]
  PIN la_iena[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1180.450 816.000 1180.730 820.000 ;
    END
  END la_iena[68]
  PIN la_iena[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.930 816.000 1198.210 820.000 ;
    END
  END la_iena[69]
  PIN la_iena[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 816.000 106.170 820.000 ;
    END
  END la_iena[6]
  PIN la_iena[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1215.410 816.000 1215.690 820.000 ;
    END
  END la_iena[70]
  PIN la_iena[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1232.430 816.000 1232.710 820.000 ;
    END
  END la_iena[71]
  PIN la_iena[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.910 816.000 1250.190 820.000 ;
    END
  END la_iena[72]
  PIN la_iena[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1267.390 816.000 1267.670 820.000 ;
    END
  END la_iena[73]
  PIN la_iena[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1284.410 816.000 1284.690 820.000 ;
    END
  END la_iena[74]
  PIN la_iena[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1301.890 816.000 1302.170 820.000 ;
    END
  END la_iena[75]
  PIN la_iena[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1319.370 816.000 1319.650 820.000 ;
    END
  END la_iena[76]
  PIN la_iena[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1336.850 816.000 1337.130 820.000 ;
    END
  END la_iena[77]
  PIN la_iena[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1353.870 816.000 1354.150 820.000 ;
    END
  END la_iena[78]
  PIN la_iena[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1371.350 816.000 1371.630 820.000 ;
    END
  END la_iena[79]
  PIN la_iena[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 816.000 123.190 820.000 ;
    END
  END la_iena[7]
  PIN la_iena[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1388.830 816.000 1389.110 820.000 ;
    END
  END la_iena[80]
  PIN la_iena[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1405.850 816.000 1406.130 820.000 ;
    END
  END la_iena[81]
  PIN la_iena[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1423.330 816.000 1423.610 820.000 ;
    END
  END la_iena[82]
  PIN la_iena[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1440.810 816.000 1441.090 820.000 ;
    END
  END la_iena[83]
  PIN la_iena[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1457.830 816.000 1458.110 820.000 ;
    END
  END la_iena[84]
  PIN la_iena[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1475.310 816.000 1475.590 820.000 ;
    END
  END la_iena[85]
  PIN la_iena[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1492.790 816.000 1493.070 820.000 ;
    END
  END la_iena[86]
  PIN la_iena[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1509.810 816.000 1510.090 820.000 ;
    END
  END la_iena[87]
  PIN la_iena[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1527.290 816.000 1527.570 820.000 ;
    END
  END la_iena[88]
  PIN la_iena[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1544.770 816.000 1545.050 820.000 ;
    END
  END la_iena[89]
  PIN la_iena[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 816.000 140.670 820.000 ;
    END
  END la_iena[8]
  PIN la_iena[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1561.790 816.000 1562.070 820.000 ;
    END
  END la_iena[90]
  PIN la_iena[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1579.270 816.000 1579.550 820.000 ;
    END
  END la_iena[91]
  PIN la_iena[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1596.750 816.000 1597.030 820.000 ;
    END
  END la_iena[92]
  PIN la_iena[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1614.230 816.000 1614.510 820.000 ;
    END
  END la_iena[93]
  PIN la_iena[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1631.250 816.000 1631.530 820.000 ;
    END
  END la_iena[94]
  PIN la_iena[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1648.730 816.000 1649.010 820.000 ;
    END
  END la_iena[95]
  PIN la_iena[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1666.210 816.000 1666.490 820.000 ;
    END
  END la_iena[96]
  PIN la_iena[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1683.230 816.000 1683.510 820.000 ;
    END
  END la_iena[97]
  PIN la_iena[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1700.710 816.000 1700.990 820.000 ;
    END
  END la_iena[98]
  PIN la_iena[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1718.190 816.000 1718.470 820.000 ;
    END
  END la_iena[99]
  PIN la_iena[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 816.000 158.150 820.000 ;
    END
  END la_iena[9]
  PIN la_input[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 816.000 6.350 820.000 ;
    END
  END la_input[0]
  PIN la_input[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1739.810 816.000 1740.090 820.000 ;
    END
  END la_input[100]
  PIN la_input[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1756.830 816.000 1757.110 820.000 ;
    END
  END la_input[101]
  PIN la_input[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1774.310 816.000 1774.590 820.000 ;
    END
  END la_input[102]
  PIN la_input[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1791.790 816.000 1792.070 820.000 ;
    END
  END la_input[103]
  PIN la_input[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1809.270 816.000 1809.550 820.000 ;
    END
  END la_input[104]
  PIN la_input[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1826.290 816.000 1826.570 820.000 ;
    END
  END la_input[105]
  PIN la_input[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1843.770 816.000 1844.050 820.000 ;
    END
  END la_input[106]
  PIN la_input[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1861.250 816.000 1861.530 820.000 ;
    END
  END la_input[107]
  PIN la_input[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1878.270 816.000 1878.550 820.000 ;
    END
  END la_input[108]
  PIN la_input[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1895.750 816.000 1896.030 820.000 ;
    END
  END la_input[109]
  PIN la_input[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 816.000 179.770 820.000 ;
    END
  END la_input[10]
  PIN la_input[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1913.230 816.000 1913.510 820.000 ;
    END
  END la_input[110]
  PIN la_input[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1930.250 816.000 1930.530 820.000 ;
    END
  END la_input[111]
  PIN la_input[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1947.730 816.000 1948.010 820.000 ;
    END
  END la_input[112]
  PIN la_input[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1965.210 816.000 1965.490 820.000 ;
    END
  END la_input[113]
  PIN la_input[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1982.230 816.000 1982.510 820.000 ;
    END
  END la_input[114]
  PIN la_input[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1999.710 816.000 1999.990 820.000 ;
    END
  END la_input[115]
  PIN la_input[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2017.190 816.000 2017.470 820.000 ;
    END
  END la_input[116]
  PIN la_input[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2034.210 816.000 2034.490 820.000 ;
    END
  END la_input[117]
  PIN la_input[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2051.690 816.000 2051.970 820.000 ;
    END
  END la_input[118]
  PIN la_input[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2069.170 816.000 2069.450 820.000 ;
    END
  END la_input[119]
  PIN la_input[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 816.000 196.790 820.000 ;
    END
  END la_input[11]
  PIN la_input[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2086.650 816.000 2086.930 820.000 ;
    END
  END la_input[120]
  PIN la_input[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2103.670 816.000 2103.950 820.000 ;
    END
  END la_input[121]
  PIN la_input[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2121.150 816.000 2121.430 820.000 ;
    END
  END la_input[122]
  PIN la_input[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2138.630 816.000 2138.910 820.000 ;
    END
  END la_input[123]
  PIN la_input[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2155.650 816.000 2155.930 820.000 ;
    END
  END la_input[124]
  PIN la_input[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2173.130 816.000 2173.410 820.000 ;
    END
  END la_input[125]
  PIN la_input[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2190.610 816.000 2190.890 820.000 ;
    END
  END la_input[126]
  PIN la_input[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2207.630 816.000 2207.910 820.000 ;
    END
  END la_input[127]
  PIN la_input[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 816.000 214.270 820.000 ;
    END
  END la_input[12]
  PIN la_input[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 816.000 231.750 820.000 ;
    END
  END la_input[13]
  PIN la_input[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 816.000 249.230 820.000 ;
    END
  END la_input[14]
  PIN la_input[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 816.000 266.250 820.000 ;
    END
  END la_input[15]
  PIN la_input[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 816.000 283.730 820.000 ;
    END
  END la_input[16]
  PIN la_input[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 816.000 301.210 820.000 ;
    END
  END la_input[17]
  PIN la_input[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 816.000 318.230 820.000 ;
    END
  END la_input[18]
  PIN la_input[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 816.000 335.710 820.000 ;
    END
  END la_input[19]
  PIN la_input[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 816.000 23.830 820.000 ;
    END
  END la_input[1]
  PIN la_input[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.910 816.000 353.190 820.000 ;
    END
  END la_input[20]
  PIN la_input[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.930 816.000 370.210 820.000 ;
    END
  END la_input[21]
  PIN la_input[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.410 816.000 387.690 820.000 ;
    END
  END la_input[22]
  PIN la_input[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.890 816.000 405.170 820.000 ;
    END
  END la_input[23]
  PIN la_input[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 816.000 422.190 820.000 ;
    END
  END la_input[24]
  PIN la_input[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 816.000 439.670 820.000 ;
    END
  END la_input[25]
  PIN la_input[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.870 816.000 457.150 820.000 ;
    END
  END la_input[26]
  PIN la_input[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.350 816.000 474.630 820.000 ;
    END
  END la_input[27]
  PIN la_input[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.370 816.000 491.650 820.000 ;
    END
  END la_input[28]
  PIN la_input[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 816.000 509.130 820.000 ;
    END
  END la_input[29]
  PIN la_input[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 816.000 40.850 820.000 ;
    END
  END la_input[2]
  PIN la_input[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.330 816.000 526.610 820.000 ;
    END
  END la_input[30]
  PIN la_input[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.350 816.000 543.630 820.000 ;
    END
  END la_input[31]
  PIN la_input[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.830 816.000 561.110 820.000 ;
    END
  END la_input[32]
  PIN la_input[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.310 816.000 578.590 820.000 ;
    END
  END la_input[33]
  PIN la_input[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.330 816.000 595.610 820.000 ;
    END
  END la_input[34]
  PIN la_input[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.810 816.000 613.090 820.000 ;
    END
  END la_input[35]
  PIN la_input[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.290 816.000 630.570 820.000 ;
    END
  END la_input[36]
  PIN la_input[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.310 816.000 647.590 820.000 ;
    END
  END la_input[37]
  PIN la_input[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.790 816.000 665.070 820.000 ;
    END
  END la_input[38]
  PIN la_input[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.270 816.000 682.550 820.000 ;
    END
  END la_input[39]
  PIN la_input[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 816.000 58.330 820.000 ;
    END
  END la_input[3]
  PIN la_input[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.290 816.000 699.570 820.000 ;
    END
  END la_input[40]
  PIN la_input[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.770 816.000 717.050 820.000 ;
    END
  END la_input[41]
  PIN la_input[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 816.000 734.530 820.000 ;
    END
  END la_input[42]
  PIN la_input[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 751.730 816.000 752.010 820.000 ;
    END
  END la_input[43]
  PIN la_input[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.750 816.000 769.030 820.000 ;
    END
  END la_input[44]
  PIN la_input[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.230 816.000 786.510 820.000 ;
    END
  END la_input[45]
  PIN la_input[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.710 816.000 803.990 820.000 ;
    END
  END la_input[46]
  PIN la_input[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.730 816.000 821.010 820.000 ;
    END
  END la_input[47]
  PIN la_input[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.210 816.000 838.490 820.000 ;
    END
  END la_input[48]
  PIN la_input[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.690 816.000 855.970 820.000 ;
    END
  END la_input[49]
  PIN la_input[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 816.000 75.810 820.000 ;
    END
  END la_input[4]
  PIN la_input[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.710 816.000 872.990 820.000 ;
    END
  END la_input[50]
  PIN la_input[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 890.190 816.000 890.470 820.000 ;
    END
  END la_input[51]
  PIN la_input[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.670 816.000 907.950 820.000 ;
    END
  END la_input[52]
  PIN la_input[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.690 816.000 924.970 820.000 ;
    END
  END la_input[53]
  PIN la_input[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.170 816.000 942.450 820.000 ;
    END
  END la_input[54]
  PIN la_input[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.650 816.000 959.930 820.000 ;
    END
  END la_input[55]
  PIN la_input[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.670 816.000 976.950 820.000 ;
    END
  END la_input[56]
  PIN la_input[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 994.150 816.000 994.430 820.000 ;
    END
  END la_input[57]
  PIN la_input[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1011.630 816.000 1011.910 820.000 ;
    END
  END la_input[58]
  PIN la_input[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1029.110 816.000 1029.390 820.000 ;
    END
  END la_input[59]
  PIN la_input[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 816.000 92.830 820.000 ;
    END
  END la_input[5]
  PIN la_input[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.130 816.000 1046.410 820.000 ;
    END
  END la_input[60]
  PIN la_input[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1063.610 816.000 1063.890 820.000 ;
    END
  END la_input[61]
  PIN la_input[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1081.090 816.000 1081.370 820.000 ;
    END
  END la_input[62]
  PIN la_input[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.110 816.000 1098.390 820.000 ;
    END
  END la_input[63]
  PIN la_input[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1115.590 816.000 1115.870 820.000 ;
    END
  END la_input[64]
  PIN la_input[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.070 816.000 1133.350 820.000 ;
    END
  END la_input[65]
  PIN la_input[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1150.090 816.000 1150.370 820.000 ;
    END
  END la_input[66]
  PIN la_input[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1167.570 816.000 1167.850 820.000 ;
    END
  END la_input[67]
  PIN la_input[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.050 816.000 1185.330 820.000 ;
    END
  END la_input[68]
  PIN la_input[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.070 816.000 1202.350 820.000 ;
    END
  END la_input[69]
  PIN la_input[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 816.000 110.310 820.000 ;
    END
  END la_input[6]
  PIN la_input[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1219.550 816.000 1219.830 820.000 ;
    END
  END la_input[70]
  PIN la_input[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1237.030 816.000 1237.310 820.000 ;
    END
  END la_input[71]
  PIN la_input[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1254.510 816.000 1254.790 820.000 ;
    END
  END la_input[72]
  PIN la_input[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.530 816.000 1271.810 820.000 ;
    END
  END la_input[73]
  PIN la_input[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1289.010 816.000 1289.290 820.000 ;
    END
  END la_input[74]
  PIN la_input[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1306.490 816.000 1306.770 820.000 ;
    END
  END la_input[75]
  PIN la_input[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.510 816.000 1323.790 820.000 ;
    END
  END la_input[76]
  PIN la_input[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.990 816.000 1341.270 820.000 ;
    END
  END la_input[77]
  PIN la_input[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.470 816.000 1358.750 820.000 ;
    END
  END la_input[78]
  PIN la_input[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.490 816.000 1375.770 820.000 ;
    END
  END la_input[79]
  PIN la_input[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 816.000 127.790 820.000 ;
    END
  END la_input[7]
  PIN la_input[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1392.970 816.000 1393.250 820.000 ;
    END
  END la_input[80]
  PIN la_input[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1410.450 816.000 1410.730 820.000 ;
    END
  END la_input[81]
  PIN la_input[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1427.470 816.000 1427.750 820.000 ;
    END
  END la_input[82]
  PIN la_input[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1444.950 816.000 1445.230 820.000 ;
    END
  END la_input[83]
  PIN la_input[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.430 816.000 1462.710 820.000 ;
    END
  END la_input[84]
  PIN la_input[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1479.450 816.000 1479.730 820.000 ;
    END
  END la_input[85]
  PIN la_input[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1496.930 816.000 1497.210 820.000 ;
    END
  END la_input[86]
  PIN la_input[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1514.410 816.000 1514.690 820.000 ;
    END
  END la_input[87]
  PIN la_input[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1531.890 816.000 1532.170 820.000 ;
    END
  END la_input[88]
  PIN la_input[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1548.910 816.000 1549.190 820.000 ;
    END
  END la_input[89]
  PIN la_input[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 816.000 144.810 820.000 ;
    END
  END la_input[8]
  PIN la_input[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1566.390 816.000 1566.670 820.000 ;
    END
  END la_input[90]
  PIN la_input[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1583.870 816.000 1584.150 820.000 ;
    END
  END la_input[91]
  PIN la_input[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1600.890 816.000 1601.170 820.000 ;
    END
  END la_input[92]
  PIN la_input[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1618.370 816.000 1618.650 820.000 ;
    END
  END la_input[93]
  PIN la_input[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1635.850 816.000 1636.130 820.000 ;
    END
  END la_input[94]
  PIN la_input[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1652.870 816.000 1653.150 820.000 ;
    END
  END la_input[95]
  PIN la_input[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1670.350 816.000 1670.630 820.000 ;
    END
  END la_input[96]
  PIN la_input[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.830 816.000 1688.110 820.000 ;
    END
  END la_input[97]
  PIN la_input[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1704.850 816.000 1705.130 820.000 ;
    END
  END la_input[98]
  PIN la_input[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1722.330 816.000 1722.610 820.000 ;
    END
  END la_input[99]
  PIN la_input[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 816.000 162.290 820.000 ;
    END
  END la_input[9]
  PIN la_oenb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 816.000 10.490 820.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.950 816.000 1744.230 820.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1761.430 816.000 1761.710 820.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1778.910 816.000 1779.190 820.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1795.930 816.000 1796.210 820.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1813.410 816.000 1813.690 820.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1830.890 816.000 1831.170 820.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1847.910 816.000 1848.190 820.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1865.390 816.000 1865.670 820.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1882.870 816.000 1883.150 820.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1899.890 816.000 1900.170 820.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 816.000 183.910 820.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1917.370 816.000 1917.650 820.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1934.850 816.000 1935.130 820.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1951.870 816.000 1952.150 820.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1969.350 816.000 1969.630 820.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1986.830 816.000 1987.110 820.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2004.310 816.000 2004.590 820.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2021.330 816.000 2021.610 820.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2038.810 816.000 2039.090 820.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2056.290 816.000 2056.570 820.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2073.310 816.000 2073.590 820.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 816.000 201.390 820.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2090.790 816.000 2091.070 820.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2108.270 816.000 2108.550 820.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2125.290 816.000 2125.570 820.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2142.770 816.000 2143.050 820.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2160.250 816.000 2160.530 820.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2177.270 816.000 2177.550 820.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2194.750 816.000 2195.030 820.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2212.230 816.000 2212.510 820.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 816.000 218.870 820.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 816.000 235.890 820.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 816.000 253.370 820.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 816.000 270.850 820.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 816.000 287.870 820.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 816.000 305.350 820.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 816.000 322.830 820.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 816.000 339.850 820.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 816.000 27.970 820.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 816.000 357.330 820.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 816.000 374.810 820.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 816.000 391.830 820.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 816.000 409.310 820.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.510 816.000 426.790 820.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 816.000 444.270 820.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 816.000 461.290 820.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.490 816.000 478.770 820.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 816.000 496.250 820.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 816.000 513.270 820.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 816.000 45.450 820.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.470 816.000 530.750 820.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.950 816.000 548.230 820.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.970 816.000 565.250 820.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.450 816.000 582.730 820.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.930 816.000 600.210 820.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.950 816.000 617.230 820.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 816.000 634.710 820.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.910 816.000 652.190 820.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.390 816.000 669.670 820.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.410 816.000 686.690 820.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 816.000 62.470 820.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.890 816.000 704.170 820.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 816.000 721.650 820.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.390 816.000 738.670 820.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.870 816.000 756.150 820.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.350 816.000 773.630 820.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.370 816.000 790.650 820.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.850 816.000 808.130 820.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 825.330 816.000 825.610 820.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 842.350 816.000 842.630 820.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.830 816.000 860.110 820.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 816.000 79.950 820.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.310 816.000 877.590 820.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.330 816.000 894.610 820.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.810 816.000 912.090 820.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.290 816.000 929.570 820.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.770 816.000 947.050 820.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.790 816.000 964.070 820.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 981.270 816.000 981.550 820.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.750 816.000 999.030 820.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1015.770 816.000 1016.050 820.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.250 816.000 1033.530 820.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 816.000 97.430 820.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1050.730 816.000 1051.010 820.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1067.750 816.000 1068.030 820.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.230 816.000 1085.510 820.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.710 816.000 1102.990 820.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1119.730 816.000 1120.010 820.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.210 816.000 1137.490 820.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1154.690 816.000 1154.970 820.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1171.710 816.000 1171.990 820.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1189.190 816.000 1189.470 820.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1206.670 816.000 1206.950 820.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 816.000 114.450 820.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1224.150 816.000 1224.430 820.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1241.170 816.000 1241.450 820.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1258.650 816.000 1258.930 820.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1276.130 816.000 1276.410 820.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1293.150 816.000 1293.430 820.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1310.630 816.000 1310.910 820.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1328.110 816.000 1328.390 820.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1345.130 816.000 1345.410 820.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.610 816.000 1362.890 820.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1380.090 816.000 1380.370 820.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 816.000 131.930 820.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.110 816.000 1397.390 820.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1414.590 816.000 1414.870 820.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.070 816.000 1432.350 820.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1449.090 816.000 1449.370 820.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1466.570 816.000 1466.850 820.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.050 816.000 1484.330 820.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1501.530 816.000 1501.810 820.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1518.550 816.000 1518.830 820.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1536.030 816.000 1536.310 820.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1553.510 816.000 1553.790 820.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 816.000 149.410 820.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1570.530 816.000 1570.810 820.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1588.010 816.000 1588.290 820.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1605.490 816.000 1605.770 820.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1622.510 816.000 1622.790 820.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.990 816.000 1640.270 820.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1657.470 816.000 1657.750 820.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1674.490 816.000 1674.770 820.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1691.970 816.000 1692.250 820.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1709.450 816.000 1709.730 820.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1726.930 816.000 1727.210 820.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 816.000 166.890 820.000 ;
    END
  END la_oenb[9]
  PIN la_output[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 816.000 15.090 820.000 ;
    END
  END la_output[0]
  PIN la_output[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1748.550 816.000 1748.830 820.000 ;
    END
  END la_output[100]
  PIN la_output[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1765.570 816.000 1765.850 820.000 ;
    END
  END la_output[101]
  PIN la_output[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1783.050 816.000 1783.330 820.000 ;
    END
  END la_output[102]
  PIN la_output[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1800.530 816.000 1800.810 820.000 ;
    END
  END la_output[103]
  PIN la_output[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1817.550 816.000 1817.830 820.000 ;
    END
  END la_output[104]
  PIN la_output[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1835.030 816.000 1835.310 820.000 ;
    END
  END la_output[105]
  PIN la_output[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1852.510 816.000 1852.790 820.000 ;
    END
  END la_output[106]
  PIN la_output[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1869.530 816.000 1869.810 820.000 ;
    END
  END la_output[107]
  PIN la_output[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1887.010 816.000 1887.290 820.000 ;
    END
  END la_output[108]
  PIN la_output[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1904.490 816.000 1904.770 820.000 ;
    END
  END la_output[109]
  PIN la_output[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 816.000 188.510 820.000 ;
    END
  END la_output[10]
  PIN la_output[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1921.970 816.000 1922.250 820.000 ;
    END
  END la_output[110]
  PIN la_output[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1938.990 816.000 1939.270 820.000 ;
    END
  END la_output[111]
  PIN la_output[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1956.470 816.000 1956.750 820.000 ;
    END
  END la_output[112]
  PIN la_output[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1973.950 816.000 1974.230 820.000 ;
    END
  END la_output[113]
  PIN la_output[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1990.970 816.000 1991.250 820.000 ;
    END
  END la_output[114]
  PIN la_output[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2008.450 816.000 2008.730 820.000 ;
    END
  END la_output[115]
  PIN la_output[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2025.930 816.000 2026.210 820.000 ;
    END
  END la_output[116]
  PIN la_output[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2042.950 816.000 2043.230 820.000 ;
    END
  END la_output[117]
  PIN la_output[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2060.430 816.000 2060.710 820.000 ;
    END
  END la_output[118]
  PIN la_output[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2077.910 816.000 2078.190 820.000 ;
    END
  END la_output[119]
  PIN la_output[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 816.000 205.530 820.000 ;
    END
  END la_output[11]
  PIN la_output[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2094.930 816.000 2095.210 820.000 ;
    END
  END la_output[120]
  PIN la_output[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2112.410 816.000 2112.690 820.000 ;
    END
  END la_output[121]
  PIN la_output[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2129.890 816.000 2130.170 820.000 ;
    END
  END la_output[122]
  PIN la_output[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2146.910 816.000 2147.190 820.000 ;
    END
  END la_output[123]
  PIN la_output[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2164.390 816.000 2164.670 820.000 ;
    END
  END la_output[124]
  PIN la_output[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2181.870 816.000 2182.150 820.000 ;
    END
  END la_output[125]
  PIN la_output[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2199.350 816.000 2199.630 820.000 ;
    END
  END la_output[126]
  PIN la_output[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2216.370 816.000 2216.650 820.000 ;
    END
  END la_output[127]
  PIN la_output[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 816.000 223.010 820.000 ;
    END
  END la_output[12]
  PIN la_output[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 816.000 240.490 820.000 ;
    END
  END la_output[13]
  PIN la_output[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 816.000 257.510 820.000 ;
    END
  END la_output[14]
  PIN la_output[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 816.000 274.990 820.000 ;
    END
  END la_output[15]
  PIN la_output[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 816.000 292.470 820.000 ;
    END
  END la_output[16]
  PIN la_output[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 816.000 309.490 820.000 ;
    END
  END la_output[17]
  PIN la_output[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 816.000 326.970 820.000 ;
    END
  END la_output[18]
  PIN la_output[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 816.000 344.450 820.000 ;
    END
  END la_output[19]
  PIN la_output[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 816.000 32.110 820.000 ;
    END
  END la_output[1]
  PIN la_output[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 816.000 361.930 820.000 ;
    END
  END la_output[20]
  PIN la_output[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.670 816.000 378.950 820.000 ;
    END
  END la_output[21]
  PIN la_output[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 816.000 396.430 820.000 ;
    END
  END la_output[22]
  PIN la_output[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.630 816.000 413.910 820.000 ;
    END
  END la_output[23]
  PIN la_output[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.650 816.000 430.930 820.000 ;
    END
  END la_output[24]
  PIN la_output[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.130 816.000 448.410 820.000 ;
    END
  END la_output[25]
  PIN la_output[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 816.000 465.890 820.000 ;
    END
  END la_output[26]
  PIN la_output[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.630 816.000 482.910 820.000 ;
    END
  END la_output[27]
  PIN la_output[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.110 816.000 500.390 820.000 ;
    END
  END la_output[28]
  PIN la_output[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.590 816.000 517.870 820.000 ;
    END
  END la_output[29]
  PIN la_output[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 816.000 49.590 820.000 ;
    END
  END la_output[2]
  PIN la_output[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 816.000 534.890 820.000 ;
    END
  END la_output[30]
  PIN la_output[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.090 816.000 552.370 820.000 ;
    END
  END la_output[31]
  PIN la_output[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 816.000 569.850 820.000 ;
    END
  END la_output[32]
  PIN la_output[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 816.000 586.870 820.000 ;
    END
  END la_output[33]
  PIN la_output[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.070 816.000 604.350 820.000 ;
    END
  END la_output[34]
  PIN la_output[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 816.000 621.830 820.000 ;
    END
  END la_output[35]
  PIN la_output[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.030 816.000 639.310 820.000 ;
    END
  END la_output[36]
  PIN la_output[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.050 816.000 656.330 820.000 ;
    END
  END la_output[37]
  PIN la_output[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.530 816.000 673.810 820.000 ;
    END
  END la_output[38]
  PIN la_output[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.010 816.000 691.290 820.000 ;
    END
  END la_output[39]
  PIN la_output[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 816.000 67.070 820.000 ;
    END
  END la_output[3]
  PIN la_output[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.030 816.000 708.310 820.000 ;
    END
  END la_output[40]
  PIN la_output[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.510 816.000 725.790 820.000 ;
    END
  END la_output[41]
  PIN la_output[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.990 816.000 743.270 820.000 ;
    END
  END la_output[42]
  PIN la_output[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 816.000 760.290 820.000 ;
    END
  END la_output[43]
  PIN la_output[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.490 816.000 777.770 820.000 ;
    END
  END la_output[44]
  PIN la_output[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.970 816.000 795.250 820.000 ;
    END
  END la_output[45]
  PIN la_output[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.990 816.000 812.270 820.000 ;
    END
  END la_output[46]
  PIN la_output[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.470 816.000 829.750 820.000 ;
    END
  END la_output[47]
  PIN la_output[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.950 816.000 847.230 820.000 ;
    END
  END la_output[48]
  PIN la_output[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.430 816.000 864.710 820.000 ;
    END
  END la_output[49]
  PIN la_output[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 816.000 84.550 820.000 ;
    END
  END la_output[4]
  PIN la_output[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.450 816.000 881.730 820.000 ;
    END
  END la_output[50]
  PIN la_output[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.930 816.000 899.210 820.000 ;
    END
  END la_output[51]
  PIN la_output[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 916.410 816.000 916.690 820.000 ;
    END
  END la_output[52]
  PIN la_output[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.430 816.000 933.710 820.000 ;
    END
  END la_output[53]
  PIN la_output[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 950.910 816.000 951.190 820.000 ;
    END
  END la_output[54]
  PIN la_output[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 968.390 816.000 968.670 820.000 ;
    END
  END la_output[55]
  PIN la_output[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.410 816.000 985.690 820.000 ;
    END
  END la_output[56]
  PIN la_output[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1002.890 816.000 1003.170 820.000 ;
    END
  END la_output[57]
  PIN la_output[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.370 816.000 1020.650 820.000 ;
    END
  END la_output[58]
  PIN la_output[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.390 816.000 1037.670 820.000 ;
    END
  END la_output[59]
  PIN la_output[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 816.000 101.570 820.000 ;
    END
  END la_output[5]
  PIN la_output[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.870 816.000 1055.150 820.000 ;
    END
  END la_output[60]
  PIN la_output[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 816.000 1072.630 820.000 ;
    END
  END la_output[61]
  PIN la_output[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1089.370 816.000 1089.650 820.000 ;
    END
  END la_output[62]
  PIN la_output[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1106.850 816.000 1107.130 820.000 ;
    END
  END la_output[63]
  PIN la_output[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1124.330 816.000 1124.610 820.000 ;
    END
  END la_output[64]
  PIN la_output[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1141.810 816.000 1142.090 820.000 ;
    END
  END la_output[65]
  PIN la_output[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1158.830 816.000 1159.110 820.000 ;
    END
  END la_output[66]
  PIN la_output[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1176.310 816.000 1176.590 820.000 ;
    END
  END la_output[67]
  PIN la_output[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1193.790 816.000 1194.070 820.000 ;
    END
  END la_output[68]
  PIN la_output[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1210.810 816.000 1211.090 820.000 ;
    END
  END la_output[69]
  PIN la_output[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 816.000 119.050 820.000 ;
    END
  END la_output[6]
  PIN la_output[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1228.290 816.000 1228.570 820.000 ;
    END
  END la_output[70]
  PIN la_output[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1245.770 816.000 1246.050 820.000 ;
    END
  END la_output[71]
  PIN la_output[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1262.790 816.000 1263.070 820.000 ;
    END
  END la_output[72]
  PIN la_output[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1280.270 816.000 1280.550 820.000 ;
    END
  END la_output[73]
  PIN la_output[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.750 816.000 1298.030 820.000 ;
    END
  END la_output[74]
  PIN la_output[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1314.770 816.000 1315.050 820.000 ;
    END
  END la_output[75]
  PIN la_output[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1332.250 816.000 1332.530 820.000 ;
    END
  END la_output[76]
  PIN la_output[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1349.730 816.000 1350.010 820.000 ;
    END
  END la_output[77]
  PIN la_output[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1366.750 816.000 1367.030 820.000 ;
    END
  END la_output[78]
  PIN la_output[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1384.230 816.000 1384.510 820.000 ;
    END
  END la_output[79]
  PIN la_output[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 816.000 136.530 820.000 ;
    END
  END la_output[7]
  PIN la_output[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1401.710 816.000 1401.990 820.000 ;
    END
  END la_output[80]
  PIN la_output[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1419.190 816.000 1419.470 820.000 ;
    END
  END la_output[81]
  PIN la_output[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1436.210 816.000 1436.490 820.000 ;
    END
  END la_output[82]
  PIN la_output[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1453.690 816.000 1453.970 820.000 ;
    END
  END la_output[83]
  PIN la_output[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.170 816.000 1471.450 820.000 ;
    END
  END la_output[84]
  PIN la_output[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1488.190 816.000 1488.470 820.000 ;
    END
  END la_output[85]
  PIN la_output[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1505.670 816.000 1505.950 820.000 ;
    END
  END la_output[86]
  PIN la_output[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1523.150 816.000 1523.430 820.000 ;
    END
  END la_output[87]
  PIN la_output[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1540.170 816.000 1540.450 820.000 ;
    END
  END la_output[88]
  PIN la_output[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1557.650 816.000 1557.930 820.000 ;
    END
  END la_output[89]
  PIN la_output[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 816.000 153.550 820.000 ;
    END
  END la_output[8]
  PIN la_output[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1575.130 816.000 1575.410 820.000 ;
    END
  END la_output[90]
  PIN la_output[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1592.150 816.000 1592.430 820.000 ;
    END
  END la_output[91]
  PIN la_output[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1609.630 816.000 1609.910 820.000 ;
    END
  END la_output[92]
  PIN la_output[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1627.110 816.000 1627.390 820.000 ;
    END
  END la_output[93]
  PIN la_output[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1644.130 816.000 1644.410 820.000 ;
    END
  END la_output[94]
  PIN la_output[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.610 816.000 1661.890 820.000 ;
    END
  END la_output[95]
  PIN la_output[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1679.090 816.000 1679.370 820.000 ;
    END
  END la_output[96]
  PIN la_output[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1696.570 816.000 1696.850 820.000 ;
    END
  END la_output[97]
  PIN la_output[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1713.590 816.000 1713.870 820.000 ;
    END
  END la_output[98]
  PIN la_output[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1731.070 816.000 1731.350 820.000 ;
    END
  END la_output[99]
  PIN la_output[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 816.000 171.030 820.000 ;
    END
  END la_output[9]
  PIN mprj_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2220.970 816.000 2221.250 820.000 ;
    END
  END mprj_ack_i
  PIN mprj_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2242.590 816.000 2242.870 820.000 ;
    END
  END mprj_adr_o[0]
  PIN mprj_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2389.790 816.000 2390.070 820.000 ;
    END
  END mprj_adr_o[10]
  PIN mprj_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2402.670 816.000 2402.950 820.000 ;
    END
  END mprj_adr_o[11]
  PIN mprj_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2416.010 816.000 2416.290 820.000 ;
    END
  END mprj_adr_o[12]
  PIN mprj_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2428.890 816.000 2429.170 820.000 ;
    END
  END mprj_adr_o[13]
  PIN mprj_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2441.770 816.000 2442.050 820.000 ;
    END
  END mprj_adr_o[14]
  PIN mprj_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2454.650 816.000 2454.930 820.000 ;
    END
  END mprj_adr_o[15]
  PIN mprj_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2467.990 816.000 2468.270 820.000 ;
    END
  END mprj_adr_o[16]
  PIN mprj_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2480.870 816.000 2481.150 820.000 ;
    END
  END mprj_adr_o[17]
  PIN mprj_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2493.750 816.000 2494.030 820.000 ;
    END
  END mprj_adr_o[18]
  PIN mprj_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2507.090 816.000 2507.370 820.000 ;
    END
  END mprj_adr_o[19]
  PIN mprj_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2259.610 816.000 2259.890 820.000 ;
    END
  END mprj_adr_o[1]
  PIN mprj_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2519.970 816.000 2520.250 820.000 ;
    END
  END mprj_adr_o[20]
  PIN mprj_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2532.850 816.000 2533.130 820.000 ;
    END
  END mprj_adr_o[21]
  PIN mprj_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2545.730 816.000 2546.010 820.000 ;
    END
  END mprj_adr_o[22]
  PIN mprj_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2559.070 816.000 2559.350 820.000 ;
    END
  END mprj_adr_o[23]
  PIN mprj_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2571.950 816.000 2572.230 820.000 ;
    END
  END mprj_adr_o[24]
  PIN mprj_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2584.830 816.000 2585.110 820.000 ;
    END
  END mprj_adr_o[25]
  PIN mprj_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2597.710 816.000 2597.990 820.000 ;
    END
  END mprj_adr_o[26]
  PIN mprj_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2611.050 816.000 2611.330 820.000 ;
    END
  END mprj_adr_o[27]
  PIN mprj_adr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2623.930 816.000 2624.210 820.000 ;
    END
  END mprj_adr_o[28]
  PIN mprj_adr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2636.810 816.000 2637.090 820.000 ;
    END
  END mprj_adr_o[29]
  PIN mprj_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2277.090 816.000 2277.370 820.000 ;
    END
  END mprj_adr_o[2]
  PIN mprj_adr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2649.690 816.000 2649.970 820.000 ;
    END
  END mprj_adr_o[30]
  PIN mprj_adr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2663.030 816.000 2663.310 820.000 ;
    END
  END mprj_adr_o[31]
  PIN mprj_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2294.570 816.000 2294.850 820.000 ;
    END
  END mprj_adr_o[3]
  PIN mprj_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2312.050 816.000 2312.330 820.000 ;
    END
  END mprj_adr_o[4]
  PIN mprj_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2324.930 816.000 2325.210 820.000 ;
    END
  END mprj_adr_o[5]
  PIN mprj_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2337.810 816.000 2338.090 820.000 ;
    END
  END mprj_adr_o[6]
  PIN mprj_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2350.690 816.000 2350.970 820.000 ;
    END
  END mprj_adr_o[7]
  PIN mprj_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2364.030 816.000 2364.310 820.000 ;
    END
  END mprj_adr_o[8]
  PIN mprj_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2376.910 816.000 2377.190 820.000 ;
    END
  END mprj_adr_o[9]
  PIN mprj_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2225.110 816.000 2225.390 820.000 ;
    END
  END mprj_cyc_o
  PIN mprj_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2246.730 816.000 2247.010 820.000 ;
    END
  END mprj_dat_i[0]
  PIN mprj_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2394.390 816.000 2394.670 820.000 ;
    END
  END mprj_dat_i[10]
  PIN mprj_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2407.270 816.000 2407.550 820.000 ;
    END
  END mprj_dat_i[11]
  PIN mprj_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2420.150 816.000 2420.430 820.000 ;
    END
  END mprj_dat_i[12]
  PIN mprj_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2433.030 816.000 2433.310 820.000 ;
    END
  END mprj_dat_i[13]
  PIN mprj_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2446.370 816.000 2446.650 820.000 ;
    END
  END mprj_dat_i[14]
  PIN mprj_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2459.250 816.000 2459.530 820.000 ;
    END
  END mprj_dat_i[15]
  PIN mprj_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2472.130 816.000 2472.410 820.000 ;
    END
  END mprj_dat_i[16]
  PIN mprj_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2485.010 816.000 2485.290 820.000 ;
    END
  END mprj_dat_i[17]
  PIN mprj_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2498.350 816.000 2498.630 820.000 ;
    END
  END mprj_dat_i[18]
  PIN mprj_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2511.230 816.000 2511.510 820.000 ;
    END
  END mprj_dat_i[19]
  PIN mprj_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2264.210 816.000 2264.490 820.000 ;
    END
  END mprj_dat_i[1]
  PIN mprj_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2524.110 816.000 2524.390 820.000 ;
    END
  END mprj_dat_i[20]
  PIN mprj_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2536.990 816.000 2537.270 820.000 ;
    END
  END mprj_dat_i[21]
  PIN mprj_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2550.330 816.000 2550.610 820.000 ;
    END
  END mprj_dat_i[22]
  PIN mprj_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2563.210 816.000 2563.490 820.000 ;
    END
  END mprj_dat_i[23]
  PIN mprj_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2576.090 816.000 2576.370 820.000 ;
    END
  END mprj_dat_i[24]
  PIN mprj_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2589.430 816.000 2589.710 820.000 ;
    END
  END mprj_dat_i[25]
  PIN mprj_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2602.310 816.000 2602.590 820.000 ;
    END
  END mprj_dat_i[26]
  PIN mprj_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2615.190 816.000 2615.470 820.000 ;
    END
  END mprj_dat_i[27]
  PIN mprj_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2628.070 816.000 2628.350 820.000 ;
    END
  END mprj_dat_i[28]
  PIN mprj_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2641.410 816.000 2641.690 820.000 ;
    END
  END mprj_dat_i[29]
  PIN mprj_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2281.690 816.000 2281.970 820.000 ;
    END
  END mprj_dat_i[2]
  PIN mprj_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2654.290 816.000 2654.570 820.000 ;
    END
  END mprj_dat_i[30]
  PIN mprj_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2667.170 816.000 2667.450 820.000 ;
    END
  END mprj_dat_i[31]
  PIN mprj_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2298.710 816.000 2298.990 820.000 ;
    END
  END mprj_dat_i[3]
  PIN mprj_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2316.190 816.000 2316.470 820.000 ;
    END
  END mprj_dat_i[4]
  PIN mprj_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2329.070 816.000 2329.350 820.000 ;
    END
  END mprj_dat_i[5]
  PIN mprj_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2341.950 816.000 2342.230 820.000 ;
    END
  END mprj_dat_i[6]
  PIN mprj_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2355.290 816.000 2355.570 820.000 ;
    END
  END mprj_dat_i[7]
  PIN mprj_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2368.170 816.000 2368.450 820.000 ;
    END
  END mprj_dat_i[8]
  PIN mprj_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2381.050 816.000 2381.330 820.000 ;
    END
  END mprj_dat_i[9]
  PIN mprj_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2251.330 816.000 2251.610 820.000 ;
    END
  END mprj_dat_o[0]
  PIN mprj_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2398.530 816.000 2398.810 820.000 ;
    END
  END mprj_dat_o[10]
  PIN mprj_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2411.410 816.000 2411.690 820.000 ;
    END
  END mprj_dat_o[11]
  PIN mprj_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2424.290 816.000 2424.570 820.000 ;
    END
  END mprj_dat_o[12]
  PIN mprj_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2437.630 816.000 2437.910 820.000 ;
    END
  END mprj_dat_o[13]
  PIN mprj_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2450.510 816.000 2450.790 820.000 ;
    END
  END mprj_dat_o[14]
  PIN mprj_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2463.390 816.000 2463.670 820.000 ;
    END
  END mprj_dat_o[15]
  PIN mprj_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2476.730 816.000 2477.010 820.000 ;
    END
  END mprj_dat_o[16]
  PIN mprj_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2489.610 816.000 2489.890 820.000 ;
    END
  END mprj_dat_o[17]
  PIN mprj_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2502.490 816.000 2502.770 820.000 ;
    END
  END mprj_dat_o[18]
  PIN mprj_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2515.370 816.000 2515.650 820.000 ;
    END
  END mprj_dat_o[19]
  PIN mprj_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2268.350 816.000 2268.630 820.000 ;
    END
  END mprj_dat_o[1]
  PIN mprj_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2528.710 816.000 2528.990 820.000 ;
    END
  END mprj_dat_o[20]
  PIN mprj_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2541.590 816.000 2541.870 820.000 ;
    END
  END mprj_dat_o[21]
  PIN mprj_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2554.470 816.000 2554.750 820.000 ;
    END
  END mprj_dat_o[22]
  PIN mprj_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2567.350 816.000 2567.630 820.000 ;
    END
  END mprj_dat_o[23]
  PIN mprj_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2580.690 816.000 2580.970 820.000 ;
    END
  END mprj_dat_o[24]
  PIN mprj_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2593.570 816.000 2593.850 820.000 ;
    END
  END mprj_dat_o[25]
  PIN mprj_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2606.450 816.000 2606.730 820.000 ;
    END
  END mprj_dat_o[26]
  PIN mprj_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2619.330 816.000 2619.610 820.000 ;
    END
  END mprj_dat_o[27]
  PIN mprj_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2632.670 816.000 2632.950 820.000 ;
    END
  END mprj_dat_o[28]
  PIN mprj_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2645.550 816.000 2645.830 820.000 ;
    END
  END mprj_dat_o[29]
  PIN mprj_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2285.830 816.000 2286.110 820.000 ;
    END
  END mprj_dat_o[2]
  PIN mprj_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2658.430 816.000 2658.710 820.000 ;
    END
  END mprj_dat_o[30]
  PIN mprj_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2671.770 816.000 2672.050 820.000 ;
    END
  END mprj_dat_o[31]
  PIN mprj_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2303.310 816.000 2303.590 820.000 ;
    END
  END mprj_dat_o[3]
  PIN mprj_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2320.330 816.000 2320.610 820.000 ;
    END
  END mprj_dat_o[4]
  PIN mprj_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2333.670 816.000 2333.950 820.000 ;
    END
  END mprj_dat_o[5]
  PIN mprj_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2346.550 816.000 2346.830 820.000 ;
    END
  END mprj_dat_o[6]
  PIN mprj_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2359.430 816.000 2359.710 820.000 ;
    END
  END mprj_dat_o[7]
  PIN mprj_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2372.310 816.000 2372.590 820.000 ;
    END
  END mprj_dat_o[8]
  PIN mprj_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2385.650 816.000 2385.930 820.000 ;
    END
  END mprj_dat_o[9]
  PIN mprj_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2255.470 816.000 2255.750 820.000 ;
    END
  END mprj_sel_o[0]
  PIN mprj_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2272.950 816.000 2273.230 820.000 ;
    END
  END mprj_sel_o[1]
  PIN mprj_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2289.970 816.000 2290.250 820.000 ;
    END
  END mprj_sel_o[2]
  PIN mprj_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2307.450 816.000 2307.730 820.000 ;
    END
  END mprj_sel_o[3]
  PIN mprj_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2229.250 816.000 2229.530 820.000 ;
    END
  END mprj_stb_o
  PIN mprj_wb_iena
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2233.850 816.000 2234.130 820.000 ;
    END
  END mprj_wb_iena
  PIN mprj_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2237.990 816.000 2238.270 820.000 ;
    END
  END mprj_we_o
  PIN qspi_enabled
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 450.880 2700.000 451.480 ;
    END
  END qspi_enabled
  PIN ser_rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 420.960 2700.000 421.560 ;
    END
  END ser_rx
  PIN ser_tx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 428.440 2700.000 429.040 ;
    END
  END ser_tx
  PIN spi_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 405.320 2700.000 405.920 ;
    END
  END spi_csb
  PIN spi_enabled
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 435.920 2700.000 436.520 ;
    END
  END spi_enabled
  PIN spi_sck
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 397.840 2700.000 398.440 ;
    END
  END spi_sck
  PIN spi_sdi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 413.480 2700.000 414.080 ;
    END
  END spi_sdi
  PIN spi_sdo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 390.360 2700.000 390.960 ;
    END
  END spi_sdo
  PIN spi_sdoenb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 382.880 2700.000 383.480 ;
    END
  END spi_sdoenb
  PIN sram_ro_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 10.920 2700.000 11.520 ;
    END
  END sram_ro_addr[0]
  PIN sram_ro_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 18.400 2700.000 19.000 ;
    END
  END sram_ro_addr[1]
  PIN sram_ro_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 25.880 2700.000 26.480 ;
    END
  END sram_ro_addr[2]
  PIN sram_ro_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 33.360 2700.000 33.960 ;
    END
  END sram_ro_addr[3]
  PIN sram_ro_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 40.840 2700.000 41.440 ;
    END
  END sram_ro_addr[4]
  PIN sram_ro_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 49.000 2700.000 49.600 ;
    END
  END sram_ro_addr[5]
  PIN sram_ro_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 56.480 2700.000 57.080 ;
    END
  END sram_ro_addr[6]
  PIN sram_ro_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 63.960 2700.000 64.560 ;
    END
  END sram_ro_addr[7]
  PIN sram_ro_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 71.440 2700.000 72.040 ;
    END
  END sram_ro_clk
  PIN sram_ro_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 3.440 2700.000 4.040 ;
    END
  END sram_ro_csb
  PIN sram_ro_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 78.920 2700.000 79.520 ;
    END
  END sram_ro_data[0]
  PIN sram_ro_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 155.080 2700.000 155.680 ;
    END
  END sram_ro_data[10]
  PIN sram_ro_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 162.560 2700.000 163.160 ;
    END
  END sram_ro_data[11]
  PIN sram_ro_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 170.040 2700.000 170.640 ;
    END
  END sram_ro_data[12]
  PIN sram_ro_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 177.520 2700.000 178.120 ;
    END
  END sram_ro_data[13]
  PIN sram_ro_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 185.680 2700.000 186.280 ;
    END
  END sram_ro_data[14]
  PIN sram_ro_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 193.160 2700.000 193.760 ;
    END
  END sram_ro_data[15]
  PIN sram_ro_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 200.640 2700.000 201.240 ;
    END
  END sram_ro_data[16]
  PIN sram_ro_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 208.120 2700.000 208.720 ;
    END
  END sram_ro_data[17]
  PIN sram_ro_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 215.600 2700.000 216.200 ;
    END
  END sram_ro_data[18]
  PIN sram_ro_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 223.080 2700.000 223.680 ;
    END
  END sram_ro_data[19]
  PIN sram_ro_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 86.400 2700.000 87.000 ;
    END
  END sram_ro_data[1]
  PIN sram_ro_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 231.240 2700.000 231.840 ;
    END
  END sram_ro_data[20]
  PIN sram_ro_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 238.720 2700.000 239.320 ;
    END
  END sram_ro_data[21]
  PIN sram_ro_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 246.200 2700.000 246.800 ;
    END
  END sram_ro_data[22]
  PIN sram_ro_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 253.680 2700.000 254.280 ;
    END
  END sram_ro_data[23]
  PIN sram_ro_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 261.160 2700.000 261.760 ;
    END
  END sram_ro_data[24]
  PIN sram_ro_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 268.640 2700.000 269.240 ;
    END
  END sram_ro_data[25]
  PIN sram_ro_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 276.800 2700.000 277.400 ;
    END
  END sram_ro_data[26]
  PIN sram_ro_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 284.280 2700.000 284.880 ;
    END
  END sram_ro_data[27]
  PIN sram_ro_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 291.760 2700.000 292.360 ;
    END
  END sram_ro_data[28]
  PIN sram_ro_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 299.240 2700.000 299.840 ;
    END
  END sram_ro_data[29]
  PIN sram_ro_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 94.560 2700.000 95.160 ;
    END
  END sram_ro_data[2]
  PIN sram_ro_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 306.720 2700.000 307.320 ;
    END
  END sram_ro_data[30]
  PIN sram_ro_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 314.200 2700.000 314.800 ;
    END
  END sram_ro_data[31]
  PIN sram_ro_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 102.040 2700.000 102.640 ;
    END
  END sram_ro_data[3]
  PIN sram_ro_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 109.520 2700.000 110.120 ;
    END
  END sram_ro_data[4]
  PIN sram_ro_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 117.000 2700.000 117.600 ;
    END
  END sram_ro_data[5]
  PIN sram_ro_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 124.480 2700.000 125.080 ;
    END
  END sram_ro_data[6]
  PIN sram_ro_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 131.960 2700.000 132.560 ;
    END
  END sram_ro_data[7]
  PIN sram_ro_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 140.120 2700.000 140.720 ;
    END
  END sram_ro_data[8]
  PIN sram_ro_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 147.600 2700.000 148.200 ;
    END
  END sram_ro_data[9]
  PIN trap
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 352.280 2700.000 352.880 ;
    END
  END trap
  PIN uart_enabled
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2696.000 443.400 2700.000 444.000 ;
    END
  END uart_enabled
  PIN user_irq_ena[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2675.910 816.000 2676.190 820.000 ;
    END
  END user_irq_ena[0]
  PIN user_irq_ena[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2680.050 816.000 2680.330 820.000 ;
    END
  END user_irq_ena[1]
  PIN user_irq_ena[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2684.650 816.000 2684.930 820.000 ;
    END
  END user_irq_ena[2]
  OBS
      LAYER li1 ;
        RECT 29.345 23.205 2697.755 819.655 ;
      LAYER met1 ;
        RECT 1.910 6.500 2697.830 819.980 ;
      LAYER met2 ;
        RECT 2.490 815.720 5.790 819.730 ;
        RECT 6.630 815.720 9.930 819.730 ;
        RECT 10.770 815.720 14.530 819.730 ;
        RECT 15.370 815.720 18.670 819.730 ;
        RECT 19.510 815.720 23.270 819.730 ;
        RECT 24.110 815.720 27.410 819.730 ;
        RECT 28.250 815.720 31.550 819.730 ;
        RECT 32.390 815.720 36.150 819.730 ;
        RECT 36.990 815.720 40.290 819.730 ;
        RECT 41.130 815.720 44.890 819.730 ;
        RECT 45.730 815.720 49.030 819.730 ;
        RECT 49.870 815.720 53.630 819.730 ;
        RECT 54.470 815.720 57.770 819.730 ;
        RECT 58.610 815.720 61.910 819.730 ;
        RECT 62.750 815.720 66.510 819.730 ;
        RECT 67.350 815.720 70.650 819.730 ;
        RECT 71.490 815.720 75.250 819.730 ;
        RECT 76.090 815.720 79.390 819.730 ;
        RECT 80.230 815.720 83.990 819.730 ;
        RECT 84.830 815.720 88.130 819.730 ;
        RECT 88.970 815.720 92.270 819.730 ;
        RECT 93.110 815.720 96.870 819.730 ;
        RECT 97.710 815.720 101.010 819.730 ;
        RECT 101.850 815.720 105.610 819.730 ;
        RECT 106.450 815.720 109.750 819.730 ;
        RECT 110.590 815.720 113.890 819.730 ;
        RECT 114.730 815.720 118.490 819.730 ;
        RECT 119.330 815.720 122.630 819.730 ;
        RECT 123.470 815.720 127.230 819.730 ;
        RECT 128.070 815.720 131.370 819.730 ;
        RECT 132.210 815.720 135.970 819.730 ;
        RECT 136.810 815.720 140.110 819.730 ;
        RECT 140.950 815.720 144.250 819.730 ;
        RECT 145.090 815.720 148.850 819.730 ;
        RECT 149.690 815.720 152.990 819.730 ;
        RECT 153.830 815.720 157.590 819.730 ;
        RECT 158.430 815.720 161.730 819.730 ;
        RECT 162.570 815.720 166.330 819.730 ;
        RECT 167.170 815.720 170.470 819.730 ;
        RECT 171.310 815.720 174.610 819.730 ;
        RECT 175.450 815.720 179.210 819.730 ;
        RECT 180.050 815.720 183.350 819.730 ;
        RECT 184.190 815.720 187.950 819.730 ;
        RECT 188.790 815.720 192.090 819.730 ;
        RECT 192.930 815.720 196.230 819.730 ;
        RECT 197.070 815.720 200.830 819.730 ;
        RECT 201.670 815.720 204.970 819.730 ;
        RECT 205.810 815.720 209.570 819.730 ;
        RECT 210.410 815.720 213.710 819.730 ;
        RECT 214.550 815.720 218.310 819.730 ;
        RECT 219.150 815.720 222.450 819.730 ;
        RECT 223.290 815.720 226.590 819.730 ;
        RECT 227.430 815.720 231.190 819.730 ;
        RECT 232.030 815.720 235.330 819.730 ;
        RECT 236.170 815.720 239.930 819.730 ;
        RECT 240.770 815.720 244.070 819.730 ;
        RECT 244.910 815.720 248.670 819.730 ;
        RECT 249.510 815.720 252.810 819.730 ;
        RECT 253.650 815.720 256.950 819.730 ;
        RECT 257.790 815.720 261.550 819.730 ;
        RECT 262.390 815.720 265.690 819.730 ;
        RECT 266.530 815.720 270.290 819.730 ;
        RECT 271.130 815.720 274.430 819.730 ;
        RECT 275.270 815.720 279.030 819.730 ;
        RECT 279.870 815.720 283.170 819.730 ;
        RECT 284.010 815.720 287.310 819.730 ;
        RECT 288.150 815.720 291.910 819.730 ;
        RECT 292.750 815.720 296.050 819.730 ;
        RECT 296.890 815.720 300.650 819.730 ;
        RECT 301.490 815.720 304.790 819.730 ;
        RECT 305.630 815.720 308.930 819.730 ;
        RECT 309.770 815.720 313.530 819.730 ;
        RECT 314.370 815.720 317.670 819.730 ;
        RECT 318.510 815.720 322.270 819.730 ;
        RECT 323.110 815.720 326.410 819.730 ;
        RECT 327.250 815.720 331.010 819.730 ;
        RECT 331.850 815.720 335.150 819.730 ;
        RECT 335.990 815.720 339.290 819.730 ;
        RECT 340.130 815.720 343.890 819.730 ;
        RECT 344.730 815.720 348.030 819.730 ;
        RECT 348.870 815.720 352.630 819.730 ;
        RECT 353.470 815.720 356.770 819.730 ;
        RECT 357.610 815.720 361.370 819.730 ;
        RECT 362.210 815.720 365.510 819.730 ;
        RECT 366.350 815.720 369.650 819.730 ;
        RECT 370.490 815.720 374.250 819.730 ;
        RECT 375.090 815.720 378.390 819.730 ;
        RECT 379.230 815.720 382.990 819.730 ;
        RECT 383.830 815.720 387.130 819.730 ;
        RECT 387.970 815.720 391.270 819.730 ;
        RECT 392.110 815.720 395.870 819.730 ;
        RECT 396.710 815.720 400.010 819.730 ;
        RECT 400.850 815.720 404.610 819.730 ;
        RECT 405.450 815.720 408.750 819.730 ;
        RECT 409.590 815.720 413.350 819.730 ;
        RECT 414.190 815.720 417.490 819.730 ;
        RECT 418.330 815.720 421.630 819.730 ;
        RECT 422.470 815.720 426.230 819.730 ;
        RECT 427.070 815.720 430.370 819.730 ;
        RECT 431.210 815.720 434.970 819.730 ;
        RECT 435.810 815.720 439.110 819.730 ;
        RECT 439.950 815.720 443.710 819.730 ;
        RECT 444.550 815.720 447.850 819.730 ;
        RECT 448.690 815.720 451.990 819.730 ;
        RECT 452.830 815.720 456.590 819.730 ;
        RECT 457.430 815.720 460.730 819.730 ;
        RECT 461.570 815.720 465.330 819.730 ;
        RECT 466.170 815.720 469.470 819.730 ;
        RECT 470.310 815.720 474.070 819.730 ;
        RECT 474.910 815.720 478.210 819.730 ;
        RECT 479.050 815.720 482.350 819.730 ;
        RECT 483.190 815.720 486.950 819.730 ;
        RECT 487.790 815.720 491.090 819.730 ;
        RECT 491.930 815.720 495.690 819.730 ;
        RECT 496.530 815.720 499.830 819.730 ;
        RECT 500.670 815.720 503.970 819.730 ;
        RECT 504.810 815.720 508.570 819.730 ;
        RECT 509.410 815.720 512.710 819.730 ;
        RECT 513.550 815.720 517.310 819.730 ;
        RECT 518.150 815.720 521.450 819.730 ;
        RECT 522.290 815.720 526.050 819.730 ;
        RECT 526.890 815.720 530.190 819.730 ;
        RECT 531.030 815.720 534.330 819.730 ;
        RECT 535.170 815.720 538.930 819.730 ;
        RECT 539.770 815.720 543.070 819.730 ;
        RECT 543.910 815.720 547.670 819.730 ;
        RECT 548.510 815.720 551.810 819.730 ;
        RECT 552.650 815.720 556.410 819.730 ;
        RECT 557.250 815.720 560.550 819.730 ;
        RECT 561.390 815.720 564.690 819.730 ;
        RECT 565.530 815.720 569.290 819.730 ;
        RECT 570.130 815.720 573.430 819.730 ;
        RECT 574.270 815.720 578.030 819.730 ;
        RECT 578.870 815.720 582.170 819.730 ;
        RECT 583.010 815.720 586.310 819.730 ;
        RECT 587.150 815.720 590.910 819.730 ;
        RECT 591.750 815.720 595.050 819.730 ;
        RECT 595.890 815.720 599.650 819.730 ;
        RECT 600.490 815.720 603.790 819.730 ;
        RECT 604.630 815.720 608.390 819.730 ;
        RECT 609.230 815.720 612.530 819.730 ;
        RECT 613.370 815.720 616.670 819.730 ;
        RECT 617.510 815.720 621.270 819.730 ;
        RECT 622.110 815.720 625.410 819.730 ;
        RECT 626.250 815.720 630.010 819.730 ;
        RECT 630.850 815.720 634.150 819.730 ;
        RECT 634.990 815.720 638.750 819.730 ;
        RECT 639.590 815.720 642.890 819.730 ;
        RECT 643.730 815.720 647.030 819.730 ;
        RECT 647.870 815.720 651.630 819.730 ;
        RECT 652.470 815.720 655.770 819.730 ;
        RECT 656.610 815.720 660.370 819.730 ;
        RECT 661.210 815.720 664.510 819.730 ;
        RECT 665.350 815.720 669.110 819.730 ;
        RECT 669.950 815.720 673.250 819.730 ;
        RECT 674.090 815.720 677.390 819.730 ;
        RECT 678.230 815.720 681.990 819.730 ;
        RECT 682.830 815.720 686.130 819.730 ;
        RECT 686.970 815.720 690.730 819.730 ;
        RECT 691.570 815.720 694.870 819.730 ;
        RECT 695.710 815.720 699.010 819.730 ;
        RECT 699.850 815.720 703.610 819.730 ;
        RECT 704.450 815.720 707.750 819.730 ;
        RECT 708.590 815.720 712.350 819.730 ;
        RECT 713.190 815.720 716.490 819.730 ;
        RECT 717.330 815.720 721.090 819.730 ;
        RECT 721.930 815.720 725.230 819.730 ;
        RECT 726.070 815.720 729.370 819.730 ;
        RECT 730.210 815.720 733.970 819.730 ;
        RECT 734.810 815.720 738.110 819.730 ;
        RECT 738.950 815.720 742.710 819.730 ;
        RECT 743.550 815.720 746.850 819.730 ;
        RECT 747.690 815.720 751.450 819.730 ;
        RECT 752.290 815.720 755.590 819.730 ;
        RECT 756.430 815.720 759.730 819.730 ;
        RECT 760.570 815.720 764.330 819.730 ;
        RECT 765.170 815.720 768.470 819.730 ;
        RECT 769.310 815.720 773.070 819.730 ;
        RECT 773.910 815.720 777.210 819.730 ;
        RECT 778.050 815.720 781.350 819.730 ;
        RECT 782.190 815.720 785.950 819.730 ;
        RECT 786.790 815.720 790.090 819.730 ;
        RECT 790.930 815.720 794.690 819.730 ;
        RECT 795.530 815.720 798.830 819.730 ;
        RECT 799.670 815.720 803.430 819.730 ;
        RECT 804.270 815.720 807.570 819.730 ;
        RECT 808.410 815.720 811.710 819.730 ;
        RECT 812.550 815.720 816.310 819.730 ;
        RECT 817.150 815.720 820.450 819.730 ;
        RECT 821.290 815.720 825.050 819.730 ;
        RECT 825.890 815.720 829.190 819.730 ;
        RECT 830.030 815.720 833.790 819.730 ;
        RECT 834.630 815.720 837.930 819.730 ;
        RECT 838.770 815.720 842.070 819.730 ;
        RECT 842.910 815.720 846.670 819.730 ;
        RECT 847.510 815.720 850.810 819.730 ;
        RECT 851.650 815.720 855.410 819.730 ;
        RECT 856.250 815.720 859.550 819.730 ;
        RECT 860.390 815.720 864.150 819.730 ;
        RECT 864.990 815.720 868.290 819.730 ;
        RECT 869.130 815.720 872.430 819.730 ;
        RECT 873.270 815.720 877.030 819.730 ;
        RECT 877.870 815.720 881.170 819.730 ;
        RECT 882.010 815.720 885.770 819.730 ;
        RECT 886.610 815.720 889.910 819.730 ;
        RECT 890.750 815.720 894.050 819.730 ;
        RECT 894.890 815.720 898.650 819.730 ;
        RECT 899.490 815.720 902.790 819.730 ;
        RECT 903.630 815.720 907.390 819.730 ;
        RECT 908.230 815.720 911.530 819.730 ;
        RECT 912.370 815.720 916.130 819.730 ;
        RECT 916.970 815.720 920.270 819.730 ;
        RECT 921.110 815.720 924.410 819.730 ;
        RECT 925.250 815.720 929.010 819.730 ;
        RECT 929.850 815.720 933.150 819.730 ;
        RECT 933.990 815.720 937.750 819.730 ;
        RECT 938.590 815.720 941.890 819.730 ;
        RECT 942.730 815.720 946.490 819.730 ;
        RECT 947.330 815.720 950.630 819.730 ;
        RECT 951.470 815.720 954.770 819.730 ;
        RECT 955.610 815.720 959.370 819.730 ;
        RECT 960.210 815.720 963.510 819.730 ;
        RECT 964.350 815.720 968.110 819.730 ;
        RECT 968.950 815.720 972.250 819.730 ;
        RECT 973.090 815.720 976.390 819.730 ;
        RECT 977.230 815.720 980.990 819.730 ;
        RECT 981.830 815.720 985.130 819.730 ;
        RECT 985.970 815.720 989.730 819.730 ;
        RECT 990.570 815.720 993.870 819.730 ;
        RECT 994.710 815.720 998.470 819.730 ;
        RECT 999.310 815.720 1002.610 819.730 ;
        RECT 1003.450 815.720 1006.750 819.730 ;
        RECT 1007.590 815.720 1011.350 819.730 ;
        RECT 1012.190 815.720 1015.490 819.730 ;
        RECT 1016.330 815.720 1020.090 819.730 ;
        RECT 1020.930 815.720 1024.230 819.730 ;
        RECT 1025.070 815.720 1028.830 819.730 ;
        RECT 1029.670 815.720 1032.970 819.730 ;
        RECT 1033.810 815.720 1037.110 819.730 ;
        RECT 1037.950 815.720 1041.710 819.730 ;
        RECT 1042.550 815.720 1045.850 819.730 ;
        RECT 1046.690 815.720 1050.450 819.730 ;
        RECT 1051.290 815.720 1054.590 819.730 ;
        RECT 1055.430 815.720 1059.190 819.730 ;
        RECT 1060.030 815.720 1063.330 819.730 ;
        RECT 1064.170 815.720 1067.470 819.730 ;
        RECT 1068.310 815.720 1072.070 819.730 ;
        RECT 1072.910 815.720 1076.210 819.730 ;
        RECT 1077.050 815.720 1080.810 819.730 ;
        RECT 1081.650 815.720 1084.950 819.730 ;
        RECT 1085.790 815.720 1089.090 819.730 ;
        RECT 1089.930 815.720 1093.690 819.730 ;
        RECT 1094.530 815.720 1097.830 819.730 ;
        RECT 1098.670 815.720 1102.430 819.730 ;
        RECT 1103.270 815.720 1106.570 819.730 ;
        RECT 1107.410 815.720 1111.170 819.730 ;
        RECT 1112.010 815.720 1115.310 819.730 ;
        RECT 1116.150 815.720 1119.450 819.730 ;
        RECT 1120.290 815.720 1124.050 819.730 ;
        RECT 1124.890 815.720 1128.190 819.730 ;
        RECT 1129.030 815.720 1132.790 819.730 ;
        RECT 1133.630 815.720 1136.930 819.730 ;
        RECT 1137.770 815.720 1141.530 819.730 ;
        RECT 1142.370 815.720 1145.670 819.730 ;
        RECT 1146.510 815.720 1149.810 819.730 ;
        RECT 1150.650 815.720 1154.410 819.730 ;
        RECT 1155.250 815.720 1158.550 819.730 ;
        RECT 1159.390 815.720 1163.150 819.730 ;
        RECT 1163.990 815.720 1167.290 819.730 ;
        RECT 1168.130 815.720 1171.430 819.730 ;
        RECT 1172.270 815.720 1176.030 819.730 ;
        RECT 1176.870 815.720 1180.170 819.730 ;
        RECT 1181.010 815.720 1184.770 819.730 ;
        RECT 1185.610 815.720 1188.910 819.730 ;
        RECT 1189.750 815.720 1193.510 819.730 ;
        RECT 1194.350 815.720 1197.650 819.730 ;
        RECT 1198.490 815.720 1201.790 819.730 ;
        RECT 1202.630 815.720 1206.390 819.730 ;
        RECT 1207.230 815.720 1210.530 819.730 ;
        RECT 1211.370 815.720 1215.130 819.730 ;
        RECT 1215.970 815.720 1219.270 819.730 ;
        RECT 1220.110 815.720 1223.870 819.730 ;
        RECT 1224.710 815.720 1228.010 819.730 ;
        RECT 1228.850 815.720 1232.150 819.730 ;
        RECT 1232.990 815.720 1236.750 819.730 ;
        RECT 1237.590 815.720 1240.890 819.730 ;
        RECT 1241.730 815.720 1245.490 819.730 ;
        RECT 1246.330 815.720 1249.630 819.730 ;
        RECT 1250.470 815.720 1254.230 819.730 ;
        RECT 1255.070 815.720 1258.370 819.730 ;
        RECT 1259.210 815.720 1262.510 819.730 ;
        RECT 1263.350 815.720 1267.110 819.730 ;
        RECT 1267.950 815.720 1271.250 819.730 ;
        RECT 1272.090 815.720 1275.850 819.730 ;
        RECT 1276.690 815.720 1279.990 819.730 ;
        RECT 1280.830 815.720 1284.130 819.730 ;
        RECT 1284.970 815.720 1288.730 819.730 ;
        RECT 1289.570 815.720 1292.870 819.730 ;
        RECT 1293.710 815.720 1297.470 819.730 ;
        RECT 1298.310 815.720 1301.610 819.730 ;
        RECT 1302.450 815.720 1306.210 819.730 ;
        RECT 1307.050 815.720 1310.350 819.730 ;
        RECT 1311.190 815.720 1314.490 819.730 ;
        RECT 1315.330 815.720 1319.090 819.730 ;
        RECT 1319.930 815.720 1323.230 819.730 ;
        RECT 1324.070 815.720 1327.830 819.730 ;
        RECT 1328.670 815.720 1331.970 819.730 ;
        RECT 1332.810 815.720 1336.570 819.730 ;
        RECT 1337.410 815.720 1340.710 819.730 ;
        RECT 1341.550 815.720 1344.850 819.730 ;
        RECT 1345.690 815.720 1349.450 819.730 ;
        RECT 1350.290 815.720 1353.590 819.730 ;
        RECT 1354.430 815.720 1358.190 819.730 ;
        RECT 1359.030 815.720 1362.330 819.730 ;
        RECT 1363.170 815.720 1366.470 819.730 ;
        RECT 1367.310 815.720 1371.070 819.730 ;
        RECT 1371.910 815.720 1375.210 819.730 ;
        RECT 1376.050 815.720 1379.810 819.730 ;
        RECT 1380.650 815.720 1383.950 819.730 ;
        RECT 1384.790 815.720 1388.550 819.730 ;
        RECT 1389.390 815.720 1392.690 819.730 ;
        RECT 1393.530 815.720 1396.830 819.730 ;
        RECT 1397.670 815.720 1401.430 819.730 ;
        RECT 1402.270 815.720 1405.570 819.730 ;
        RECT 1406.410 815.720 1410.170 819.730 ;
        RECT 1411.010 815.720 1414.310 819.730 ;
        RECT 1415.150 815.720 1418.910 819.730 ;
        RECT 1419.750 815.720 1423.050 819.730 ;
        RECT 1423.890 815.720 1427.190 819.730 ;
        RECT 1428.030 815.720 1431.790 819.730 ;
        RECT 1432.630 815.720 1435.930 819.730 ;
        RECT 1436.770 815.720 1440.530 819.730 ;
        RECT 1441.370 815.720 1444.670 819.730 ;
        RECT 1445.510 815.720 1448.810 819.730 ;
        RECT 1449.650 815.720 1453.410 819.730 ;
        RECT 1454.250 815.720 1457.550 819.730 ;
        RECT 1458.390 815.720 1462.150 819.730 ;
        RECT 1462.990 815.720 1466.290 819.730 ;
        RECT 1467.130 815.720 1470.890 819.730 ;
        RECT 1471.730 815.720 1475.030 819.730 ;
        RECT 1475.870 815.720 1479.170 819.730 ;
        RECT 1480.010 815.720 1483.770 819.730 ;
        RECT 1484.610 815.720 1487.910 819.730 ;
        RECT 1488.750 815.720 1492.510 819.730 ;
        RECT 1493.350 815.720 1496.650 819.730 ;
        RECT 1497.490 815.720 1501.250 819.730 ;
        RECT 1502.090 815.720 1505.390 819.730 ;
        RECT 1506.230 815.720 1509.530 819.730 ;
        RECT 1510.370 815.720 1514.130 819.730 ;
        RECT 1514.970 815.720 1518.270 819.730 ;
        RECT 1519.110 815.720 1522.870 819.730 ;
        RECT 1523.710 815.720 1527.010 819.730 ;
        RECT 1527.850 815.720 1531.610 819.730 ;
        RECT 1532.450 815.720 1535.750 819.730 ;
        RECT 1536.590 815.720 1539.890 819.730 ;
        RECT 1540.730 815.720 1544.490 819.730 ;
        RECT 1545.330 815.720 1548.630 819.730 ;
        RECT 1549.470 815.720 1553.230 819.730 ;
        RECT 1554.070 815.720 1557.370 819.730 ;
        RECT 1558.210 815.720 1561.510 819.730 ;
        RECT 1562.350 815.720 1566.110 819.730 ;
        RECT 1566.950 815.720 1570.250 819.730 ;
        RECT 1571.090 815.720 1574.850 819.730 ;
        RECT 1575.690 815.720 1578.990 819.730 ;
        RECT 1579.830 815.720 1583.590 819.730 ;
        RECT 1584.430 815.720 1587.730 819.730 ;
        RECT 1588.570 815.720 1591.870 819.730 ;
        RECT 1592.710 815.720 1596.470 819.730 ;
        RECT 1597.310 815.720 1600.610 819.730 ;
        RECT 1601.450 815.720 1605.210 819.730 ;
        RECT 1606.050 815.720 1609.350 819.730 ;
        RECT 1610.190 815.720 1613.950 819.730 ;
        RECT 1614.790 815.720 1618.090 819.730 ;
        RECT 1618.930 815.720 1622.230 819.730 ;
        RECT 1623.070 815.720 1626.830 819.730 ;
        RECT 1627.670 815.720 1630.970 819.730 ;
        RECT 1631.810 815.720 1635.570 819.730 ;
        RECT 1636.410 815.720 1639.710 819.730 ;
        RECT 1640.550 815.720 1643.850 819.730 ;
        RECT 1644.690 815.720 1648.450 819.730 ;
        RECT 1649.290 815.720 1652.590 819.730 ;
        RECT 1653.430 815.720 1657.190 819.730 ;
        RECT 1658.030 815.720 1661.330 819.730 ;
        RECT 1662.170 815.720 1665.930 819.730 ;
        RECT 1666.770 815.720 1670.070 819.730 ;
        RECT 1670.910 815.720 1674.210 819.730 ;
        RECT 1675.050 815.720 1678.810 819.730 ;
        RECT 1679.650 815.720 1682.950 819.730 ;
        RECT 1683.790 815.720 1687.550 819.730 ;
        RECT 1688.390 815.720 1691.690 819.730 ;
        RECT 1692.530 815.720 1696.290 819.730 ;
        RECT 1697.130 815.720 1700.430 819.730 ;
        RECT 1701.270 815.720 1704.570 819.730 ;
        RECT 1705.410 815.720 1709.170 819.730 ;
        RECT 1710.010 815.720 1713.310 819.730 ;
        RECT 1714.150 815.720 1717.910 819.730 ;
        RECT 1718.750 815.720 1722.050 819.730 ;
        RECT 1722.890 815.720 1726.650 819.730 ;
        RECT 1727.490 815.720 1730.790 819.730 ;
        RECT 1731.630 815.720 1734.930 819.730 ;
        RECT 1735.770 815.720 1739.530 819.730 ;
        RECT 1740.370 815.720 1743.670 819.730 ;
        RECT 1744.510 815.720 1748.270 819.730 ;
        RECT 1749.110 815.720 1752.410 819.730 ;
        RECT 1753.250 815.720 1756.550 819.730 ;
        RECT 1757.390 815.720 1761.150 819.730 ;
        RECT 1761.990 815.720 1765.290 819.730 ;
        RECT 1766.130 815.720 1769.890 819.730 ;
        RECT 1770.730 815.720 1774.030 819.730 ;
        RECT 1774.870 815.720 1778.630 819.730 ;
        RECT 1779.470 815.720 1782.770 819.730 ;
        RECT 1783.610 815.720 1786.910 819.730 ;
        RECT 1787.750 815.720 1791.510 819.730 ;
        RECT 1792.350 815.720 1795.650 819.730 ;
        RECT 1796.490 815.720 1800.250 819.730 ;
        RECT 1801.090 815.720 1804.390 819.730 ;
        RECT 1805.230 815.720 1808.990 819.730 ;
        RECT 1809.830 815.720 1813.130 819.730 ;
        RECT 1813.970 815.720 1817.270 819.730 ;
        RECT 1818.110 815.720 1821.870 819.730 ;
        RECT 1822.710 815.720 1826.010 819.730 ;
        RECT 1826.850 815.720 1830.610 819.730 ;
        RECT 1831.450 815.720 1834.750 819.730 ;
        RECT 1835.590 815.720 1838.890 819.730 ;
        RECT 1839.730 815.720 1843.490 819.730 ;
        RECT 1844.330 815.720 1847.630 819.730 ;
        RECT 1848.470 815.720 1852.230 819.730 ;
        RECT 1853.070 815.720 1856.370 819.730 ;
        RECT 1857.210 815.720 1860.970 819.730 ;
        RECT 1861.810 815.720 1865.110 819.730 ;
        RECT 1865.950 815.720 1869.250 819.730 ;
        RECT 1870.090 815.720 1873.850 819.730 ;
        RECT 1874.690 815.720 1877.990 819.730 ;
        RECT 1878.830 815.720 1882.590 819.730 ;
        RECT 1883.430 815.720 1886.730 819.730 ;
        RECT 1887.570 815.720 1891.330 819.730 ;
        RECT 1892.170 815.720 1895.470 819.730 ;
        RECT 1896.310 815.720 1899.610 819.730 ;
        RECT 1900.450 815.720 1904.210 819.730 ;
        RECT 1905.050 815.720 1908.350 819.730 ;
        RECT 1909.190 815.720 1912.950 819.730 ;
        RECT 1913.790 815.720 1917.090 819.730 ;
        RECT 1917.930 815.720 1921.690 819.730 ;
        RECT 1922.530 815.720 1925.830 819.730 ;
        RECT 1926.670 815.720 1929.970 819.730 ;
        RECT 1930.810 815.720 1934.570 819.730 ;
        RECT 1935.410 815.720 1938.710 819.730 ;
        RECT 1939.550 815.720 1943.310 819.730 ;
        RECT 1944.150 815.720 1947.450 819.730 ;
        RECT 1948.290 815.720 1951.590 819.730 ;
        RECT 1952.430 815.720 1956.190 819.730 ;
        RECT 1957.030 815.720 1960.330 819.730 ;
        RECT 1961.170 815.720 1964.930 819.730 ;
        RECT 1965.770 815.720 1969.070 819.730 ;
        RECT 1969.910 815.720 1973.670 819.730 ;
        RECT 1974.510 815.720 1977.810 819.730 ;
        RECT 1978.650 815.720 1981.950 819.730 ;
        RECT 1982.790 815.720 1986.550 819.730 ;
        RECT 1987.390 815.720 1990.690 819.730 ;
        RECT 1991.530 815.720 1995.290 819.730 ;
        RECT 1996.130 815.720 1999.430 819.730 ;
        RECT 2000.270 815.720 2004.030 819.730 ;
        RECT 2004.870 815.720 2008.170 819.730 ;
        RECT 2009.010 815.720 2012.310 819.730 ;
        RECT 2013.150 815.720 2016.910 819.730 ;
        RECT 2017.750 815.720 2021.050 819.730 ;
        RECT 2021.890 815.720 2025.650 819.730 ;
        RECT 2026.490 815.720 2029.790 819.730 ;
        RECT 2030.630 815.720 2033.930 819.730 ;
        RECT 2034.770 815.720 2038.530 819.730 ;
        RECT 2039.370 815.720 2042.670 819.730 ;
        RECT 2043.510 815.720 2047.270 819.730 ;
        RECT 2048.110 815.720 2051.410 819.730 ;
        RECT 2052.250 815.720 2056.010 819.730 ;
        RECT 2056.850 815.720 2060.150 819.730 ;
        RECT 2060.990 815.720 2064.290 819.730 ;
        RECT 2065.130 815.720 2068.890 819.730 ;
        RECT 2069.730 815.720 2073.030 819.730 ;
        RECT 2073.870 815.720 2077.630 819.730 ;
        RECT 2078.470 815.720 2081.770 819.730 ;
        RECT 2082.610 815.720 2086.370 819.730 ;
        RECT 2087.210 815.720 2090.510 819.730 ;
        RECT 2091.350 815.720 2094.650 819.730 ;
        RECT 2095.490 815.720 2099.250 819.730 ;
        RECT 2100.090 815.720 2103.390 819.730 ;
        RECT 2104.230 815.720 2107.990 819.730 ;
        RECT 2108.830 815.720 2112.130 819.730 ;
        RECT 2112.970 815.720 2116.730 819.730 ;
        RECT 2117.570 815.720 2120.870 819.730 ;
        RECT 2121.710 815.720 2125.010 819.730 ;
        RECT 2125.850 815.720 2129.610 819.730 ;
        RECT 2130.450 815.720 2133.750 819.730 ;
        RECT 2134.590 815.720 2138.350 819.730 ;
        RECT 2139.190 815.720 2142.490 819.730 ;
        RECT 2143.330 815.720 2146.630 819.730 ;
        RECT 2147.470 815.720 2151.230 819.730 ;
        RECT 2152.070 815.720 2155.370 819.730 ;
        RECT 2156.210 815.720 2159.970 819.730 ;
        RECT 2160.810 815.720 2164.110 819.730 ;
        RECT 2164.950 815.720 2168.710 819.730 ;
        RECT 2169.550 815.720 2172.850 819.730 ;
        RECT 2173.690 815.720 2176.990 819.730 ;
        RECT 2177.830 815.720 2181.590 819.730 ;
        RECT 2182.430 815.720 2185.730 819.730 ;
        RECT 2186.570 815.720 2190.330 819.730 ;
        RECT 2191.170 815.720 2194.470 819.730 ;
        RECT 2195.310 815.720 2199.070 819.730 ;
        RECT 2199.910 815.720 2203.210 819.730 ;
        RECT 2204.050 815.720 2207.350 819.730 ;
        RECT 2208.190 815.720 2211.950 819.730 ;
        RECT 2212.790 815.720 2216.090 819.730 ;
        RECT 2216.930 815.720 2220.690 819.730 ;
        RECT 2221.530 815.720 2224.830 819.730 ;
        RECT 2225.670 815.720 2228.970 819.730 ;
        RECT 2229.810 815.720 2233.570 819.730 ;
        RECT 2234.410 815.720 2237.710 819.730 ;
        RECT 2238.550 815.720 2242.310 819.730 ;
        RECT 2243.150 815.720 2246.450 819.730 ;
        RECT 2247.290 815.720 2251.050 819.730 ;
        RECT 2251.890 815.720 2255.190 819.730 ;
        RECT 2256.030 815.720 2259.330 819.730 ;
        RECT 2260.170 815.720 2263.930 819.730 ;
        RECT 2264.770 815.720 2268.070 819.730 ;
        RECT 2268.910 815.720 2272.670 819.730 ;
        RECT 2273.510 815.720 2276.810 819.730 ;
        RECT 2277.650 815.720 2281.410 819.730 ;
        RECT 2282.250 815.720 2285.550 819.730 ;
        RECT 2286.390 815.720 2289.690 819.730 ;
        RECT 2290.530 815.720 2294.290 819.730 ;
        RECT 2295.130 815.720 2298.430 819.730 ;
        RECT 2299.270 815.720 2303.030 819.730 ;
        RECT 2303.870 815.720 2307.170 819.730 ;
        RECT 2308.010 815.720 2311.770 819.730 ;
        RECT 2312.610 815.720 2315.910 819.730 ;
        RECT 2316.750 815.720 2320.050 819.730 ;
        RECT 2320.890 815.720 2324.650 819.730 ;
        RECT 2325.490 815.720 2328.790 819.730 ;
        RECT 2329.630 815.720 2333.390 819.730 ;
        RECT 2334.230 815.720 2337.530 819.730 ;
        RECT 2338.370 815.720 2341.670 819.730 ;
        RECT 2342.510 815.720 2346.270 819.730 ;
        RECT 2347.110 815.720 2350.410 819.730 ;
        RECT 2351.250 815.720 2355.010 819.730 ;
        RECT 2355.850 815.720 2359.150 819.730 ;
        RECT 2359.990 815.720 2363.750 819.730 ;
        RECT 2364.590 815.720 2367.890 819.730 ;
        RECT 2368.730 815.720 2372.030 819.730 ;
        RECT 2372.870 815.720 2376.630 819.730 ;
        RECT 2377.470 815.720 2380.770 819.730 ;
        RECT 2381.610 815.720 2385.370 819.730 ;
        RECT 2386.210 815.720 2389.510 819.730 ;
        RECT 2390.350 815.720 2394.110 819.730 ;
        RECT 2394.950 815.720 2398.250 819.730 ;
        RECT 2399.090 815.720 2402.390 819.730 ;
        RECT 2403.230 815.720 2406.990 819.730 ;
        RECT 2407.830 815.720 2411.130 819.730 ;
        RECT 2411.970 815.720 2415.730 819.730 ;
        RECT 2416.570 815.720 2419.870 819.730 ;
        RECT 2420.710 815.720 2424.010 819.730 ;
        RECT 2424.850 815.720 2428.610 819.730 ;
        RECT 2429.450 815.720 2432.750 819.730 ;
        RECT 2433.590 815.720 2437.350 819.730 ;
        RECT 2438.190 815.720 2441.490 819.730 ;
        RECT 2442.330 815.720 2446.090 819.730 ;
        RECT 2446.930 815.720 2450.230 819.730 ;
        RECT 2451.070 815.720 2454.370 819.730 ;
        RECT 2455.210 815.720 2458.970 819.730 ;
        RECT 2459.810 815.720 2463.110 819.730 ;
        RECT 2463.950 815.720 2467.710 819.730 ;
        RECT 2468.550 815.720 2471.850 819.730 ;
        RECT 2472.690 815.720 2476.450 819.730 ;
        RECT 2477.290 815.720 2480.590 819.730 ;
        RECT 2481.430 815.720 2484.730 819.730 ;
        RECT 2485.570 815.720 2489.330 819.730 ;
        RECT 2490.170 815.720 2493.470 819.730 ;
        RECT 2494.310 815.720 2498.070 819.730 ;
        RECT 2498.910 815.720 2502.210 819.730 ;
        RECT 2503.050 815.720 2506.810 819.730 ;
        RECT 2507.650 815.720 2510.950 819.730 ;
        RECT 2511.790 815.720 2515.090 819.730 ;
        RECT 2515.930 815.720 2519.690 819.730 ;
        RECT 2520.530 815.720 2523.830 819.730 ;
        RECT 2524.670 815.720 2528.430 819.730 ;
        RECT 2529.270 815.720 2532.570 819.730 ;
        RECT 2533.410 815.720 2536.710 819.730 ;
        RECT 2537.550 815.720 2541.310 819.730 ;
        RECT 2542.150 815.720 2545.450 819.730 ;
        RECT 2546.290 815.720 2550.050 819.730 ;
        RECT 2550.890 815.720 2554.190 819.730 ;
        RECT 2555.030 815.720 2558.790 819.730 ;
        RECT 2559.630 815.720 2562.930 819.730 ;
        RECT 2563.770 815.720 2567.070 819.730 ;
        RECT 2567.910 815.720 2571.670 819.730 ;
        RECT 2572.510 815.720 2575.810 819.730 ;
        RECT 2576.650 815.720 2580.410 819.730 ;
        RECT 2581.250 815.720 2584.550 819.730 ;
        RECT 2585.390 815.720 2589.150 819.730 ;
        RECT 2589.990 815.720 2593.290 819.730 ;
        RECT 2594.130 815.720 2597.430 819.730 ;
        RECT 2598.270 815.720 2602.030 819.730 ;
        RECT 2602.870 815.720 2606.170 819.730 ;
        RECT 2607.010 815.720 2610.770 819.730 ;
        RECT 2611.610 815.720 2614.910 819.730 ;
        RECT 2615.750 815.720 2619.050 819.730 ;
        RECT 2619.890 815.720 2623.650 819.730 ;
        RECT 2624.490 815.720 2627.790 819.730 ;
        RECT 2628.630 815.720 2632.390 819.730 ;
        RECT 2633.230 815.720 2636.530 819.730 ;
        RECT 2637.370 815.720 2641.130 819.730 ;
        RECT 2641.970 815.720 2645.270 819.730 ;
        RECT 2646.110 815.720 2649.410 819.730 ;
        RECT 2650.250 815.720 2654.010 819.730 ;
        RECT 2654.850 815.720 2658.150 819.730 ;
        RECT 2658.990 815.720 2662.750 819.730 ;
        RECT 2663.590 815.720 2666.890 819.730 ;
        RECT 2667.730 815.720 2671.490 819.730 ;
        RECT 2672.330 815.720 2675.630 819.730 ;
        RECT 2676.470 815.720 2679.770 819.730 ;
        RECT 2680.610 815.720 2684.370 819.730 ;
        RECT 2685.210 815.720 2688.510 819.730 ;
        RECT 2689.350 815.720 2693.110 819.730 ;
        RECT 2693.950 815.720 2697.250 819.730 ;
        RECT 1.940 4.280 2697.800 815.720 ;
        RECT 1.940 3.555 168.170 4.280 ;
        RECT 169.010 3.555 505.350 4.280 ;
        RECT 506.190 3.555 842.990 4.280 ;
        RECT 843.830 3.555 1180.630 4.280 ;
        RECT 1181.470 3.555 1518.270 4.280 ;
        RECT 1519.110 3.555 1855.450 4.280 ;
        RECT 1856.290 3.555 2193.090 4.280 ;
        RECT 2193.930 3.555 2530.730 4.280 ;
        RECT 2531.570 3.555 2697.800 4.280 ;
      LAYER met3 ;
        RECT 29.965 814.960 2695.600 815.825 ;
        RECT 29.965 808.880 2696.000 814.960 ;
        RECT 29.965 807.480 2695.600 808.880 ;
        RECT 29.965 801.400 2696.000 807.480 ;
        RECT 29.965 800.000 2695.600 801.400 ;
        RECT 29.965 793.920 2696.000 800.000 ;
        RECT 29.965 792.520 2695.600 793.920 ;
        RECT 29.965 786.440 2696.000 792.520 ;
        RECT 29.965 785.040 2695.600 786.440 ;
        RECT 29.965 778.960 2696.000 785.040 ;
        RECT 29.965 777.560 2695.600 778.960 ;
        RECT 29.965 770.800 2696.000 777.560 ;
        RECT 29.965 769.400 2695.600 770.800 ;
        RECT 29.965 763.320 2696.000 769.400 ;
        RECT 29.965 761.920 2695.600 763.320 ;
        RECT 29.965 755.840 2696.000 761.920 ;
        RECT 29.965 754.440 2695.600 755.840 ;
        RECT 29.965 748.360 2696.000 754.440 ;
        RECT 29.965 746.960 2695.600 748.360 ;
        RECT 29.965 740.880 2696.000 746.960 ;
        RECT 29.965 739.480 2695.600 740.880 ;
        RECT 29.965 733.400 2696.000 739.480 ;
        RECT 29.965 732.000 2695.600 733.400 ;
        RECT 29.965 725.240 2696.000 732.000 ;
        RECT 29.965 723.840 2695.600 725.240 ;
        RECT 29.965 717.760 2696.000 723.840 ;
        RECT 29.965 716.360 2695.600 717.760 ;
        RECT 29.965 710.280 2696.000 716.360 ;
        RECT 29.965 708.880 2695.600 710.280 ;
        RECT 29.965 702.800 2696.000 708.880 ;
        RECT 29.965 701.400 2695.600 702.800 ;
        RECT 29.965 695.320 2696.000 701.400 ;
        RECT 29.965 693.920 2695.600 695.320 ;
        RECT 29.965 687.840 2696.000 693.920 ;
        RECT 29.965 686.440 2695.600 687.840 ;
        RECT 29.965 679.680 2696.000 686.440 ;
        RECT 29.965 678.280 2695.600 679.680 ;
        RECT 29.965 672.200 2696.000 678.280 ;
        RECT 29.965 670.800 2695.600 672.200 ;
        RECT 29.965 664.720 2696.000 670.800 ;
        RECT 29.965 663.320 2695.600 664.720 ;
        RECT 29.965 657.240 2696.000 663.320 ;
        RECT 29.965 655.840 2695.600 657.240 ;
        RECT 29.965 649.760 2696.000 655.840 ;
        RECT 29.965 648.360 2695.600 649.760 ;
        RECT 29.965 642.280 2696.000 648.360 ;
        RECT 29.965 640.880 2695.600 642.280 ;
        RECT 29.965 634.120 2696.000 640.880 ;
        RECT 29.965 632.720 2695.600 634.120 ;
        RECT 29.965 626.640 2696.000 632.720 ;
        RECT 29.965 625.240 2695.600 626.640 ;
        RECT 29.965 619.160 2696.000 625.240 ;
        RECT 29.965 617.760 2695.600 619.160 ;
        RECT 29.965 611.680 2696.000 617.760 ;
        RECT 29.965 610.280 2695.600 611.680 ;
        RECT 29.965 604.200 2696.000 610.280 ;
        RECT 29.965 602.800 2695.600 604.200 ;
        RECT 29.965 596.720 2696.000 602.800 ;
        RECT 29.965 595.320 2695.600 596.720 ;
        RECT 29.965 588.560 2696.000 595.320 ;
        RECT 29.965 587.160 2695.600 588.560 ;
        RECT 29.965 581.080 2696.000 587.160 ;
        RECT 29.965 579.680 2695.600 581.080 ;
        RECT 29.965 573.600 2696.000 579.680 ;
        RECT 29.965 572.200 2695.600 573.600 ;
        RECT 29.965 566.120 2696.000 572.200 ;
        RECT 29.965 564.720 2695.600 566.120 ;
        RECT 29.965 558.640 2696.000 564.720 ;
        RECT 29.965 557.240 2695.600 558.640 ;
        RECT 29.965 551.160 2696.000 557.240 ;
        RECT 29.965 549.760 2695.600 551.160 ;
        RECT 29.965 543.000 2696.000 549.760 ;
        RECT 29.965 541.600 2695.600 543.000 ;
        RECT 29.965 535.520 2696.000 541.600 ;
        RECT 29.965 534.120 2695.600 535.520 ;
        RECT 29.965 528.040 2696.000 534.120 ;
        RECT 29.965 526.640 2695.600 528.040 ;
        RECT 29.965 520.560 2696.000 526.640 ;
        RECT 29.965 519.160 2695.600 520.560 ;
        RECT 29.965 513.080 2696.000 519.160 ;
        RECT 29.965 511.680 2695.600 513.080 ;
        RECT 29.965 505.600 2696.000 511.680 ;
        RECT 29.965 504.200 2695.600 505.600 ;
        RECT 29.965 497.440 2696.000 504.200 ;
        RECT 29.965 496.040 2695.600 497.440 ;
        RECT 29.965 489.960 2696.000 496.040 ;
        RECT 29.965 488.560 2695.600 489.960 ;
        RECT 29.965 482.480 2696.000 488.560 ;
        RECT 29.965 481.080 2695.600 482.480 ;
        RECT 29.965 475.000 2696.000 481.080 ;
        RECT 29.965 473.600 2695.600 475.000 ;
        RECT 29.965 467.520 2696.000 473.600 ;
        RECT 29.965 466.120 2695.600 467.520 ;
        RECT 29.965 460.040 2696.000 466.120 ;
        RECT 29.965 458.640 2695.600 460.040 ;
        RECT 29.965 451.880 2696.000 458.640 ;
        RECT 29.965 450.480 2695.600 451.880 ;
        RECT 29.965 444.400 2696.000 450.480 ;
        RECT 29.965 443.000 2695.600 444.400 ;
        RECT 29.965 436.920 2696.000 443.000 ;
        RECT 29.965 435.520 2695.600 436.920 ;
        RECT 29.965 429.440 2696.000 435.520 ;
        RECT 29.965 428.040 2695.600 429.440 ;
        RECT 29.965 421.960 2696.000 428.040 ;
        RECT 29.965 420.560 2695.600 421.960 ;
        RECT 29.965 414.480 2696.000 420.560 ;
        RECT 29.965 413.080 2695.600 414.480 ;
        RECT 29.965 406.320 2696.000 413.080 ;
        RECT 29.965 404.920 2695.600 406.320 ;
        RECT 29.965 398.840 2696.000 404.920 ;
        RECT 29.965 397.440 2695.600 398.840 ;
        RECT 29.965 391.360 2696.000 397.440 ;
        RECT 29.965 389.960 2695.600 391.360 ;
        RECT 29.965 383.880 2696.000 389.960 ;
        RECT 29.965 382.480 2695.600 383.880 ;
        RECT 29.965 376.400 2696.000 382.480 ;
        RECT 29.965 375.000 2695.600 376.400 ;
        RECT 29.965 368.920 2696.000 375.000 ;
        RECT 29.965 367.520 2695.600 368.920 ;
        RECT 29.965 360.760 2696.000 367.520 ;
        RECT 29.965 359.360 2695.600 360.760 ;
        RECT 29.965 353.280 2696.000 359.360 ;
        RECT 29.965 351.880 2695.600 353.280 ;
        RECT 29.965 345.800 2696.000 351.880 ;
        RECT 29.965 344.400 2695.600 345.800 ;
        RECT 29.965 338.320 2696.000 344.400 ;
        RECT 29.965 336.920 2695.600 338.320 ;
        RECT 29.965 330.840 2696.000 336.920 ;
        RECT 29.965 329.440 2695.600 330.840 ;
        RECT 29.965 323.360 2696.000 329.440 ;
        RECT 29.965 321.960 2695.600 323.360 ;
        RECT 29.965 315.200 2696.000 321.960 ;
        RECT 29.965 313.800 2695.600 315.200 ;
        RECT 29.965 307.720 2696.000 313.800 ;
        RECT 29.965 306.320 2695.600 307.720 ;
        RECT 29.965 300.240 2696.000 306.320 ;
        RECT 29.965 298.840 2695.600 300.240 ;
        RECT 29.965 292.760 2696.000 298.840 ;
        RECT 29.965 291.360 2695.600 292.760 ;
        RECT 29.965 285.280 2696.000 291.360 ;
        RECT 29.965 283.880 2695.600 285.280 ;
        RECT 29.965 277.800 2696.000 283.880 ;
        RECT 29.965 276.400 2695.600 277.800 ;
        RECT 29.965 269.640 2696.000 276.400 ;
        RECT 29.965 268.240 2695.600 269.640 ;
        RECT 29.965 262.160 2696.000 268.240 ;
        RECT 29.965 260.760 2695.600 262.160 ;
        RECT 29.965 254.680 2696.000 260.760 ;
        RECT 29.965 253.280 2695.600 254.680 ;
        RECT 29.965 247.200 2696.000 253.280 ;
        RECT 29.965 245.800 2695.600 247.200 ;
        RECT 29.965 239.720 2696.000 245.800 ;
        RECT 29.965 238.320 2695.600 239.720 ;
        RECT 29.965 232.240 2696.000 238.320 ;
        RECT 29.965 230.840 2695.600 232.240 ;
        RECT 29.965 224.080 2696.000 230.840 ;
        RECT 29.965 222.680 2695.600 224.080 ;
        RECT 29.965 216.600 2696.000 222.680 ;
        RECT 29.965 215.200 2695.600 216.600 ;
        RECT 29.965 209.120 2696.000 215.200 ;
        RECT 29.965 207.720 2695.600 209.120 ;
        RECT 29.965 201.640 2696.000 207.720 ;
        RECT 29.965 200.240 2695.600 201.640 ;
        RECT 29.965 194.160 2696.000 200.240 ;
        RECT 29.965 192.760 2695.600 194.160 ;
        RECT 29.965 186.680 2696.000 192.760 ;
        RECT 29.965 185.280 2695.600 186.680 ;
        RECT 29.965 178.520 2696.000 185.280 ;
        RECT 29.965 177.120 2695.600 178.520 ;
        RECT 29.965 171.040 2696.000 177.120 ;
        RECT 29.965 169.640 2695.600 171.040 ;
        RECT 29.965 163.560 2696.000 169.640 ;
        RECT 29.965 162.160 2695.600 163.560 ;
        RECT 29.965 156.080 2696.000 162.160 ;
        RECT 29.965 154.680 2695.600 156.080 ;
        RECT 29.965 148.600 2696.000 154.680 ;
        RECT 29.965 147.200 2695.600 148.600 ;
        RECT 29.965 141.120 2696.000 147.200 ;
        RECT 29.965 139.720 2695.600 141.120 ;
        RECT 29.965 132.960 2696.000 139.720 ;
        RECT 29.965 131.560 2695.600 132.960 ;
        RECT 29.965 125.480 2696.000 131.560 ;
        RECT 29.965 124.080 2695.600 125.480 ;
        RECT 29.965 118.000 2696.000 124.080 ;
        RECT 29.965 116.600 2695.600 118.000 ;
        RECT 29.965 110.520 2696.000 116.600 ;
        RECT 29.965 109.120 2695.600 110.520 ;
        RECT 29.965 103.040 2696.000 109.120 ;
        RECT 29.965 101.640 2695.600 103.040 ;
        RECT 29.965 95.560 2696.000 101.640 ;
        RECT 29.965 94.160 2695.600 95.560 ;
        RECT 29.965 87.400 2696.000 94.160 ;
        RECT 29.965 86.000 2695.600 87.400 ;
        RECT 29.965 79.920 2696.000 86.000 ;
        RECT 29.965 78.520 2695.600 79.920 ;
        RECT 29.965 72.440 2696.000 78.520 ;
        RECT 29.965 71.040 2695.600 72.440 ;
        RECT 29.965 64.960 2696.000 71.040 ;
        RECT 29.965 63.560 2695.600 64.960 ;
        RECT 29.965 57.480 2696.000 63.560 ;
        RECT 29.965 56.080 2695.600 57.480 ;
        RECT 29.965 50.000 2696.000 56.080 ;
        RECT 29.965 48.600 2695.600 50.000 ;
        RECT 29.965 41.840 2696.000 48.600 ;
        RECT 29.965 40.440 2695.600 41.840 ;
        RECT 29.965 34.360 2696.000 40.440 ;
        RECT 29.965 32.960 2695.600 34.360 ;
        RECT 29.965 26.880 2696.000 32.960 ;
        RECT 29.965 25.480 2695.600 26.880 ;
        RECT 29.965 19.400 2696.000 25.480 ;
        RECT 29.965 18.000 2695.600 19.400 ;
        RECT 29.965 11.920 2696.000 18.000 ;
        RECT 29.965 10.520 2695.600 11.920 ;
        RECT 29.965 4.440 2696.000 10.520 ;
        RECT 29.965 3.575 2695.600 4.440 ;
      LAYER met4 ;
        RECT 20.020 20.780 2640.090 794.490 ;
      LAYER met5 ;
        RECT 20.020 744.930 2644.100 794.700 ;
        RECT 20.020 740.130 578.400 744.930 ;
        RECT 641.600 740.130 2644.100 744.930 ;
        RECT 20.020 679.930 2644.100 740.130 ;
        RECT 20.020 675.130 578.400 679.930 ;
        RECT 641.600 675.130 2644.100 679.930 ;
        RECT 20.020 614.930 2644.100 675.130 ;
        RECT 20.020 610.130 578.400 614.930 ;
        RECT 641.600 610.130 2644.100 614.930 ;
        RECT 20.020 549.930 2644.100 610.130 ;
        RECT 20.020 545.130 578.400 549.930 ;
        RECT 641.600 545.130 2644.100 549.930 ;
        RECT 20.020 484.930 2644.100 545.130 ;
        RECT 20.020 480.130 578.400 484.930 ;
        RECT 641.600 480.130 2644.100 484.930 ;
        RECT 20.020 419.930 2644.100 480.130 ;
        RECT 20.020 415.130 578.400 419.930 ;
        RECT 641.600 415.130 2644.100 419.930 ;
        RECT 20.020 354.930 2644.100 415.130 ;
        RECT 20.020 350.130 578.400 354.930 ;
        RECT 641.600 350.130 2644.100 354.930 ;
        RECT 20.020 289.930 2644.100 350.130 ;
        RECT 20.020 285.130 578.400 289.930 ;
        RECT 641.600 285.130 2644.100 289.930 ;
        RECT 20.020 224.930 2644.100 285.130 ;
        RECT 20.020 220.130 578.400 224.930 ;
        RECT 641.600 220.130 2644.100 224.930 ;
        RECT 20.020 159.930 2644.100 220.130 ;
        RECT 20.020 155.130 578.400 159.930 ;
        RECT 641.600 155.130 2644.100 159.930 ;
        RECT 20.020 94.930 2644.100 155.130 ;
        RECT 20.020 90.130 578.400 94.930 ;
        RECT 641.600 90.130 2644.100 94.930 ;
        RECT 20.020 29.930 2644.100 90.130 ;
        RECT 20.020 25.130 578.400 29.930 ;
        RECT 641.600 25.130 2644.100 29.930 ;
        RECT 20.020 20.780 2644.100 25.130 ;
  END
END mgmt_core_wrapper
END LIBRARY

