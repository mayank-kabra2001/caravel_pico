magic
tech sky130A
magscale 1 2
timestamp 1637331822
<< metal1 >>
rect 43254 162596 43260 162648
rect 43312 162636 43318 162648
rect 151906 162636 151912 162648
rect 43312 162608 151912 162636
rect 43312 162596 43318 162608
rect 151906 162596 151912 162608
rect 151964 162596 151970 162648
rect 39850 162528 39856 162580
rect 39908 162568 39914 162580
rect 149422 162568 149428 162580
rect 39908 162540 149428 162568
rect 39908 162528 39914 162540
rect 149422 162528 149428 162540
rect 149480 162528 149486 162580
rect 102134 162460 102140 162512
rect 102192 162500 102198 162512
rect 196894 162500 196900 162512
rect 102192 162472 196900 162500
rect 102192 162460 102198 162472
rect 196894 162460 196900 162472
rect 196952 162460 196958 162512
rect 108850 162392 108856 162444
rect 108908 162432 108914 162444
rect 202046 162432 202052 162444
rect 108908 162404 202052 162432
rect 108908 162392 108914 162404
rect 202046 162392 202052 162404
rect 202104 162392 202110 162444
rect 95418 162324 95424 162376
rect 95476 162364 95482 162376
rect 190730 162364 190736 162376
rect 95476 162336 190736 162364
rect 95476 162324 95482 162336
rect 190730 162324 190736 162336
rect 190788 162324 190794 162376
rect 98730 162256 98736 162308
rect 98788 162296 98794 162308
rect 193398 162296 193404 162308
rect 98788 162268 193404 162296
rect 98788 162256 98794 162268
rect 193398 162256 193404 162268
rect 193456 162256 193462 162308
rect 92014 162188 92020 162240
rect 92072 162228 92078 162240
rect 189166 162228 189172 162240
rect 92072 162200 189172 162228
rect 92072 162188 92078 162200
rect 189166 162188 189172 162200
rect 189224 162188 189230 162240
rect 88702 162120 88708 162172
rect 88760 162160 88766 162172
rect 186314 162160 186320 162172
rect 88760 162132 186320 162160
rect 88760 162120 88766 162132
rect 186314 162120 186320 162132
rect 186372 162120 186378 162172
rect 81894 162052 81900 162104
rect 81952 162092 81958 162104
rect 181070 162092 181076 162104
rect 81952 162064 181076 162092
rect 81952 162052 81958 162064
rect 181070 162052 181076 162064
rect 181128 162052 181134 162104
rect 71866 161984 71872 162036
rect 71924 162024 71930 162036
rect 172698 162024 172704 162036
rect 71924 161996 172704 162024
rect 71924 161984 71930 161996
rect 172698 161984 172704 161996
rect 172756 161984 172762 162036
rect 78582 161916 78588 161968
rect 78640 161956 78646 161968
rect 178218 161956 178224 161968
rect 78640 161928 178224 161956
rect 78640 161916 78646 161928
rect 178218 161916 178224 161928
rect 178276 161916 178282 161968
rect 75178 161848 75184 161900
rect 75236 161888 75242 161900
rect 175550 161888 175556 161900
rect 75236 161860 175556 161888
rect 75236 161848 75242 161860
rect 175550 161848 175556 161860
rect 175608 161848 175614 161900
rect 65150 161780 65156 161832
rect 65208 161820 65214 161832
rect 168466 161820 168472 161832
rect 65208 161792 168472 161820
rect 65208 161780 65214 161792
rect 168466 161780 168472 161792
rect 168524 161780 168530 161832
rect 68462 161712 68468 161764
rect 68520 161752 68526 161764
rect 171318 161752 171324 161764
rect 68520 161724 171324 161752
rect 68520 161712 68526 161724
rect 171318 161712 171324 161724
rect 171376 161712 171382 161764
rect 61746 161644 61752 161696
rect 61804 161684 61810 161696
rect 165614 161684 165620 161696
rect 61804 161656 165620 161684
rect 61804 161644 61810 161656
rect 165614 161644 165620 161656
rect 165672 161644 165678 161696
rect 56686 161576 56692 161628
rect 56744 161616 56750 161628
rect 161474 161616 161480 161628
rect 56744 161588 161480 161616
rect 56744 161576 56750 161588
rect 161474 161576 161480 161588
rect 161532 161576 161538 161628
rect 115566 161508 115572 161560
rect 115624 161548 115630 161560
rect 207198 161548 207204 161560
rect 115624 161520 207204 161548
rect 115624 161508 115630 161520
rect 207198 161508 207204 161520
rect 207256 161508 207262 161560
rect 112254 161440 112260 161492
rect 112312 161480 112318 161492
rect 204254 161480 204260 161492
rect 112312 161452 204260 161480
rect 112312 161440 112318 161452
rect 204254 161440 204260 161452
rect 204312 161440 204318 161492
rect 114738 161372 114744 161424
rect 114796 161412 114802 161424
rect 206186 161412 206192 161424
rect 114796 161384 206192 161412
rect 114796 161372 114802 161384
rect 206186 161372 206192 161384
rect 206244 161372 206250 161424
rect 108022 161304 108028 161356
rect 108080 161344 108086 161356
rect 200298 161344 200304 161356
rect 108080 161316 200304 161344
rect 108080 161304 108086 161316
rect 200298 161304 200304 161316
rect 200356 161304 200362 161356
rect 101306 161236 101312 161288
rect 101364 161276 101370 161288
rect 196250 161276 196256 161288
rect 101364 161248 196256 161276
rect 101364 161236 101370 161248
rect 196250 161236 196256 161248
rect 196308 161236 196314 161288
rect 94590 161168 94596 161220
rect 94648 161208 94654 161220
rect 191098 161208 191104 161220
rect 94648 161180 191104 161208
rect 94648 161168 94654 161180
rect 191098 161168 191104 161180
rect 191156 161168 191162 161220
rect 205542 161168 205548 161220
rect 205600 161208 205606 161220
rect 275186 161208 275192 161220
rect 205600 161180 275192 161208
rect 205600 161168 205606 161180
rect 275186 161168 275192 161180
rect 275244 161168 275250 161220
rect 81066 161100 81072 161152
rect 81124 161140 81130 161152
rect 180886 161140 180892 161152
rect 81124 161112 180892 161140
rect 81124 161100 81130 161112
rect 180886 161100 180892 161112
rect 180944 161100 180950 161152
rect 198826 161100 198832 161152
rect 198884 161140 198890 161152
rect 270494 161140 270500 161152
rect 198884 161112 270500 161140
rect 198884 161100 198890 161112
rect 270494 161100 270500 161112
rect 270552 161100 270558 161152
rect 67634 161032 67640 161084
rect 67692 161072 67698 161084
rect 169754 161072 169760 161084
rect 67692 161044 169760 161072
rect 67692 161032 67698 161044
rect 169754 161032 169760 161044
rect 169812 161032 169818 161084
rect 183738 161032 183744 161084
rect 183796 161072 183802 161084
rect 258074 161072 258080 161084
rect 183796 161044 258080 161072
rect 183796 161032 183802 161044
rect 258074 161032 258080 161044
rect 258132 161032 258138 161084
rect 60918 160964 60924 161016
rect 60976 161004 60982 161016
rect 165430 161004 165436 161016
rect 60976 160976 165436 161004
rect 60976 160964 60982 160976
rect 165430 160964 165436 160976
rect 165488 160964 165494 161016
rect 175274 160964 175280 161016
rect 175332 161004 175338 161016
rect 252738 161004 252744 161016
rect 175332 160976 252744 161004
rect 175332 160964 175338 160976
rect 252738 160964 252744 160976
rect 252796 160964 252802 161016
rect 54202 160896 54208 160948
rect 54260 160936 54266 160948
rect 160370 160936 160376 160948
rect 54260 160908 160376 160936
rect 54260 160896 54266 160908
rect 160370 160896 160376 160908
rect 160428 160896 160434 160948
rect 166074 160896 166080 160948
rect 166132 160936 166138 160948
rect 245746 160936 245752 160948
rect 166132 160908 245752 160936
rect 166132 160896 166138 160908
rect 245746 160896 245752 160908
rect 245804 160896 245810 160948
rect 47486 160828 47492 160880
rect 47544 160868 47550 160880
rect 155034 160868 155040 160880
rect 47544 160840 155040 160868
rect 47544 160828 47550 160840
rect 155034 160828 155040 160840
rect 155092 160828 155098 160880
rect 161842 160828 161848 160880
rect 161900 160868 161906 160880
rect 242066 160868 242072 160880
rect 161900 160840 242072 160868
rect 161900 160828 161906 160840
rect 242066 160828 242072 160840
rect 242124 160828 242130 160880
rect 40678 160760 40684 160812
rect 40736 160800 40742 160812
rect 149146 160800 149152 160812
rect 40736 160772 149152 160800
rect 40736 160760 40742 160772
rect 149146 160760 149152 160772
rect 149204 160760 149210 160812
rect 155126 160760 155132 160812
rect 155184 160800 155190 160812
rect 237374 160800 237380 160812
rect 155184 160772 237380 160800
rect 155184 160760 155190 160772
rect 237374 160760 237380 160772
rect 237432 160760 237438 160812
rect 36538 160692 36544 160744
rect 36596 160732 36602 160744
rect 146846 160732 146852 160744
rect 36596 160704 146852 160732
rect 36596 160692 36602 160704
rect 146846 160692 146852 160704
rect 146904 160692 146910 160744
rect 148410 160692 148416 160744
rect 148468 160732 148474 160744
rect 232222 160732 232228 160744
rect 148468 160704 232228 160732
rect 148468 160692 148474 160704
rect 232222 160692 232228 160704
rect 232280 160692 232286 160744
rect 124858 160624 124864 160676
rect 124916 160664 124922 160676
rect 213914 160664 213920 160676
rect 124916 160636 213920 160664
rect 124916 160624 124922 160636
rect 213914 160624 213920 160636
rect 213972 160624 213978 160676
rect 141694 160556 141700 160608
rect 141752 160596 141758 160608
rect 227070 160596 227076 160608
rect 141752 160568 227076 160596
rect 141752 160556 141758 160568
rect 227070 160556 227076 160568
rect 227128 160556 227134 160608
rect 149238 160488 149244 160540
rect 149296 160528 149302 160540
rect 231946 160528 231952 160540
rect 149296 160500 231952 160528
rect 149296 160488 149302 160500
rect 231946 160488 231952 160500
rect 232004 160488 232010 160540
rect 49970 160012 49976 160064
rect 50028 160052 50034 160064
rect 109218 160052 109224 160064
rect 50028 160024 109224 160052
rect 50028 160012 50034 160024
rect 109218 160012 109224 160024
rect 109276 160012 109282 160064
rect 120626 160012 120632 160064
rect 120684 160052 120690 160064
rect 183278 160052 183284 160064
rect 120684 160024 183284 160052
rect 120684 160012 120690 160024
rect 183278 160012 183284 160024
rect 183336 160012 183342 160064
rect 187878 160012 187884 160064
rect 187936 160052 187942 160064
rect 210142 160052 210148 160064
rect 187936 160024 210148 160052
rect 187936 160012 187942 160024
rect 210142 160012 210148 160024
rect 210200 160012 210206 160064
rect 217318 160012 217324 160064
rect 217376 160052 217382 160064
rect 223482 160052 223488 160064
rect 217376 160024 223488 160052
rect 217376 160012 217382 160024
rect 223482 160012 223488 160024
rect 223540 160012 223546 160064
rect 228266 160012 228272 160064
rect 228324 160052 228330 160064
rect 239950 160052 239956 160064
rect 228324 160024 239956 160052
rect 228324 160012 228330 160024
rect 239950 160012 239956 160024
rect 240008 160012 240014 160064
rect 240870 160012 240876 160064
rect 240928 160052 240934 160064
rect 263870 160052 263876 160064
rect 240928 160024 263876 160052
rect 240928 160012 240934 160024
rect 263870 160012 263876 160024
rect 263928 160012 263934 160064
rect 265342 160012 265348 160064
rect 265400 160052 265406 160064
rect 311066 160052 311072 160064
rect 265400 160024 311072 160052
rect 265400 160012 265406 160024
rect 311066 160012 311072 160024
rect 311124 160012 311130 160064
rect 318334 160012 318340 160064
rect 318392 160052 318398 160064
rect 336642 160052 336648 160064
rect 318392 160024 336648 160052
rect 318392 160012 318398 160024
rect 336642 160012 336648 160024
rect 336700 160012 336706 160064
rect 342714 160012 342720 160064
rect 342772 160052 342778 160064
rect 372614 160052 372620 160064
rect 342772 160024 372620 160052
rect 342772 160012 342778 160024
rect 372614 160012 372620 160024
rect 372672 160012 372678 160064
rect 409138 160012 409144 160064
rect 409196 160052 409202 160064
rect 431218 160052 431224 160064
rect 409196 160024 431224 160052
rect 409196 160012 409202 160024
rect 431218 160012 431224 160024
rect 431276 160012 431282 160064
rect 457070 160012 457076 160064
rect 457128 160052 457134 160064
rect 464338 160052 464344 160064
rect 457128 160024 464344 160052
rect 457128 160012 457134 160024
rect 464338 160012 464344 160024
rect 464396 160012 464402 160064
rect 66806 159944 66812 159996
rect 66864 159984 66870 159996
rect 135622 159984 135628 159996
rect 66864 159956 135628 159984
rect 66864 159944 66870 159956
rect 135622 159944 135628 159956
rect 135680 159944 135686 159996
rect 164326 159944 164332 159996
rect 164384 159984 164390 159996
rect 221918 159984 221924 159996
rect 164384 159956 221924 159984
rect 164384 159944 164390 159956
rect 221918 159944 221924 159956
rect 221976 159944 221982 159996
rect 234154 159944 234160 159996
rect 234212 159984 234218 159996
rect 255498 159984 255504 159996
rect 234212 159956 255504 159984
rect 234212 159944 234218 159956
rect 255498 159944 255504 159956
rect 255556 159944 255562 159996
rect 258534 159944 258540 159996
rect 258592 159984 258598 159996
rect 304994 159984 305000 159996
rect 258592 159956 305000 159984
rect 258592 159944 258598 159956
rect 304994 159944 305000 159956
rect 305052 159944 305058 159996
rect 311526 159944 311532 159996
rect 311584 159984 311590 159996
rect 330202 159984 330208 159996
rect 311584 159956 330208 159984
rect 311584 159944 311590 159956
rect 330202 159944 330208 159956
rect 330260 159944 330266 159996
rect 332594 159944 332600 159996
rect 332652 159984 332658 159996
rect 368474 159984 368480 159996
rect 332652 159956 368480 159984
rect 332652 159944 332658 159956
rect 368474 159944 368480 159956
rect 368532 159944 368538 159996
rect 393130 159944 393136 159996
rect 393188 159984 393194 159996
rect 419074 159984 419080 159996
rect 393188 159956 419080 159984
rect 393188 159944 393194 159956
rect 419074 159944 419080 159956
rect 419132 159944 419138 159996
rect 425974 159944 425980 159996
rect 426032 159984 426038 159996
rect 426434 159984 426440 159996
rect 426032 159956 426440 159984
rect 426032 159944 426038 159956
rect 426434 159944 426440 159956
rect 426492 159944 426498 159996
rect 430206 159944 430212 159996
rect 430264 159984 430270 159996
rect 433058 159984 433064 159996
rect 430264 159956 433064 159984
rect 430264 159944 430270 159956
rect 433058 159944 433064 159956
rect 433116 159944 433122 159996
rect 450354 159944 450360 159996
rect 450412 159984 450418 159996
rect 456058 159984 456064 159996
rect 450412 159956 456064 159984
rect 450412 159944 450418 159956
rect 456058 159944 456064 159956
rect 456116 159944 456122 159996
rect 457898 159944 457904 159996
rect 457956 159984 457962 159996
rect 464706 159984 464712 159996
rect 457956 159956 464712 159984
rect 457956 159944 457962 159956
rect 464706 159944 464712 159956
rect 464764 159944 464770 159996
rect 76926 159876 76932 159928
rect 76984 159916 76990 159928
rect 147766 159916 147772 159928
rect 76984 159888 147772 159916
rect 76984 159876 76990 159888
rect 147766 159876 147772 159888
rect 147824 159876 147830 159928
rect 150894 159876 150900 159928
rect 150952 159916 150958 159928
rect 207014 159916 207020 159928
rect 150952 159888 207020 159916
rect 150952 159876 150958 159888
rect 207014 159876 207020 159888
rect 207072 159876 207078 159928
rect 208946 159876 208952 159928
rect 209004 159916 209010 159928
rect 220170 159916 220176 159928
rect 209004 159888 220176 159916
rect 209004 159876 209010 159888
rect 220170 159876 220176 159888
rect 220228 159876 220234 159928
rect 222378 159876 222384 159928
rect 222436 159916 222442 159928
rect 225690 159916 225696 159928
rect 222436 159888 225696 159916
rect 222436 159876 222442 159888
rect 225690 159876 225696 159888
rect 225748 159876 225754 159928
rect 238386 159876 238392 159928
rect 238444 159916 238450 159928
rect 288342 159916 288348 159928
rect 238444 159888 288348 159916
rect 238444 159876 238450 159888
rect 288342 159876 288348 159888
rect 288400 159876 288406 159928
rect 291378 159876 291384 159928
rect 291436 159916 291442 159928
rect 311894 159916 311900 159928
rect 291436 159888 311900 159916
rect 291436 159876 291442 159888
rect 311894 159876 311900 159888
rect 311952 159876 311958 159928
rect 325878 159876 325884 159928
rect 325936 159916 325942 159928
rect 362126 159916 362132 159928
rect 325936 159888 362132 159916
rect 325936 159876 325942 159888
rect 362126 159876 362132 159888
rect 362184 159876 362190 159928
rect 386414 159876 386420 159928
rect 386472 159916 386478 159928
rect 412818 159916 412824 159928
rect 386472 159888 412824 159916
rect 386472 159876 386478 159888
rect 412818 159876 412824 159888
rect 412876 159876 412882 159928
rect 86954 159808 86960 159860
rect 87012 159848 87018 159860
rect 160278 159848 160284 159860
rect 87012 159820 160284 159848
rect 87012 159808 87018 159820
rect 160278 159808 160284 159820
rect 160336 159808 160342 159860
rect 171134 159808 171140 159860
rect 171192 159848 171198 159860
rect 230382 159848 230388 159860
rect 171192 159820 230388 159848
rect 171192 159808 171198 159820
rect 230382 159808 230388 159820
rect 230440 159808 230446 159860
rect 231670 159808 231676 159860
rect 231728 159848 231734 159860
rect 284386 159848 284392 159860
rect 231728 159820 284392 159848
rect 231728 159808 231734 159820
rect 284386 159808 284392 159820
rect 284444 159808 284450 159860
rect 305638 159808 305644 159860
rect 305696 159848 305702 159860
rect 346302 159848 346308 159860
rect 305696 159820 346308 159848
rect 305696 159808 305702 159820
rect 346302 159808 346308 159820
rect 346360 159808 346366 159860
rect 375466 159808 375472 159860
rect 375524 159848 375530 159860
rect 405550 159848 405556 159860
rect 375524 159820 405556 159848
rect 375524 159808 375530 159820
rect 405550 159808 405556 159820
rect 405608 159808 405614 159860
rect 406654 159808 406660 159860
rect 406712 159848 406718 159860
rect 429378 159848 429384 159860
rect 406712 159820 429384 159848
rect 406712 159808 406718 159820
rect 429378 159808 429384 159820
rect 429436 159808 429442 159860
rect 472250 159808 472256 159860
rect 472308 159848 472314 159860
rect 479426 159848 479432 159860
rect 472308 159820 479432 159848
rect 472308 159808 472314 159820
rect 479426 159808 479432 159820
rect 479484 159808 479490 159860
rect 479794 159808 479800 159860
rect 479852 159848 479858 159860
rect 485222 159848 485228 159860
rect 479852 159820 485228 159848
rect 479852 159808 479858 159820
rect 485222 159808 485228 159820
rect 485280 159808 485286 159860
rect 60090 159740 60096 159792
rect 60148 159780 60154 159792
rect 133506 159780 133512 159792
rect 60148 159752 133512 159780
rect 60148 159740 60154 159752
rect 133506 159740 133512 159752
rect 133564 159740 133570 159792
rect 157610 159740 157616 159792
rect 157668 159780 157674 159792
rect 216766 159780 216772 159792
rect 157668 159752 216772 159780
rect 157668 159740 157674 159752
rect 216766 159740 216772 159752
rect 216824 159740 216830 159792
rect 218238 159740 218244 159792
rect 218296 159780 218302 159792
rect 272518 159780 272524 159792
rect 218296 159752 272524 159780
rect 218296 159740 218302 159752
rect 272518 159740 272524 159752
rect 272576 159740 272582 159792
rect 277946 159740 277952 159792
rect 278004 159780 278010 159792
rect 287054 159780 287060 159792
rect 278004 159752 287060 159780
rect 278004 159740 278010 159752
rect 287054 159740 287060 159752
rect 287112 159740 287118 159792
rect 287974 159740 287980 159792
rect 288032 159780 288038 159792
rect 288618 159780 288624 159792
rect 288032 159752 288624 159780
rect 288032 159740 288038 159752
rect 288618 159740 288624 159752
rect 288676 159740 288682 159792
rect 298922 159740 298928 159792
rect 298980 159780 298986 159792
rect 343634 159780 343640 159792
rect 298980 159752 343640 159780
rect 298980 159740 298986 159752
rect 343634 159740 343640 159752
rect 343692 159740 343698 159792
rect 366266 159740 366272 159792
rect 366324 159780 366330 159792
rect 398466 159780 398472 159792
rect 366324 159752 398472 159780
rect 366324 159740 366330 159752
rect 398466 159740 398472 159752
rect 398524 159740 398530 159792
rect 399846 159740 399852 159792
rect 399904 159780 399910 159792
rect 424226 159780 424232 159792
rect 399904 159752 424232 159780
rect 399904 159740 399910 159752
rect 424226 159740 424232 159752
rect 424284 159740 424290 159792
rect 451182 159740 451188 159792
rect 451240 159780 451246 159792
rect 462866 159780 462872 159792
rect 451240 159752 462872 159780
rect 451240 159740 451246 159752
rect 462866 159740 462872 159752
rect 462924 159740 462930 159792
rect 463786 159740 463792 159792
rect 463844 159780 463850 159792
rect 471790 159780 471796 159792
rect 463844 159752 471796 159780
rect 463844 159740 463850 159752
rect 471790 159740 471796 159752
rect 471848 159740 471854 159792
rect 478966 159740 478972 159792
rect 479024 159780 479030 159792
rect 484578 159780 484584 159792
rect 479024 159752 484584 159780
rect 479024 159740 479030 159752
rect 484578 159740 484584 159752
rect 484636 159740 484642 159792
rect 46566 159672 46572 159724
rect 46624 159712 46630 159724
rect 120166 159712 120172 159724
rect 46624 159684 120172 159712
rect 46624 159672 46630 159684
rect 120166 159672 120172 159684
rect 120224 159672 120230 159724
rect 124030 159672 124036 159724
rect 124088 159712 124094 159724
rect 187694 159712 187700 159724
rect 124088 159684 187700 159712
rect 124088 159672 124094 159684
rect 187694 159672 187700 159684
rect 187752 159672 187758 159724
rect 194686 159672 194692 159724
rect 194744 159712 194750 159724
rect 213638 159712 213644 159724
rect 194744 159684 213644 159712
rect 194744 159672 194750 159684
rect 213638 159672 213644 159684
rect 213696 159672 213702 159724
rect 214834 159672 214840 159724
rect 214892 159712 214898 159724
rect 224586 159712 224592 159724
rect 214892 159684 224592 159712
rect 214892 159672 214898 159684
rect 224586 159672 224592 159684
rect 224644 159672 224650 159724
rect 224954 159672 224960 159724
rect 225012 159712 225018 159724
rect 281442 159712 281448 159724
rect 225012 159684 281448 159712
rect 225012 159672 225018 159684
rect 281442 159672 281448 159684
rect 281500 159672 281506 159724
rect 282086 159672 282092 159724
rect 282144 159712 282150 159724
rect 289906 159712 289912 159724
rect 282144 159684 289912 159712
rect 282144 159672 282150 159684
rect 289906 159672 289912 159684
rect 289964 159672 289970 159724
rect 292206 159672 292212 159724
rect 292264 159712 292270 159724
rect 338758 159712 338764 159724
rect 292264 159684 338764 159712
rect 292264 159672 292270 159684
rect 338758 159672 338764 159684
rect 338816 159672 338822 159724
rect 352742 159672 352748 159724
rect 352800 159712 352806 159724
rect 385954 159712 385960 159724
rect 352800 159684 385960 159712
rect 352800 159672 352806 159684
rect 385954 159672 385960 159684
rect 386012 159672 386018 159724
rect 388990 159672 388996 159724
rect 389048 159712 389054 159724
rect 414290 159712 414296 159724
rect 389048 159684 414296 159712
rect 389048 159672 389054 159684
rect 414290 159672 414296 159684
rect 414348 159672 414354 159724
rect 420086 159672 420092 159724
rect 420144 159712 420150 159724
rect 435818 159712 435824 159724
rect 420144 159684 435824 159712
rect 420144 159672 420150 159684
rect 435818 159672 435824 159684
rect 435876 159672 435882 159724
rect 458726 159672 458732 159724
rect 458784 159712 458790 159724
rect 465074 159712 465080 159724
rect 458784 159684 465080 159712
rect 458784 159672 458790 159684
rect 465074 159672 465080 159684
rect 465132 159672 465138 159724
rect 53374 159604 53380 159656
rect 53432 159644 53438 159656
rect 128354 159644 128360 159656
rect 53432 159616 128360 159644
rect 53432 159604 53438 159616
rect 128354 159604 128360 159616
rect 128412 159604 128418 159656
rect 130746 159604 130752 159656
rect 130804 159644 130810 159656
rect 195238 159644 195244 159656
rect 130804 159616 195244 159644
rect 130804 159604 130810 159616
rect 195238 159604 195244 159616
rect 195296 159604 195302 159656
rect 211430 159604 211436 159656
rect 211488 159644 211494 159656
rect 268930 159644 268936 159656
rect 211488 159616 268936 159644
rect 211488 159604 211494 159616
rect 268930 159604 268936 159616
rect 268988 159604 268994 159656
rect 285490 159604 285496 159656
rect 285548 159644 285554 159656
rect 332594 159644 332600 159656
rect 285548 159616 332600 159644
rect 285548 159604 285554 159616
rect 332594 159604 332600 159616
rect 332652 159604 332658 159656
rect 346026 159604 346032 159656
rect 346084 159644 346090 159656
rect 378134 159644 378140 159656
rect 346084 159616 378140 159644
rect 346084 159604 346090 159616
rect 378134 159604 378140 159616
rect 378192 159604 378198 159656
rect 382182 159604 382188 159656
rect 382240 159644 382246 159656
rect 408494 159644 408500 159656
rect 382240 159616 408500 159644
rect 382240 159604 382246 159616
rect 408494 159604 408500 159616
rect 408552 159604 408558 159656
rect 413370 159604 413376 159656
rect 413428 159644 413434 159656
rect 434438 159644 434444 159656
rect 413428 159616 434444 159644
rect 413428 159604 413434 159616
rect 434438 159604 434444 159616
rect 434496 159604 434502 159656
rect 441062 159604 441068 159656
rect 441120 159644 441126 159656
rect 445662 159644 445668 159656
rect 441120 159616 445668 159644
rect 441120 159604 441126 159616
rect 445662 159604 445668 159616
rect 445720 159604 445726 159656
rect 447870 159604 447876 159656
rect 447928 159644 447934 159656
rect 460198 159644 460204 159656
rect 447928 159616 460204 159644
rect 447928 159604 447934 159616
rect 460198 159604 460204 159616
rect 460256 159604 460262 159656
rect 468018 159604 468024 159656
rect 468076 159644 468082 159656
rect 476022 159644 476028 159656
rect 468076 159616 476028 159644
rect 468076 159604 468082 159616
rect 476022 159604 476028 159616
rect 476080 159604 476086 159656
rect 80238 159536 80244 159588
rect 80296 159576 80302 159588
rect 158438 159576 158444 159588
rect 80296 159548 158444 159576
rect 80296 159536 80302 159548
rect 158438 159536 158444 159548
rect 158496 159536 158502 159588
rect 170214 159536 170220 159588
rect 170272 159576 170278 159588
rect 176654 159576 176660 159588
rect 170272 159548 176660 159576
rect 170272 159536 170278 159548
rect 176654 159536 176660 159548
rect 176712 159536 176718 159588
rect 197998 159536 198004 159588
rect 198056 159576 198062 159588
rect 259638 159576 259644 159588
rect 198056 159548 259644 159576
rect 198056 159536 198062 159548
rect 259638 159536 259644 159548
rect 259696 159536 259702 159588
rect 272058 159536 272064 159588
rect 272116 159576 272122 159588
rect 320726 159576 320732 159588
rect 272116 159548 320732 159576
rect 272116 159536 272122 159548
rect 320726 159536 320732 159548
rect 320784 159536 320790 159588
rect 339310 159536 339316 159588
rect 339368 159576 339374 159588
rect 377950 159576 377956 159588
rect 339368 159548 377956 159576
rect 339368 159536 339374 159548
rect 377950 159536 377956 159548
rect 378008 159536 378014 159588
rect 379698 159536 379704 159588
rect 379756 159576 379762 159588
rect 408770 159576 408776 159588
rect 379756 159548 408776 159576
rect 379756 159536 379762 159548
rect 408770 159536 408776 159548
rect 408828 159536 408834 159588
rect 431862 159536 431868 159588
rect 431920 159576 431926 159588
rect 436370 159576 436376 159588
rect 431920 159548 436376 159576
rect 431920 159536 431926 159548
rect 436370 159536 436376 159548
rect 436428 159536 436434 159588
rect 449526 159536 449532 159588
rect 449584 159576 449590 159588
rect 461486 159576 461492 159588
rect 449584 159548 461492 159576
rect 449584 159536 449590 159548
rect 461486 159536 461492 159548
rect 461544 159536 461550 159588
rect 470502 159536 470508 159588
rect 470560 159576 470566 159588
rect 476114 159576 476120 159588
rect 470560 159548 476120 159576
rect 470560 159536 470566 159548
rect 476114 159536 476120 159548
rect 476172 159536 476178 159588
rect 100478 159468 100484 159520
rect 100536 159508 100542 159520
rect 179414 159508 179420 159520
rect 100536 159480 179420 159508
rect 100536 159468 100542 159480
rect 179414 159468 179420 159480
rect 179472 159468 179478 159520
rect 184566 159468 184572 159520
rect 184624 159508 184630 159520
rect 247218 159508 247224 159520
rect 184624 159480 247224 159508
rect 184624 159468 184630 159480
rect 247218 159468 247224 159480
rect 247276 159468 247282 159520
rect 251818 159468 251824 159520
rect 251876 159508 251882 159520
rect 301682 159508 301688 159520
rect 251876 159480 301688 159508
rect 251876 159468 251882 159480
rect 301682 159468 301688 159480
rect 301740 159468 301746 159520
rect 308214 159468 308220 159520
rect 308272 159508 308278 159520
rect 317782 159508 317788 159520
rect 308272 159480 317788 159508
rect 308272 159468 308278 159480
rect 317782 159468 317788 159480
rect 317840 159468 317846 159520
rect 319162 159468 319168 159520
rect 319220 159508 319226 159520
rect 361574 159508 361580 159520
rect 319220 159480 361580 159508
rect 319220 159468 319226 159480
rect 361574 159468 361580 159480
rect 361632 159468 361638 159520
rect 368750 159468 368756 159520
rect 368808 159508 368814 159520
rect 400398 159508 400404 159520
rect 368808 159480 400404 159508
rect 368808 159468 368814 159480
rect 400398 159468 400404 159480
rect 400456 159468 400462 159520
rect 402422 159468 402428 159520
rect 402480 159508 402486 159520
rect 426158 159508 426164 159520
rect 402480 159480 426164 159508
rect 402480 159468 402486 159480
rect 426158 159468 426164 159480
rect 426216 159468 426222 159520
rect 433518 159468 433524 159520
rect 433576 159508 433582 159520
rect 449802 159508 449808 159520
rect 433576 159480 449808 159508
rect 433576 159468 433582 159480
rect 449802 159468 449808 159480
rect 449860 159468 449866 159520
rect 453758 159468 453764 159520
rect 453816 159508 453822 159520
rect 465258 159508 465264 159520
rect 453816 159480 465264 159508
rect 453816 159468 453822 159480
rect 465258 159468 465264 159480
rect 465316 159468 465322 159520
rect 467190 159468 467196 159520
rect 467248 159508 467254 159520
rect 473354 159508 473360 159520
rect 467248 159480 473360 159508
rect 467248 159468 467254 159480
rect 473354 159468 473360 159480
rect 473412 159468 473418 159520
rect 482278 159468 482284 159520
rect 482336 159508 482342 159520
rect 487246 159508 487252 159520
rect 482336 159480 487252 159508
rect 482336 159468 482342 159480
rect 487246 159468 487252 159480
rect 487304 159468 487310 159520
rect 26418 159400 26424 159452
rect 26476 159440 26482 159452
rect 129826 159440 129832 159452
rect 26476 159412 129832 159440
rect 26476 159400 26482 159412
rect 129826 159400 129832 159412
rect 129884 159400 129890 159452
rect 139118 159400 139124 159452
rect 139176 159440 139182 159452
rect 157334 159440 157340 159452
rect 139176 159412 157340 159440
rect 139176 159400 139182 159412
rect 157334 159400 157340 159412
rect 157392 159400 157398 159452
rect 177850 159400 177856 159452
rect 177908 159440 177914 159452
rect 241698 159440 241704 159452
rect 177908 159412 241704 159440
rect 177908 159400 177914 159412
rect 241698 159400 241704 159412
rect 241756 159400 241762 159452
rect 245102 159400 245108 159452
rect 245160 159440 245166 159452
rect 298738 159440 298744 159452
rect 245160 159412 298744 159440
rect 245160 159400 245166 159412
rect 298738 159400 298744 159412
rect 298796 159400 298802 159452
rect 312446 159400 312452 159452
rect 312504 159440 312510 159452
rect 355226 159440 355232 159452
rect 312504 159412 355232 159440
rect 312504 159400 312510 159412
rect 355226 159400 355232 159412
rect 355284 159400 355290 159452
rect 359550 159400 359556 159452
rect 359608 159440 359614 159452
rect 393406 159440 393412 159452
rect 359608 159412 393412 159440
rect 359608 159400 359614 159412
rect 393406 159400 393412 159412
rect 393464 159400 393470 159452
rect 395706 159400 395712 159452
rect 395764 159440 395770 159452
rect 421098 159440 421104 159452
rect 395764 159412 421104 159440
rect 395764 159400 395770 159412
rect 421098 159400 421104 159412
rect 421156 159400 421162 159452
rect 432690 159400 432696 159452
rect 432748 159440 432754 159452
rect 447134 159440 447140 159452
rect 432748 159412 447140 159440
rect 432748 159400 432754 159412
rect 447134 159400 447140 159412
rect 447192 159400 447198 159452
rect 448698 159400 448704 159452
rect 448756 159440 448762 159452
rect 460934 159440 460940 159452
rect 448756 159412 460940 159440
rect 448756 159400 448762 159412
rect 460934 159400 460940 159412
rect 460992 159400 460998 159452
rect 468846 159400 468852 159452
rect 468904 159440 468910 159452
rect 474826 159440 474832 159452
rect 468904 159412 474832 159440
rect 468904 159400 468910 159412
rect 474826 159400 474832 159412
rect 474884 159400 474890 159452
rect 477310 159400 477316 159452
rect 477368 159440 477374 159452
rect 483290 159440 483296 159452
rect 477368 159412 483296 159440
rect 477368 159400 477374 159412
rect 483290 159400 483296 159412
rect 483348 159400 483354 159452
rect 518066 159400 518072 159452
rect 518124 159440 518130 159452
rect 522666 159440 522672 159452
rect 518124 159412 522672 159440
rect 518124 159400 518130 159412
rect 522666 159400 522672 159412
rect 522724 159400 522730 159452
rect 12986 159332 12992 159384
rect 13044 159372 13050 159384
rect 123938 159372 123944 159384
rect 13044 159344 123944 159372
rect 13044 159332 13050 159344
rect 123938 159332 123944 159344
rect 123996 159332 124002 159384
rect 132402 159332 132408 159384
rect 132460 159372 132466 159384
rect 136082 159372 136088 159384
rect 132460 159344 136088 159372
rect 132460 159332 132466 159344
rect 136082 159332 136088 159344
rect 136140 159332 136146 159384
rect 140774 159332 140780 159384
rect 140832 159372 140838 159384
rect 173986 159372 173992 159384
rect 140832 159344 173992 159372
rect 140832 159332 140838 159344
rect 173986 159332 173992 159344
rect 174044 159332 174050 159384
rect 191282 159332 191288 159384
rect 191340 159372 191346 159384
rect 257338 159372 257344 159384
rect 191340 159344 257344 159372
rect 191340 159332 191346 159344
rect 257338 159332 257344 159344
rect 257396 159332 257402 159384
rect 287054 159332 287060 159384
rect 287112 159372 287118 159384
rect 291470 159372 291476 159384
rect 287112 159344 291476 159372
rect 287112 159332 287118 159344
rect 291470 159332 291476 159344
rect 291528 159332 291534 159384
rect 331766 159332 331772 159384
rect 331824 159372 331830 159384
rect 372062 159372 372068 159384
rect 331824 159344 372068 159372
rect 331824 159332 331830 159344
rect 372062 159332 372068 159344
rect 372120 159332 372126 159384
rect 372982 159332 372988 159384
rect 373040 159372 373046 159384
rect 403158 159372 403164 159384
rect 373040 159344 403164 159372
rect 373040 159332 373046 159344
rect 403158 159332 403164 159344
rect 403216 159332 403222 159384
rect 426802 159332 426808 159384
rect 426860 159372 426866 159384
rect 433242 159372 433248 159384
rect 426860 159344 433248 159372
rect 426860 159332 426866 159344
rect 433242 159332 433248 159344
rect 433300 159332 433306 159384
rect 434346 159332 434352 159384
rect 434404 159372 434410 159384
rect 450078 159372 450084 159384
rect 434404 159344 450084 159372
rect 434404 159332 434410 159344
rect 450078 159332 450084 159344
rect 450136 159332 450142 159384
rect 452010 159332 452016 159384
rect 452068 159372 452074 159384
rect 463970 159372 463976 159384
rect 452068 159344 463976 159372
rect 452068 159332 452074 159344
rect 463970 159332 463976 159344
rect 464028 159332 464034 159384
rect 469674 159332 469680 159384
rect 469732 159372 469738 159384
rect 477402 159372 477408 159384
rect 469732 159344 477408 159372
rect 469732 159332 469738 159344
rect 477402 159332 477408 159344
rect 477460 159332 477466 159384
rect 478138 159332 478144 159384
rect 478196 159372 478202 159384
rect 483934 159372 483940 159384
rect 478196 159344 483940 159372
rect 478196 159332 478202 159344
rect 483934 159332 483940 159344
rect 483992 159332 483998 159384
rect 518710 159332 518716 159384
rect 518768 159372 518774 159384
rect 523494 159372 523500 159384
rect 518768 159344 523500 159372
rect 518768 159332 518774 159344
rect 523494 159332 523500 159344
rect 523552 159332 523558 159384
rect 93670 159264 93676 159316
rect 93728 159304 93734 159316
rect 146018 159304 146024 159316
rect 93728 159276 146024 159304
rect 93728 159264 93734 159276
rect 146018 159264 146024 159276
rect 146076 159264 146082 159316
rect 181162 159264 181168 159316
rect 181220 159304 181226 159316
rect 230658 159304 230664 159316
rect 181220 159276 230664 159304
rect 181220 159264 181226 159276
rect 230658 159264 230664 159276
rect 230716 159264 230722 159316
rect 237558 159264 237564 159316
rect 237616 159304 237622 159316
rect 251726 159304 251732 159316
rect 237616 159276 251732 159304
rect 237616 159264 237622 159276
rect 251726 159264 251732 159276
rect 251784 159264 251790 159316
rect 271230 159264 271236 159316
rect 271288 159304 271294 159316
rect 296806 159304 296812 159316
rect 271288 159276 296812 159304
rect 271288 159264 271294 159276
rect 296806 159264 296812 159276
rect 296864 159264 296870 159316
rect 298094 159264 298100 159316
rect 298152 159304 298158 159316
rect 311986 159304 311992 159316
rect 298152 159276 311992 159304
rect 298152 159264 298158 159276
rect 311986 159264 311992 159276
rect 312044 159264 312050 159316
rect 325050 159264 325056 159316
rect 325108 159304 325114 159316
rect 352006 159304 352012 159316
rect 325108 159276 352012 159304
rect 325108 159264 325114 159276
rect 352006 159264 352012 159276
rect 352064 159264 352070 159316
rect 461302 159264 461308 159316
rect 461360 159304 461366 159316
rect 467926 159304 467932 159316
rect 461360 159276 467932 159304
rect 461360 159264 461366 159276
rect 467926 159264 467932 159276
rect 467984 159264 467990 159316
rect 109678 159196 109684 159248
rect 109736 159236 109742 159248
rect 118694 159236 118700 159248
rect 109736 159208 118700 159236
rect 109736 159196 109742 159208
rect 118694 159196 118700 159208
rect 118752 159196 118758 159248
rect 144178 159196 144184 159248
rect 144236 159236 144242 159248
rect 192570 159236 192576 159248
rect 144236 159208 192576 159236
rect 144236 159196 144242 159208
rect 192570 159196 192576 159208
rect 192628 159196 192634 159248
rect 208118 159196 208124 159248
rect 208176 159236 208182 159248
rect 222102 159236 222108 159248
rect 208176 159208 222108 159236
rect 208176 159196 208182 159208
rect 222102 159196 222108 159208
rect 222160 159196 222166 159248
rect 227438 159196 227444 159248
rect 227496 159236 227502 159248
rect 247034 159236 247040 159248
rect 227496 159208 247040 159236
rect 227496 159196 227502 159208
rect 247034 159196 247040 159208
rect 247092 159196 247098 159248
rect 250990 159196 250996 159248
rect 251048 159236 251054 159248
rect 274634 159236 274640 159248
rect 251048 159208 274640 159236
rect 251048 159196 251054 159208
rect 274634 159196 274640 159208
rect 274692 159196 274698 159248
rect 284662 159196 284668 159248
rect 284720 159236 284726 159248
rect 305454 159236 305460 159248
rect 284720 159208 305460 159236
rect 284720 159196 284726 159208
rect 305454 159196 305460 159208
rect 305512 159196 305518 159248
rect 460474 159196 460480 159248
rect 460532 159236 460538 159248
rect 466638 159236 466644 159248
rect 460532 159208 466644 159236
rect 460532 159196 460538 159208
rect 466638 159196 466644 159208
rect 466696 159196 466702 159248
rect 110506 159128 110512 159180
rect 110564 159168 110570 159180
rect 146110 159168 146116 159180
rect 110564 159140 146116 159168
rect 110564 159128 110570 159140
rect 146110 159128 146116 159140
rect 146168 159128 146174 159180
rect 155954 159128 155960 159180
rect 156012 159168 156018 159180
rect 197630 159168 197636 159180
rect 156012 159140 197636 159168
rect 156012 159128 156018 159140
rect 197630 159128 197636 159140
rect 197688 159128 197694 159180
rect 201402 159128 201408 159180
rect 201460 159168 201466 159180
rect 211890 159168 211896 159180
rect 201460 159140 211896 159168
rect 201460 159128 201466 159140
rect 211890 159128 211896 159140
rect 211948 159128 211954 159180
rect 257706 159128 257712 159180
rect 257764 159168 257770 159180
rect 280062 159168 280068 159180
rect 257764 159140 280068 159168
rect 257764 159128 257770 159140
rect 280062 159128 280068 159140
rect 280120 159128 280126 159180
rect 304810 159128 304816 159180
rect 304868 159168 304874 159180
rect 324314 159168 324320 159180
rect 304868 159140 324320 159168
rect 304868 159128 304874 159140
rect 324314 159128 324320 159140
rect 324372 159128 324378 159180
rect 446122 159128 446128 159180
rect 446180 159168 446186 159180
rect 458358 159168 458364 159180
rect 446180 159140 458364 159168
rect 446180 159128 446186 159140
rect 458358 159128 458364 159140
rect 458416 159128 458422 159180
rect 462958 159128 462964 159180
rect 463016 159168 463022 159180
rect 469214 159168 469220 159180
rect 463016 159140 469220 159168
rect 463016 159128 463022 159140
rect 469214 159128 469220 159140
rect 469272 159128 469278 159180
rect 37366 159060 37372 159112
rect 37424 159100 37430 159112
rect 38562 159100 38568 159112
rect 37424 159072 38568 159100
rect 37424 159060 37430 159072
rect 38562 159060 38568 159072
rect 38620 159060 38626 159112
rect 91186 159060 91192 159112
rect 91244 159100 91250 159112
rect 92382 159100 92388 159112
rect 91244 159072 92388 159100
rect 91244 159060 91250 159072
rect 92382 159060 92388 159072
rect 92440 159060 92446 159112
rect 127342 159060 127348 159112
rect 127400 159100 127406 159112
rect 147674 159100 147680 159112
rect 127400 159072 147680 159100
rect 127400 159060 127406 159072
rect 147674 159060 147680 159072
rect 147732 159060 147738 159112
rect 174446 159060 174452 159112
rect 174504 159100 174510 159112
rect 202966 159100 202972 159112
rect 174504 159072 202972 159100
rect 174504 159060 174510 159072
rect 202966 159060 202972 159072
rect 203024 159060 203030 159112
rect 214006 159060 214012 159112
rect 214064 159100 214070 159112
rect 216674 159100 216680 159112
rect 214064 159072 216680 159100
rect 214064 159060 214070 159072
rect 216674 159060 216680 159072
rect 216732 159060 216738 159112
rect 247678 159060 247684 159112
rect 247736 159100 247742 159112
rect 262122 159100 262128 159112
rect 247736 159072 262128 159100
rect 247736 159060 247742 159072
rect 262122 159060 262128 159072
rect 262180 159060 262186 159112
rect 264422 159060 264428 159112
rect 264480 159100 264486 159112
rect 284294 159100 284300 159112
rect 264480 159072 284300 159100
rect 264480 159060 264486 159072
rect 284294 159060 284300 159072
rect 284352 159060 284358 159112
rect 459646 159060 459652 159112
rect 459704 159100 459710 159112
rect 466454 159100 466460 159112
rect 459704 159072 466460 159100
rect 459704 159060 459710 159072
rect 466454 159060 466460 159072
rect 466512 159060 466518 159112
rect 471422 159060 471428 159112
rect 471480 159100 471486 159112
rect 477678 159100 477684 159112
rect 471480 159072 477684 159100
rect 471480 159060 471486 159072
rect 477678 159060 477684 159072
rect 477736 159060 477742 159112
rect 210602 158992 210608 159044
rect 210660 159032 210666 159044
rect 215018 159032 215024 159044
rect 210660 159004 215024 159032
rect 210660 158992 210666 159004
rect 215018 158992 215024 159004
rect 215076 158992 215082 159044
rect 267826 158992 267832 159044
rect 267884 159032 267890 159044
rect 279510 159032 279516 159044
rect 267884 159004 279516 159032
rect 267884 158992 267890 159004
rect 279510 158992 279516 159004
rect 279568 158992 279574 159044
rect 288894 158992 288900 159044
rect 288952 159032 288958 159044
rect 292298 159032 292304 159044
rect 288952 159004 292304 159032
rect 288952 158992 288958 159004
rect 292298 158992 292304 159004
rect 292356 158992 292362 159044
rect 455414 158992 455420 159044
rect 455472 159032 455478 159044
rect 462958 159032 462964 159044
rect 455472 159004 462964 159032
rect 455472 158992 455478 159004
rect 462958 158992 462964 159004
rect 463016 158992 463022 159044
rect 473906 158992 473912 159044
rect 473964 159032 473970 159044
rect 480714 159032 480720 159044
rect 473964 159004 480720 159032
rect 473964 158992 473970 159004
rect 480714 158992 480720 159004
rect 480772 158992 480778 159044
rect 507118 158992 507124 159044
rect 507176 159032 507182 159044
rect 508406 159032 508412 159044
rect 507176 159004 508412 159032
rect 507176 158992 507182 159004
rect 508406 158992 508412 159004
rect 508464 158992 508470 159044
rect 118970 158924 118976 158976
rect 119028 158964 119034 158976
rect 125502 158964 125508 158976
rect 119028 158936 125508 158964
rect 119028 158924 119034 158936
rect 125502 158924 125508 158936
rect 125560 158924 125566 158976
rect 224126 158924 224132 158976
rect 224184 158964 224190 158976
rect 227714 158964 227720 158976
rect 224184 158936 227720 158964
rect 224184 158924 224190 158936
rect 227714 158924 227720 158936
rect 227772 158924 227778 158976
rect 278774 158924 278780 158976
rect 278832 158964 278838 158976
rect 278832 158936 316034 158964
rect 278832 158924 278838 158936
rect 275370 158856 275376 158908
rect 275428 158896 275434 158908
rect 278314 158896 278320 158908
rect 275428 158868 278320 158896
rect 275428 158856 275434 158868
rect 278314 158856 278320 158868
rect 278372 158856 278378 158908
rect 316006 158896 316034 158936
rect 327534 158924 327540 158976
rect 327592 158964 327598 158976
rect 328362 158964 328368 158976
rect 327592 158936 328368 158964
rect 327592 158924 327598 158936
rect 328362 158924 328368 158936
rect 328420 158924 328426 158976
rect 362034 158924 362040 158976
rect 362092 158964 362098 158976
rect 366818 158964 366824 158976
rect 362092 158936 366824 158964
rect 362092 158924 362098 158936
rect 366818 158924 366824 158936
rect 366876 158924 366882 158976
rect 372154 158924 372160 158976
rect 372212 158964 372218 158976
rect 374270 158964 374276 158976
rect 372212 158936 374276 158964
rect 372212 158924 372218 158936
rect 374270 158924 374276 158936
rect 374328 158924 374334 158976
rect 405734 158924 405740 158976
rect 405792 158964 405798 158976
rect 407022 158964 407028 158976
rect 405792 158936 407028 158964
rect 405792 158924 405798 158936
rect 407022 158924 407028 158936
rect 407080 158924 407086 158976
rect 437750 158924 437756 158976
rect 437808 158964 437814 158976
rect 444282 158964 444288 158976
rect 437808 158936 444288 158964
rect 437808 158924 437814 158936
rect 444282 158924 444288 158936
rect 444340 158924 444346 158976
rect 454586 158924 454592 158976
rect 454644 158964 454650 158976
rect 461578 158964 461584 158976
rect 454644 158936 461584 158964
rect 454644 158924 454650 158936
rect 461578 158924 461584 158936
rect 461636 158924 461642 158976
rect 466362 158924 466368 158976
rect 466420 158964 466426 158976
rect 472802 158964 472808 158976
rect 466420 158936 472808 158964
rect 466420 158924 466426 158936
rect 472802 158924 472808 158936
rect 472860 158924 472866 158976
rect 475562 158924 475568 158976
rect 475620 158964 475626 158976
rect 482002 158964 482008 158976
rect 475620 158936 482008 158964
rect 475620 158924 475626 158936
rect 482002 158924 482008 158936
rect 482060 158924 482066 158976
rect 331766 158896 331772 158908
rect 316006 158868 331772 158896
rect 331766 158856 331772 158868
rect 331824 158856 331830 158908
rect 456242 158856 456248 158908
rect 456300 158896 456306 158908
rect 463142 158896 463148 158908
rect 456300 158868 463148 158896
rect 456300 158856 456306 158868
rect 463142 158856 463148 158868
rect 463200 158856 463206 158908
rect 465534 158856 465540 158908
rect 465592 158896 465598 158908
rect 471974 158896 471980 158908
rect 465592 158868 471980 158896
rect 465592 158856 465598 158868
rect 471974 158856 471980 158868
rect 472032 158856 472038 158908
rect 474734 158856 474740 158908
rect 474792 158896 474798 158908
rect 480254 158896 480260 158908
rect 474792 158868 480260 158896
rect 474792 158856 474798 158868
rect 480254 158856 480260 158868
rect 480312 158856 480318 158908
rect 480622 158856 480628 158908
rect 480680 158896 480686 158908
rect 485958 158896 485964 158908
rect 480680 158868 485964 158896
rect 480680 158856 480686 158868
rect 485958 158856 485964 158868
rect 486016 158856 486022 158908
rect 508406 158856 508412 158908
rect 508464 158896 508470 158908
rect 510062 158896 510068 158908
rect 508464 158868 510068 158896
rect 508464 158856 508470 158868
rect 510062 158856 510068 158868
rect 510120 158856 510126 158908
rect 145834 158788 145840 158840
rect 145892 158828 145898 158840
rect 150434 158828 150440 158840
rect 145892 158800 150440 158828
rect 145892 158788 145898 158800
rect 150434 158788 150440 158800
rect 150492 158788 150498 158840
rect 196342 158788 196348 158840
rect 196400 158828 196406 158840
rect 198734 158828 198740 158840
rect 196400 158800 198740 158828
rect 196400 158788 196406 158800
rect 198734 158788 198740 158800
rect 198792 158788 198798 158840
rect 261938 158788 261944 158840
rect 261996 158828 262002 158840
rect 263410 158828 263416 158840
rect 261996 158800 263416 158828
rect 261996 158788 262002 158800
rect 263410 158788 263416 158800
rect 263468 158788 263474 158840
rect 268654 158788 268660 158840
rect 268712 158828 268718 158840
rect 271690 158828 271696 158840
rect 268712 158800 271696 158828
rect 268712 158788 268718 158800
rect 271690 158788 271696 158800
rect 271748 158788 271754 158840
rect 315758 158788 315764 158840
rect 315816 158828 315822 158840
rect 318702 158828 318708 158840
rect 315816 158800 318708 158828
rect 315816 158788 315822 158800
rect 318702 158788 318708 158800
rect 318760 158788 318766 158840
rect 335998 158788 336004 158840
rect 336056 158828 336062 158840
rect 337930 158828 337936 158840
rect 336056 158800 337936 158828
rect 336056 158788 336062 158800
rect 337930 158788 337936 158800
rect 337988 158788 337994 158840
rect 436094 158788 436100 158840
rect 436152 158828 436158 158840
rect 438854 158828 438860 158840
rect 436152 158800 438860 158828
rect 436152 158788 436158 158800
rect 438854 158788 438860 158800
rect 438912 158788 438918 158840
rect 464614 158788 464620 158840
rect 464672 158828 464678 158840
rect 471606 158828 471612 158840
rect 464672 158800 471612 158828
rect 464672 158788 464678 158800
rect 471606 158788 471612 158800
rect 471664 158788 471670 158840
rect 476390 158788 476396 158840
rect 476448 158828 476454 158840
rect 481634 158828 481640 158840
rect 476448 158800 481640 158828
rect 476448 158788 476454 158800
rect 481634 158788 481640 158800
rect 481692 158788 481698 158840
rect 499942 158788 499948 158840
rect 500000 158828 500006 158840
rect 500586 158828 500592 158840
rect 500000 158800 500592 158828
rect 500000 158788 500006 158800
rect 500586 158788 500592 158800
rect 500644 158788 500650 158840
rect 506382 158788 506388 158840
rect 506440 158828 506446 158840
rect 507578 158828 507584 158840
rect 506440 158800 507584 158828
rect 506440 158788 506446 158800
rect 507578 158788 507584 158800
rect 507636 158788 507642 158840
rect 382 158720 388 158772
rect 440 158760 446 158772
rect 2038 158760 2044 158772
rect 440 158732 2044 158760
rect 440 158720 446 158732
rect 2038 158720 2044 158732
rect 2096 158720 2102 158772
rect 64230 158720 64236 158772
rect 64288 158760 64294 158772
rect 64782 158760 64788 158772
rect 64288 158732 64788 158760
rect 64288 158720 64294 158732
rect 64782 158720 64788 158732
rect 64840 158720 64846 158772
rect 71038 158720 71044 158772
rect 71096 158760 71102 158772
rect 71682 158760 71688 158772
rect 71096 158732 71688 158760
rect 71096 158720 71102 158732
rect 71682 158720 71688 158732
rect 71740 158720 71746 158772
rect 77754 158720 77760 158772
rect 77812 158760 77818 158772
rect 78582 158760 78588 158772
rect 77812 158732 78588 158760
rect 77812 158720 77818 158732
rect 78582 158720 78588 158732
rect 78640 158720 78646 158772
rect 84470 158720 84476 158772
rect 84528 158760 84534 158772
rect 85482 158760 85488 158772
rect 84528 158732 85488 158760
rect 84528 158720 84534 158732
rect 85482 158720 85488 158732
rect 85540 158720 85546 158772
rect 103790 158720 103796 158772
rect 103848 158760 103854 158772
rect 109034 158760 109040 158772
rect 103848 158732 109040 158760
rect 103848 158720 103854 158732
rect 109034 158720 109040 158732
rect 109092 158720 109098 158772
rect 121454 158720 121460 158772
rect 121512 158760 121518 158772
rect 122742 158760 122748 158772
rect 121512 158732 122748 158760
rect 121512 158720 121518 158732
rect 122742 158720 122748 158732
rect 122800 158720 122806 158772
rect 128998 158720 129004 158772
rect 129056 158760 129062 158772
rect 131114 158760 131120 158772
rect 129056 158732 131120 158760
rect 129056 158720 129062 158732
rect 131114 158720 131120 158732
rect 131172 158720 131178 158772
rect 131574 158720 131580 158772
rect 131632 158760 131638 158772
rect 132402 158760 132408 158772
rect 131632 158732 132408 158760
rect 131632 158720 131638 158732
rect 132402 158720 132408 158732
rect 132460 158720 132466 158772
rect 145006 158720 145012 158772
rect 145064 158760 145070 158772
rect 146202 158760 146208 158772
rect 145064 158732 146208 158760
rect 145064 158720 145070 158732
rect 146202 158720 146208 158732
rect 146260 158720 146266 158772
rect 152550 158720 152556 158772
rect 152608 158760 152614 158772
rect 153102 158760 153108 158772
rect 152608 158732 153108 158760
rect 152608 158720 152614 158732
rect 153102 158720 153108 158732
rect 153160 158720 153166 158772
rect 165246 158720 165252 158772
rect 165304 158760 165310 158772
rect 167638 158760 167644 158772
rect 165304 158732 167644 158760
rect 165304 158720 165310 158732
rect 167638 158720 167644 158732
rect 167696 158720 167702 158772
rect 202230 158720 202236 158772
rect 202288 158760 202294 158772
rect 202782 158760 202788 158772
rect 202288 158732 202788 158760
rect 202288 158720 202294 158732
rect 202782 158720 202788 158732
rect 202840 158720 202846 158772
rect 203058 158720 203064 158772
rect 203116 158760 203122 158772
rect 208486 158760 208492 158772
rect 203116 158732 208492 158760
rect 203116 158720 203122 158732
rect 208486 158720 208492 158732
rect 208544 158720 208550 158772
rect 220722 158720 220728 158772
rect 220780 158760 220786 158772
rect 227898 158760 227904 158772
rect 220780 158732 227904 158760
rect 220780 158720 220786 158732
rect 227898 158720 227904 158732
rect 227956 158720 227962 158772
rect 230842 158720 230848 158772
rect 230900 158760 230906 158772
rect 238662 158760 238668 158772
rect 230900 158732 238668 158760
rect 230900 158720 230906 158732
rect 238662 158720 238668 158732
rect 238720 158720 238726 158772
rect 241790 158720 241796 158772
rect 241848 158760 241854 158772
rect 244642 158760 244648 158772
rect 241848 158732 244648 158760
rect 241848 158720 241854 158732
rect 244642 158720 244648 158732
rect 244700 158720 244706 158772
rect 256878 158720 256884 158772
rect 256936 158760 256942 158772
rect 257982 158760 257988 158772
rect 256936 158732 257988 158760
rect 256936 158720 256942 158732
rect 257982 158720 257988 158732
rect 258040 158720 258046 158772
rect 261110 158720 261116 158772
rect 261168 158760 261174 158772
rect 269022 158760 269028 158772
rect 261168 158732 269028 158760
rect 261168 158720 261174 158732
rect 269022 158720 269028 158732
rect 269080 158720 269086 158772
rect 281258 158720 281264 158772
rect 281316 158760 281322 158772
rect 282546 158760 282552 158772
rect 281316 158732 282552 158760
rect 281316 158720 281322 158732
rect 282546 158720 282552 158732
rect 282604 158720 282610 158772
rect 286318 158720 286324 158772
rect 286376 158760 286382 158772
rect 286870 158760 286876 158772
rect 286376 158732 286876 158760
rect 286376 158720 286382 158732
rect 286870 158720 286876 158732
rect 286928 158720 286934 158772
rect 301498 158720 301504 158772
rect 301556 158760 301562 158772
rect 304810 158760 304816 158772
rect 301556 158732 304816 158760
rect 301556 158720 301562 158732
rect 304810 158720 304816 158732
rect 304868 158720 304874 158772
rect 378870 158720 378876 158772
rect 378928 158760 378934 158772
rect 380986 158760 380992 158772
rect 378928 158732 380992 158760
rect 378928 158720 378934 158732
rect 380986 158720 380992 158732
rect 381044 158720 381050 158772
rect 385586 158720 385592 158772
rect 385644 158760 385650 158772
rect 389082 158760 389088 158772
rect 385644 158732 389088 158760
rect 385644 158720 385650 158732
rect 389082 158720 389088 158732
rect 389140 158720 389146 158772
rect 389818 158720 389824 158772
rect 389876 158760 389882 158772
rect 391566 158760 391572 158772
rect 389876 158732 391572 158760
rect 389876 158720 389882 158732
rect 391566 158720 391572 158732
rect 391624 158720 391630 158772
rect 452838 158720 452844 158772
rect 452896 158760 452902 158772
rect 460106 158760 460112 158772
rect 452896 158732 460112 158760
rect 452896 158720 452902 158732
rect 460106 158720 460112 158732
rect 460164 158720 460170 158772
rect 462130 158720 462136 158772
rect 462188 158760 462194 158772
rect 467834 158760 467840 158772
rect 462188 158732 467840 158760
rect 462188 158720 462194 158732
rect 467834 158720 467840 158732
rect 467892 158720 467898 158772
rect 473078 158720 473084 158772
rect 473136 158760 473142 158772
rect 478966 158760 478972 158772
rect 473136 158732 478972 158760
rect 473136 158720 473142 158732
rect 478966 158720 478972 158732
rect 479024 158720 479030 158772
rect 481450 158720 481456 158772
rect 481508 158760 481514 158772
rect 486418 158760 486424 158772
rect 481508 158732 486424 158760
rect 481508 158720 481514 158732
rect 486418 158720 486424 158732
rect 486476 158720 486482 158772
rect 504450 158720 504456 158772
rect 504508 158760 504514 158772
rect 505002 158760 505008 158772
rect 504508 158732 505008 158760
rect 504508 158720 504514 158732
rect 505002 158720 505008 158732
rect 505060 158720 505066 158772
rect 505830 158720 505836 158772
rect 505888 158760 505894 158772
rect 506750 158760 506756 158772
rect 505888 158732 506756 158760
rect 505888 158720 505894 158732
rect 506750 158720 506756 158732
rect 506808 158720 506814 158772
rect 509694 158720 509700 158772
rect 509752 158760 509758 158772
rect 511718 158760 511724 158772
rect 509752 158732 511724 158760
rect 509752 158720 509758 158732
rect 511718 158720 511724 158732
rect 511776 158720 511782 158772
rect 514846 158720 514852 158772
rect 514904 158760 514910 158772
rect 518526 158760 518532 158772
rect 514904 158732 518532 158760
rect 514904 158720 514910 158732
rect 518526 158720 518532 158732
rect 518584 158720 518590 158772
rect 99558 158652 99564 158704
rect 99616 158692 99622 158704
rect 194962 158692 194968 158704
rect 99616 158664 194968 158692
rect 99616 158652 99622 158664
rect 194962 158652 194968 158664
rect 195020 158652 195026 158704
rect 220170 158652 220176 158704
rect 220228 158692 220234 158704
rect 277946 158692 277952 158704
rect 220228 158664 277952 158692
rect 220228 158652 220234 158664
rect 277946 158652 277952 158664
rect 278004 158652 278010 158704
rect 279602 158652 279608 158704
rect 279660 158692 279666 158704
rect 331306 158692 331312 158704
rect 279660 158664 331312 158692
rect 279660 158652 279666 158664
rect 331306 158652 331312 158664
rect 331364 158652 331370 158704
rect 86126 158584 86132 158636
rect 86184 158624 86190 158636
rect 183554 158624 183560 158636
rect 86184 158596 183560 158624
rect 86184 158584 86190 158596
rect 183554 158584 183560 158596
rect 183612 158584 183618 158636
rect 200574 158584 200580 158636
rect 200632 158624 200638 158636
rect 272058 158624 272064 158636
rect 200632 158596 272064 158624
rect 200632 158584 200638 158596
rect 272058 158584 272064 158596
rect 272116 158584 272122 158636
rect 274542 158584 274548 158636
rect 274600 158624 274606 158636
rect 328546 158624 328552 158636
rect 274600 158596 328552 158624
rect 274600 158584 274606 158596
rect 328546 158584 328552 158596
rect 328604 158584 328610 158636
rect 351914 158584 351920 158636
rect 351972 158624 351978 158636
rect 386506 158624 386512 158636
rect 351972 158596 386512 158624
rect 351972 158584 351978 158596
rect 386506 158584 386512 158596
rect 386564 158584 386570 158636
rect 62574 158516 62580 158568
rect 62632 158556 62638 158568
rect 166718 158556 166724 158568
rect 62632 158528 166724 158556
rect 62632 158516 62638 158528
rect 166718 158516 166724 158528
rect 166776 158516 166782 158568
rect 197170 158516 197176 158568
rect 197228 158556 197234 158568
rect 269390 158556 269396 158568
rect 197228 158528 269396 158556
rect 197228 158516 197234 158528
rect 269390 158516 269396 158528
rect 269448 158516 269454 158568
rect 272886 158516 272892 158568
rect 272944 158556 272950 158568
rect 327074 158556 327080 158568
rect 272944 158528 327080 158556
rect 272944 158516 272950 158528
rect 327074 158516 327080 158528
rect 327132 158516 327138 158568
rect 350258 158516 350264 158568
rect 350316 158556 350322 158568
rect 385218 158556 385224 158568
rect 350316 158528 385224 158556
rect 350316 158516 350322 158528
rect 385218 158516 385224 158528
rect 385276 158516 385282 158568
rect 65978 158448 65984 158500
rect 66036 158488 66042 158500
rect 168374 158488 168380 158500
rect 66036 158460 168380 158488
rect 66036 158448 66042 158460
rect 168374 158448 168380 158460
rect 168432 158448 168438 158500
rect 190454 158448 190460 158500
rect 190512 158488 190518 158500
rect 263778 158488 263784 158500
rect 190512 158460 263784 158488
rect 190512 158448 190518 158460
rect 263778 158448 263784 158460
rect 263836 158448 263842 158500
rect 266170 158448 266176 158500
rect 266228 158488 266234 158500
rect 322106 158488 322112 158500
rect 266228 158460 322112 158488
rect 266228 158448 266234 158460
rect 322106 158448 322112 158460
rect 322164 158448 322170 158500
rect 338482 158448 338488 158500
rect 338540 158488 338546 158500
rect 376846 158488 376852 158500
rect 338540 158460 376852 158488
rect 338540 158448 338546 158460
rect 376846 158448 376852 158460
rect 376904 158448 376910 158500
rect 377214 158448 377220 158500
rect 377272 158488 377278 158500
rect 406838 158488 406844 158500
rect 377272 158460 406844 158488
rect 377272 158448 377278 158460
rect 406838 158448 406844 158460
rect 406896 158448 406902 158500
rect 59262 158380 59268 158432
rect 59320 158420 59326 158432
rect 163038 158420 163044 158432
rect 59320 158392 163044 158420
rect 59320 158380 59326 158392
rect 163038 158380 163044 158392
rect 163096 158380 163102 158432
rect 187050 158380 187056 158432
rect 187108 158420 187114 158432
rect 260834 158420 260840 158432
rect 187108 158392 260840 158420
rect 187108 158380 187114 158392
rect 260834 158380 260840 158392
rect 260892 158380 260898 158432
rect 262766 158380 262772 158432
rect 262824 158420 262830 158432
rect 319530 158420 319536 158432
rect 262824 158392 319536 158420
rect 262824 158380 262830 158392
rect 319530 158380 319536 158392
rect 319588 158380 319594 158432
rect 330110 158380 330116 158432
rect 330168 158420 330174 158432
rect 370866 158420 370872 158432
rect 330168 158392 370872 158420
rect 330168 158380 330174 158392
rect 370866 158380 370872 158392
rect 370924 158380 370930 158432
rect 52454 158312 52460 158364
rect 52512 158352 52518 158364
rect 158990 158352 158996 158364
rect 52512 158324 158996 158352
rect 52512 158312 52518 158324
rect 158990 158312 158996 158324
rect 159048 158312 159054 158364
rect 177022 158312 177028 158364
rect 177080 158352 177086 158364
rect 254026 158352 254032 158364
rect 177080 158324 254032 158352
rect 177080 158312 177086 158324
rect 254026 158312 254032 158324
rect 254084 158312 254090 158364
rect 256050 158312 256056 158364
rect 256108 158352 256114 158364
rect 314378 158352 314384 158364
rect 256108 158324 314384 158352
rect 256108 158312 256114 158324
rect 314378 158312 314384 158324
rect 314436 158312 314442 158364
rect 317414 158312 317420 158364
rect 317472 158352 317478 158364
rect 360194 158352 360200 158364
rect 317472 158324 360200 158352
rect 317472 158312 317478 158324
rect 360194 158312 360200 158324
rect 360252 158312 360258 158364
rect 378042 158312 378048 158364
rect 378100 158352 378106 158364
rect 407390 158352 407396 158364
rect 378100 158324 407396 158352
rect 378100 158312 378106 158324
rect 407390 158312 407396 158324
rect 407448 158312 407454 158364
rect 427354 158352 427360 158364
rect 412606 158324 427360 158352
rect 45738 158244 45744 158296
rect 45796 158284 45802 158296
rect 153378 158284 153384 158296
rect 45796 158256 153384 158284
rect 45796 158244 45802 158256
rect 153378 158244 153384 158256
rect 153436 158244 153442 158296
rect 173618 158244 173624 158296
rect 173676 158284 173682 158296
rect 251450 158284 251456 158296
rect 173676 158256 251456 158284
rect 173676 158244 173682 158256
rect 251450 158244 251456 158256
rect 251508 158244 251514 158296
rect 252646 158244 252652 158296
rect 252704 158284 252710 158296
rect 310606 158284 310612 158296
rect 252704 158256 310612 158284
rect 252704 158244 252710 158256
rect 310606 158244 310612 158256
rect 310664 158244 310670 158296
rect 320818 158244 320824 158296
rect 320876 158284 320882 158296
rect 363506 158284 363512 158296
rect 320876 158256 363512 158284
rect 320876 158244 320882 158256
rect 363506 158244 363512 158256
rect 363564 158244 363570 158296
rect 367094 158244 367100 158296
rect 367152 158284 367158 158296
rect 399110 158284 399116 158296
rect 367152 158256 399116 158284
rect 367152 158244 367158 158256
rect 399110 158244 399116 158256
rect 399168 158244 399174 158296
rect 31478 158176 31484 158228
rect 31536 158216 31542 158228
rect 139486 158216 139492 158228
rect 31536 158188 139492 158216
rect 31536 158176 31542 158188
rect 139486 158176 139492 158188
rect 139544 158176 139550 158228
rect 163498 158176 163504 158228
rect 163556 158216 163562 158228
rect 242894 158216 242900 158228
rect 163556 158188 242900 158216
rect 163556 158176 163562 158188
rect 242894 158176 242900 158188
rect 242952 158176 242958 158228
rect 245930 158176 245936 158228
rect 245988 158216 245994 158228
rect 306374 158216 306380 158228
rect 245988 158188 306380 158216
rect 245988 158176 245994 158188
rect 306374 158176 306380 158188
rect 306432 158176 306438 158228
rect 314102 158176 314108 158228
rect 314160 158216 314166 158228
rect 357618 158216 357624 158228
rect 314160 158188 357624 158216
rect 314160 158176 314166 158188
rect 357618 158176 357624 158188
rect 357676 158176 357682 158228
rect 361206 158176 361212 158228
rect 361264 158216 361270 158228
rect 394694 158216 394700 158228
rect 361264 158188 394700 158216
rect 361264 158176 361270 158188
rect 394694 158176 394700 158188
rect 394752 158176 394758 158228
rect 404078 158176 404084 158228
rect 404136 158216 404142 158228
rect 412606 158216 412634 158324
rect 427354 158312 427360 158324
rect 427412 158312 427418 158364
rect 439406 158244 439412 158296
rect 439464 158284 439470 158296
rect 454402 158284 454408 158296
rect 439464 158256 454408 158284
rect 439464 158244 439470 158256
rect 454402 158244 454408 158256
rect 454460 158244 454466 158296
rect 404136 158188 412634 158216
rect 404136 158176 404142 158188
rect 426434 158176 426440 158228
rect 426492 158216 426498 158228
rect 442994 158216 443000 158228
rect 426492 158188 443000 158216
rect 426492 158176 426498 158188
rect 442994 158176 443000 158188
rect 443052 158176 443058 158228
rect 35710 158108 35716 158160
rect 35768 158148 35774 158160
rect 145098 158148 145104 158160
rect 35768 158120 145104 158148
rect 35768 158108 35774 158120
rect 145098 158108 145104 158120
rect 145156 158108 145162 158160
rect 153470 158108 153476 158160
rect 153528 158148 153534 158160
rect 236086 158148 236092 158160
rect 153528 158120 236092 158148
rect 153528 158108 153534 158120
rect 236086 158108 236092 158120
rect 236144 158108 236150 158160
rect 242618 158108 242624 158160
rect 242676 158148 242682 158160
rect 304074 158148 304080 158160
rect 242676 158120 304080 158148
rect 242676 158108 242682 158120
rect 304074 158108 304080 158120
rect 304132 158108 304138 158160
rect 307386 158108 307392 158160
rect 307444 158148 307450 158160
rect 353294 158148 353300 158160
rect 307444 158120 353300 158148
rect 307444 158108 307450 158120
rect 353294 158108 353300 158120
rect 353352 158108 353358 158160
rect 358630 158108 358636 158160
rect 358688 158148 358694 158160
rect 391934 158148 391940 158160
rect 358688 158120 391940 158148
rect 358688 158108 358694 158120
rect 391934 158108 391940 158120
rect 391992 158108 391998 158160
rect 404906 158108 404912 158160
rect 404964 158148 404970 158160
rect 427998 158148 428004 158160
rect 404964 158120 428004 158148
rect 404964 158108 404970 158120
rect 427998 158108 428004 158120
rect 428056 158108 428062 158160
rect 428458 158108 428464 158160
rect 428516 158148 428522 158160
rect 445754 158148 445760 158160
rect 428516 158120 445760 158148
rect 428516 158108 428522 158120
rect 445754 158108 445760 158120
rect 445812 158108 445818 158160
rect 18874 158040 18880 158092
rect 18932 158080 18938 158092
rect 132494 158080 132500 158092
rect 18932 158052 132500 158080
rect 18932 158040 18938 158052
rect 132494 158040 132500 158052
rect 132552 158040 132558 158092
rect 139946 158040 139952 158092
rect 140004 158080 140010 158092
rect 224954 158080 224960 158092
rect 140004 158052 224960 158080
rect 140004 158040 140010 158052
rect 224954 158040 224960 158052
rect 225012 158040 225018 158092
rect 229094 158040 229100 158092
rect 229152 158080 229158 158092
rect 292758 158080 292764 158092
rect 229152 158052 292764 158080
rect 229152 158040 229158 158052
rect 292758 158040 292764 158052
rect 292816 158040 292822 158092
rect 293034 158040 293040 158092
rect 293092 158080 293098 158092
rect 342254 158080 342260 158092
rect 293092 158052 342260 158080
rect 293092 158040 293098 158052
rect 342254 158040 342260 158052
rect 342312 158040 342318 158092
rect 351086 158040 351092 158092
rect 351144 158080 351150 158092
rect 386966 158080 386972 158092
rect 351144 158052 386972 158080
rect 351144 158040 351150 158052
rect 386966 158040 386972 158052
rect 387024 158040 387030 158092
rect 393958 158040 393964 158092
rect 394016 158080 394022 158092
rect 419534 158080 419540 158092
rect 394016 158052 419540 158080
rect 394016 158040 394022 158052
rect 419534 158040 419540 158052
rect 419592 158040 419598 158092
rect 420914 158040 420920 158092
rect 420972 158080 420978 158092
rect 440326 158080 440332 158092
rect 420972 158052 440332 158080
rect 420972 158040 420978 158052
rect 440326 158040 440332 158052
rect 440384 158040 440390 158092
rect 443638 158040 443644 158092
rect 443696 158080 443702 158092
rect 456794 158080 456800 158092
rect 443696 158052 456800 158080
rect 443696 158040 443702 158052
rect 456794 158040 456800 158052
rect 456852 158040 456858 158092
rect 2130 157972 2136 158024
rect 2188 158012 2194 158024
rect 120074 158012 120080 158024
rect 2188 157984 120080 158012
rect 2188 157972 2194 157984
rect 120074 157972 120080 157984
rect 120132 157972 120138 158024
rect 133230 157972 133236 158024
rect 133288 158012 133294 158024
rect 220630 158012 220636 158024
rect 133288 157984 220636 158012
rect 133288 157972 133294 157984
rect 220630 157972 220636 157984
rect 220688 157972 220694 158024
rect 225690 157972 225696 158024
rect 225748 158012 225754 158024
rect 288434 158012 288440 158024
rect 225748 157984 288440 158012
rect 225748 157972 225754 157984
rect 288434 157972 288440 157984
rect 288492 157972 288498 158024
rect 289722 157972 289728 158024
rect 289780 158012 289786 158024
rect 340046 158012 340052 158024
rect 289780 157984 340052 158012
rect 289780 157972 289786 157984
rect 340046 157972 340052 157984
rect 340104 157972 340110 158024
rect 340138 157972 340144 158024
rect 340196 158012 340202 158024
rect 378594 158012 378600 158024
rect 340196 157984 378600 158012
rect 340196 157972 340202 157984
rect 378594 157972 378600 157984
rect 378652 157972 378658 158024
rect 388070 157972 388076 158024
rect 388128 158012 388134 158024
rect 414566 158012 414572 158024
rect 388128 157984 414572 158012
rect 388128 157972 388134 157984
rect 414566 157972 414572 157984
rect 414624 157972 414630 158024
rect 415026 157972 415032 158024
rect 415084 158012 415090 158024
rect 434714 158012 434720 158024
rect 415084 157984 434720 158012
rect 415084 157972 415090 157984
rect 434714 157972 434720 157984
rect 434772 157972 434778 158024
rect 435174 157972 435180 158024
rect 435232 158012 435238 158024
rect 451182 158012 451188 158024
rect 435232 157984 451188 158012
rect 435232 157972 435238 157984
rect 451182 157972 451188 157984
rect 451240 157972 451246 158024
rect 106366 157904 106372 157956
rect 106424 157944 106430 157956
rect 200114 157944 200120 157956
rect 106424 157916 200120 157944
rect 106424 157904 106430 157916
rect 200114 157904 200120 157916
rect 200172 157904 200178 157956
rect 207014 157904 207020 157956
rect 207072 157944 207078 157956
rect 233234 157944 233240 157956
rect 207072 157916 233240 157944
rect 207072 157904 207078 157916
rect 233234 157904 233240 157916
rect 233292 157904 233298 157956
rect 239214 157904 239220 157956
rect 239272 157944 239278 157956
rect 252002 157944 252008 157956
rect 239272 157916 252008 157944
rect 239272 157904 239278 157916
rect 252002 157904 252008 157916
rect 252060 157904 252066 157956
rect 259454 157904 259460 157956
rect 259512 157944 259518 157956
rect 316954 157944 316960 157956
rect 259512 157916 316960 157944
rect 259512 157904 259518 157916
rect 316954 157904 316960 157916
rect 317012 157904 317018 157956
rect 321646 157904 321652 157956
rect 321704 157944 321710 157956
rect 359458 157944 359464 157956
rect 321704 157916 359464 157944
rect 321704 157904 321710 157916
rect 359458 157904 359464 157916
rect 359516 157904 359522 157956
rect 123110 157836 123116 157888
rect 123168 157876 123174 157888
rect 205634 157876 205640 157888
rect 123168 157848 205640 157876
rect 123168 157836 123174 157848
rect 205634 157836 205640 157848
rect 205692 157836 205698 157888
rect 221550 157836 221556 157888
rect 221608 157876 221614 157888
rect 245654 157876 245660 157888
rect 221608 157848 245660 157876
rect 221608 157836 221614 157848
rect 245654 157836 245660 157848
rect 245712 157836 245718 157888
rect 269482 157836 269488 157888
rect 269540 157876 269546 157888
rect 269540 157848 320496 157876
rect 269540 157836 269546 157848
rect 79410 157768 79416 157820
rect 79468 157808 79474 157820
rect 146110 157808 146116 157820
rect 79468 157780 146116 157808
rect 79468 157768 79474 157780
rect 146110 157768 146116 157780
rect 146168 157768 146174 157820
rect 147674 157768 147680 157820
rect 147732 157808 147738 157820
rect 215386 157808 215392 157820
rect 147732 157780 215392 157808
rect 147732 157768 147738 157780
rect 215386 157768 215392 157780
rect 215444 157768 215450 157820
rect 311894 157768 311900 157820
rect 311952 157808 311958 157820
rect 320468 157808 320496 157848
rect 324314 157836 324320 157888
rect 324372 157876 324378 157888
rect 350534 157876 350540 157888
rect 324372 157848 350540 157876
rect 324372 157836 324378 157848
rect 350534 157836 350540 157848
rect 350592 157836 350598 157888
rect 324682 157808 324688 157820
rect 311952 157780 316034 157808
rect 320468 157780 324688 157808
rect 311952 157768 311958 157780
rect 146018 157700 146024 157752
rect 146076 157740 146082 157752
rect 190454 157740 190460 157752
rect 146076 157712 190460 157740
rect 146076 157700 146082 157712
rect 190454 157700 190460 157712
rect 190512 157700 190518 157752
rect 201310 157700 201316 157752
rect 201368 157740 201374 157752
rect 223850 157740 223856 157752
rect 201368 157712 223856 157740
rect 201368 157700 201374 157712
rect 223850 157700 223856 157712
rect 223908 157700 223914 157752
rect 316006 157672 316034 157780
rect 324682 157768 324688 157780
rect 324740 157768 324746 157820
rect 341334 157808 341340 157820
rect 325666 157780 341340 157808
rect 325666 157672 325694 157780
rect 341334 157768 341340 157780
rect 341392 157768 341398 157820
rect 316006 157644 325694 157672
rect 76006 157292 76012 157344
rect 76064 157332 76070 157344
rect 177022 157332 177028 157344
rect 76064 157304 177028 157332
rect 76064 157292 76070 157304
rect 177022 157292 177028 157304
rect 177080 157292 177086 157344
rect 193766 157292 193772 157344
rect 193824 157332 193830 157344
rect 266906 157332 266912 157344
rect 193824 157304 266912 157332
rect 193824 157292 193830 157304
rect 266906 157292 266912 157304
rect 266964 157292 266970 157344
rect 296438 157292 296444 157344
rect 296496 157332 296502 157344
rect 345014 157332 345020 157344
rect 296496 157304 345020 157332
rect 296496 157292 296502 157304
rect 345014 157292 345020 157304
rect 345072 157292 345078 157344
rect 356146 157292 356152 157344
rect 356204 157332 356210 157344
rect 358814 157332 358820 157344
rect 356204 157304 358820 157332
rect 356204 157292 356210 157304
rect 358814 157292 358820 157304
rect 358872 157292 358878 157344
rect 69290 157224 69296 157276
rect 69348 157264 69354 157276
rect 171134 157264 171140 157276
rect 69348 157236 171140 157264
rect 69348 157224 69354 157236
rect 171134 157224 171140 157236
rect 171192 157224 171198 157276
rect 179506 157224 179512 157276
rect 179564 157264 179570 157276
rect 255866 157264 255872 157276
rect 179564 157236 255872 157264
rect 179564 157224 179570 157236
rect 255866 157224 255872 157236
rect 255924 157224 255930 157276
rect 276198 157224 276204 157276
rect 276256 157264 276262 157276
rect 329834 157264 329840 157276
rect 276256 157236 329840 157264
rect 276256 157224 276262 157236
rect 329834 157224 329840 157236
rect 329892 157224 329898 157276
rect 352006 157224 352012 157276
rect 352064 157264 352070 157276
rect 365898 157264 365904 157276
rect 352064 157236 365904 157264
rect 352064 157224 352070 157236
rect 365898 157224 365904 157236
rect 365956 157224 365962 157276
rect 4522 157156 4528 157208
rect 4580 157196 4586 157208
rect 109126 157196 109132 157208
rect 4580 157168 109132 157196
rect 4580 157156 4586 157168
rect 109126 157156 109132 157168
rect 109184 157156 109190 157208
rect 113082 157156 113088 157208
rect 113140 157196 113146 157208
rect 205266 157196 205272 157208
rect 113140 157168 205272 157196
rect 113140 157156 113146 157168
rect 205266 157156 205272 157168
rect 205324 157156 205330 157208
rect 209774 157156 209780 157208
rect 209832 157196 209838 157208
rect 279050 157196 279056 157208
rect 209832 157168 279056 157196
rect 209832 157156 209838 157168
rect 279050 157156 279056 157168
rect 279108 157156 279114 157208
rect 288618 157156 288624 157208
rect 288676 157196 288682 157208
rect 338666 157196 338672 157208
rect 288676 157168 338672 157196
rect 288676 157156 288682 157168
rect 338666 157156 338672 157168
rect 338724 157156 338730 157208
rect 347774 157156 347780 157208
rect 347832 157196 347838 157208
rect 384390 157196 384396 157208
rect 347832 157168 384396 157196
rect 347832 157156 347838 157168
rect 384390 157156 384396 157168
rect 384448 157156 384454 157208
rect 55858 157088 55864 157140
rect 55916 157128 55922 157140
rect 161566 157128 161572 157140
rect 55916 157100 161572 157128
rect 55916 157088 55922 157100
rect 161566 157088 161572 157100
rect 161624 157088 161630 157140
rect 172790 157088 172796 157140
rect 172848 157128 172854 157140
rect 250806 157128 250812 157140
rect 172848 157100 250812 157128
rect 172848 157088 172854 157100
rect 250806 157088 250812 157100
rect 250864 157088 250870 157140
rect 260282 157088 260288 157140
rect 260340 157128 260346 157140
rect 317414 157128 317420 157140
rect 260340 157100 317420 157128
rect 260340 157088 260346 157100
rect 317414 157088 317420 157100
rect 317472 157088 317478 157140
rect 346854 157088 346860 157140
rect 346912 157128 346918 157140
rect 383746 157128 383752 157140
rect 346912 157100 383752 157128
rect 346912 157088 346918 157100
rect 383746 157088 383752 157100
rect 383804 157088 383810 157140
rect 49142 157020 49148 157072
rect 49200 157060 49206 157072
rect 156414 157060 156420 157072
rect 49200 157032 156420 157060
rect 49200 157020 49206 157032
rect 156414 157020 156420 157032
rect 156472 157020 156478 157072
rect 176102 157020 176108 157072
rect 176160 157060 176166 157072
rect 252554 157060 252560 157072
rect 176160 157032 252560 157060
rect 176160 157020 176166 157032
rect 252554 157020 252560 157032
rect 252612 157020 252618 157072
rect 254394 157020 254400 157072
rect 254452 157060 254458 157072
rect 311894 157060 311900 157072
rect 254452 157032 311900 157060
rect 254452 157020 254458 157032
rect 311894 157020 311900 157032
rect 311952 157020 311958 157072
rect 336826 157020 336832 157072
rect 336884 157060 336890 157072
rect 376018 157060 376024 157072
rect 336884 157032 376024 157060
rect 336884 157020 336890 157032
rect 376018 157020 376024 157032
rect 376076 157020 376082 157072
rect 383102 157020 383108 157072
rect 383160 157060 383166 157072
rect 411346 157060 411352 157072
rect 383160 157032 411352 157060
rect 383160 157020 383166 157032
rect 411346 157020 411352 157032
rect 411404 157020 411410 157072
rect 39022 156952 39028 157004
rect 39080 156992 39086 157004
rect 147674 156992 147680 157004
rect 39080 156964 147680 156992
rect 39080 156952 39086 156964
rect 147674 156952 147680 156964
rect 147732 156952 147738 157004
rect 169386 156952 169392 157004
rect 169444 156992 169450 157004
rect 247126 156992 247132 157004
rect 169444 156964 247132 156992
rect 169444 156952 169450 156964
rect 247126 156952 247132 156964
rect 247184 156952 247190 157004
rect 253566 156952 253572 157004
rect 253624 156992 253630 157004
rect 307018 156992 307024 157004
rect 253624 156964 307024 156992
rect 253624 156952 253630 156964
rect 307018 156952 307024 156964
rect 307076 156952 307082 157004
rect 330938 156952 330944 157004
rect 330996 156992 331002 157004
rect 371234 156992 371240 157004
rect 330996 156964 371240 156992
rect 330996 156952 331002 156964
rect 371234 156952 371240 156964
rect 371292 156952 371298 157004
rect 373810 156952 373816 157004
rect 373868 156992 373874 157004
rect 404078 156992 404084 157004
rect 373868 156964 404084 156992
rect 373868 156952 373874 156964
rect 404078 156952 404084 156964
rect 404136 156952 404142 157004
rect 423398 156952 423404 157004
rect 423456 156992 423462 157004
rect 442166 156992 442172 157004
rect 423456 156964 442172 156992
rect 423456 156952 423462 156964
rect 442166 156952 442172 156964
rect 442224 156952 442230 157004
rect 24762 156884 24768 156936
rect 24820 156924 24826 156936
rect 137830 156924 137836 156936
rect 24820 156896 137836 156924
rect 24820 156884 24826 156896
rect 137830 156884 137836 156896
rect 137888 156884 137894 156936
rect 160186 156884 160192 156936
rect 160244 156924 160250 156936
rect 241238 156924 241244 156936
rect 160244 156896 241244 156924
rect 160244 156884 160250 156896
rect 241238 156884 241244 156896
rect 241296 156884 241302 156936
rect 249334 156884 249340 156936
rect 249392 156924 249398 156936
rect 306374 156924 306380 156936
rect 249392 156896 306380 156924
rect 249392 156884 249398 156896
rect 306374 156884 306380 156896
rect 306432 156884 306438 156936
rect 307294 156924 307300 156936
rect 306484 156896 307300 156924
rect 21358 156816 21364 156868
rect 21416 156856 21422 156868
rect 135254 156856 135260 156868
rect 21416 156828 135260 156856
rect 21416 156816 21422 156828
rect 135254 156816 135260 156828
rect 135312 156816 135318 156868
rect 150066 156816 150072 156868
rect 150124 156856 150130 156868
rect 233510 156856 233516 156868
rect 150124 156828 233516 156856
rect 150124 156816 150130 156828
rect 233510 156816 233516 156828
rect 233568 156816 233574 156868
rect 246758 156816 246764 156868
rect 246816 156856 246822 156868
rect 306484 156856 306512 156896
rect 307294 156884 307300 156896
rect 307352 156884 307358 156936
rect 310698 156884 310704 156936
rect 310756 156924 310762 156936
rect 356146 156924 356152 156936
rect 310756 156896 356152 156924
rect 310756 156884 310762 156896
rect 356146 156884 356152 156896
rect 356204 156884 356210 156936
rect 374638 156884 374644 156936
rect 374696 156924 374702 156936
rect 404446 156924 404452 156936
rect 374696 156896 404452 156924
rect 374696 156884 374702 156896
rect 404446 156884 404452 156896
rect 404504 156884 404510 156936
rect 411622 156884 411628 156936
rect 411680 156924 411686 156936
rect 433150 156924 433156 156936
rect 411680 156896 433156 156924
rect 411680 156884 411686 156896
rect 433150 156884 433156 156896
rect 433208 156884 433214 156936
rect 246816 156828 306512 156856
rect 246816 156816 246822 156828
rect 306650 156816 306656 156868
rect 306708 156856 306714 156868
rect 351914 156856 351920 156868
rect 306708 156828 351920 156856
rect 306708 156816 306714 156828
rect 351914 156816 351920 156828
rect 351972 156816 351978 156868
rect 363690 156816 363696 156868
rect 363748 156856 363754 156868
rect 396534 156856 396540 156868
rect 363748 156828 396540 156856
rect 363748 156816 363754 156828
rect 396534 156816 396540 156828
rect 396592 156816 396598 156868
rect 401594 156816 401600 156868
rect 401652 156856 401658 156868
rect 425146 156856 425152 156868
rect 401652 156828 425152 156856
rect 401652 156816 401658 156828
rect 425146 156816 425152 156828
rect 425204 156816 425210 156868
rect 433058 156816 433064 156868
rect 433116 156856 433122 156868
rect 447318 156856 447324 156868
rect 433116 156828 447324 156856
rect 433116 156816 433122 156828
rect 447318 156816 447324 156828
rect 447376 156816 447382 156868
rect 18046 156748 18052 156800
rect 18104 156788 18110 156800
rect 132678 156788 132684 156800
rect 18104 156760 132684 156788
rect 18104 156748 18110 156760
rect 132678 156748 132684 156760
rect 132736 156748 132742 156800
rect 136634 156748 136640 156800
rect 136692 156788 136698 156800
rect 222746 156788 222752 156800
rect 136692 156760 222752 156788
rect 136692 156748 136698 156760
rect 222746 156748 222752 156760
rect 222804 156748 222810 156800
rect 236730 156748 236736 156800
rect 236788 156788 236794 156800
rect 299474 156788 299480 156800
rect 236788 156760 299480 156788
rect 236788 156748 236794 156760
rect 299474 156748 299480 156760
rect 299532 156748 299538 156800
rect 299750 156748 299756 156800
rect 299808 156788 299814 156800
rect 347774 156788 347780 156800
rect 299808 156760 347780 156788
rect 299808 156748 299814 156760
rect 347774 156748 347780 156760
rect 347832 156748 347838 156800
rect 348602 156748 348608 156800
rect 348660 156788 348666 156800
rect 385034 156788 385040 156800
rect 348660 156760 385040 156788
rect 348660 156748 348666 156760
rect 385034 156748 385040 156760
rect 385092 156748 385098 156800
rect 387242 156748 387248 156800
rect 387300 156788 387306 156800
rect 414106 156788 414112 156800
rect 387300 156760 414112 156788
rect 387300 156748 387306 156760
rect 414106 156748 414112 156760
rect 414164 156748 414170 156800
rect 414198 156748 414204 156800
rect 414256 156788 414262 156800
rect 435082 156788 435088 156800
rect 414256 156760 435088 156788
rect 414256 156748 414262 156760
rect 435082 156748 435088 156760
rect 435140 156748 435146 156800
rect 436370 156748 436376 156800
rect 436428 156788 436434 156800
rect 448606 156788 448612 156800
rect 436428 156760 448612 156788
rect 436428 156748 436434 156760
rect 448606 156748 448612 156760
rect 448664 156748 448670 156800
rect 11238 156680 11244 156732
rect 11296 156720 11302 156732
rect 125686 156720 125692 156732
rect 11296 156692 125692 156720
rect 11296 156680 11302 156692
rect 125686 156680 125692 156692
rect 125744 156680 125750 156732
rect 126514 156680 126520 156732
rect 126572 156720 126578 156732
rect 215478 156720 215484 156732
rect 126572 156692 215484 156720
rect 126572 156680 126578 156692
rect 215478 156680 215484 156692
rect 215536 156680 215542 156732
rect 216674 156680 216680 156732
rect 216732 156720 216738 156732
rect 282086 156720 282092 156732
rect 216732 156692 282092 156720
rect 216732 156680 216738 156692
rect 282086 156680 282092 156692
rect 282144 156680 282150 156732
rect 283006 156680 283012 156732
rect 283064 156720 283070 156732
rect 334894 156720 334900 156732
rect 283064 156692 334900 156720
rect 283064 156680 283070 156692
rect 334894 156680 334900 156692
rect 334952 156680 334958 156732
rect 341886 156680 341892 156732
rect 341944 156720 341950 156732
rect 379882 156720 379888 156732
rect 341944 156692 379888 156720
rect 341944 156680 341950 156692
rect 379882 156680 379888 156692
rect 379940 156680 379946 156732
rect 384758 156680 384764 156732
rect 384816 156720 384822 156732
rect 412634 156720 412640 156732
rect 384816 156692 412640 156720
rect 384816 156680 384822 156692
rect 412634 156680 412640 156692
rect 412692 156680 412698 156732
rect 419258 156680 419264 156732
rect 419316 156720 419322 156732
rect 438946 156720 438952 156732
rect 419316 156692 438952 156720
rect 419316 156680 419322 156692
rect 438946 156680 438952 156692
rect 439004 156680 439010 156732
rect 14642 156612 14648 156664
rect 14700 156652 14706 156664
rect 129734 156652 129740 156664
rect 14700 156624 129740 156652
rect 14700 156612 14706 156624
rect 129734 156612 129740 156624
rect 129792 156612 129798 156664
rect 129918 156612 129924 156664
rect 129976 156652 129982 156664
rect 218054 156652 218060 156664
rect 129976 156624 218060 156652
rect 129976 156612 129982 156624
rect 218054 156612 218060 156624
rect 218112 156612 218118 156664
rect 240042 156612 240048 156664
rect 240100 156652 240106 156664
rect 302234 156652 302240 156664
rect 240100 156624 302240 156652
rect 240100 156612 240106 156624
rect 302234 156612 302240 156624
rect 302292 156612 302298 156664
rect 303982 156612 303988 156664
rect 304040 156652 304046 156664
rect 350994 156652 351000 156664
rect 304040 156624 351000 156652
rect 304040 156612 304046 156624
rect 350994 156612 351000 156624
rect 351052 156612 351058 156664
rect 357802 156612 357808 156664
rect 357860 156652 357866 156664
rect 392118 156652 392124 156664
rect 357860 156624 392124 156652
rect 357860 156612 357866 156624
rect 392118 156612 392124 156624
rect 392176 156612 392182 156664
rect 400766 156612 400772 156664
rect 400824 156652 400830 156664
rect 423766 156652 423772 156664
rect 400824 156624 423772 156652
rect 400824 156612 400830 156624
rect 423766 156612 423772 156624
rect 423824 156612 423830 156664
rect 427630 156612 427636 156664
rect 427688 156652 427694 156664
rect 444374 156652 444380 156664
rect 427688 156624 444380 156652
rect 427688 156612 427694 156624
rect 444374 156612 444380 156624
rect 444432 156612 444438 156664
rect 445294 156612 445300 156664
rect 445352 156652 445358 156664
rect 458818 156652 458824 156664
rect 445352 156624 458824 156652
rect 445352 156612 445358 156624
rect 458818 156612 458824 156624
rect 458876 156612 458882 156664
rect 96246 156544 96252 156596
rect 96304 156584 96310 156596
rect 192386 156584 192392 156596
rect 96304 156556 192392 156584
rect 96304 156544 96310 156556
rect 192386 156544 192392 156556
rect 192444 156544 192450 156596
rect 215018 156544 215024 156596
rect 215076 156584 215082 156596
rect 278774 156584 278780 156596
rect 215076 156556 278780 156584
rect 215076 156544 215082 156556
rect 278774 156544 278780 156556
rect 278832 156544 278838 156596
rect 303154 156544 303160 156596
rect 303212 156584 303218 156596
rect 349246 156584 349252 156596
rect 303212 156556 349252 156584
rect 303212 156544 303218 156556
rect 349246 156544 349252 156556
rect 349304 156544 349310 156596
rect 116394 156476 116400 156528
rect 116452 156516 116458 156528
rect 207014 156516 207020 156528
rect 116452 156488 207020 156516
rect 116452 156476 116458 156488
rect 207014 156476 207020 156488
rect 207072 156476 207078 156528
rect 227714 156476 227720 156528
rect 227772 156516 227778 156528
rect 289998 156516 290004 156528
rect 227772 156488 290004 156516
rect 227772 156476 227778 156488
rect 289998 156476 290004 156488
rect 290056 156476 290062 156528
rect 307018 156476 307024 156528
rect 307076 156516 307082 156528
rect 312446 156516 312452 156528
rect 307076 156488 312452 156516
rect 307076 156476 307082 156488
rect 312446 156476 312452 156488
rect 312504 156476 312510 156528
rect 317782 156476 317788 156528
rect 317840 156516 317846 156528
rect 354214 156516 354220 156528
rect 317840 156488 354220 156516
rect 317840 156476 317846 156488
rect 354214 156476 354220 156488
rect 354272 156476 354278 156528
rect 135622 156408 135628 156460
rect 135680 156448 135686 156460
rect 169938 156448 169944 156460
rect 135680 156420 169944 156448
rect 135680 156408 135686 156420
rect 169938 156408 169944 156420
rect 169996 156408 170002 156460
rect 176654 156408 176660 156460
rect 176712 156448 176718 156460
rect 248874 156448 248880 156460
rect 176712 156420 248880 156448
rect 176712 156408 176718 156420
rect 248874 156408 248880 156420
rect 248932 156408 248938 156460
rect 251726 156408 251732 156460
rect 251784 156448 251790 156460
rect 300302 156448 300308 156460
rect 251784 156420 300308 156448
rect 251784 156408 251790 156420
rect 300302 156408 300308 156420
rect 300360 156408 300366 156460
rect 306374 156408 306380 156460
rect 306432 156448 306438 156460
rect 309226 156448 309232 156460
rect 306432 156420 309232 156448
rect 306432 156408 306438 156420
rect 309226 156408 309232 156420
rect 309284 156408 309290 156460
rect 311986 156408 311992 156460
rect 312044 156448 312050 156460
rect 346486 156448 346492 156460
rect 312044 156420 346492 156448
rect 312044 156408 312050 156420
rect 346486 156408 346492 156420
rect 346544 156408 346550 156460
rect 133506 156340 133512 156392
rect 133564 156380 133570 156392
rect 164418 156380 164424 156392
rect 133564 156352 164424 156380
rect 133564 156340 133570 156352
rect 164418 156340 164424 156352
rect 164476 156340 164482 156392
rect 279510 156340 279516 156392
rect 279568 156380 279574 156392
rect 323394 156380 323400 156392
rect 279568 156352 323400 156380
rect 279568 156340 279574 156352
rect 323394 156340 323400 156352
rect 323452 156340 323458 156392
rect 72694 155864 72700 155916
rect 72752 155904 72758 155916
rect 174446 155904 174452 155916
rect 72752 155876 174452 155904
rect 72752 155864 72758 155876
rect 174446 155864 174452 155876
rect 174504 155864 174510 155916
rect 203886 155864 203892 155916
rect 203944 155904 203950 155916
rect 273438 155904 273444 155916
rect 203944 155876 273444 155904
rect 203944 155864 203950 155876
rect 273438 155864 273444 155876
rect 273496 155864 273502 155916
rect 324222 155864 324228 155916
rect 324280 155904 324286 155916
rect 366266 155904 366272 155916
rect 324280 155876 366272 155904
rect 324280 155864 324286 155876
rect 366266 155864 366272 155876
rect 366324 155864 366330 155916
rect 378134 155864 378140 155916
rect 378192 155904 378198 155916
rect 382274 155904 382280 155916
rect 378192 155876 382280 155904
rect 378192 155864 378198 155876
rect 382274 155864 382280 155876
rect 382332 155864 382338 155916
rect 55030 155796 55036 155848
rect 55088 155836 55094 155848
rect 160094 155836 160100 155848
rect 55088 155808 160100 155836
rect 55088 155796 55094 155808
rect 160094 155796 160100 155808
rect 160152 155796 160158 155848
rect 206462 155796 206468 155848
rect 206520 155836 206526 155848
rect 276474 155836 276480 155848
rect 206520 155808 276480 155836
rect 206520 155796 206526 155808
rect 276474 155796 276480 155808
rect 276532 155796 276538 155848
rect 287146 155796 287152 155848
rect 287204 155836 287210 155848
rect 338114 155836 338120 155848
rect 287204 155808 338120 155836
rect 287204 155796 287210 155808
rect 338114 155796 338120 155808
rect 338172 155796 338178 155848
rect 346302 155796 346308 155848
rect 346360 155836 346366 155848
rect 352282 155836 352288 155848
rect 346360 155808 352288 155836
rect 346360 155796 346366 155808
rect 352282 155796 352288 155808
rect 352340 155796 352346 155848
rect 48314 155728 48320 155780
rect 48372 155768 48378 155780
rect 154666 155768 154672 155780
rect 48372 155740 154672 155768
rect 48372 155728 48378 155740
rect 154666 155728 154672 155740
rect 154724 155728 154730 155780
rect 199654 155728 199660 155780
rect 199712 155768 199718 155780
rect 271046 155768 271052 155780
rect 199712 155740 271052 155768
rect 199712 155728 199718 155740
rect 271046 155728 271052 155740
rect 271104 155728 271110 155780
rect 280430 155728 280436 155780
rect 280488 155768 280494 155780
rect 333054 155768 333060 155780
rect 280488 155740 333060 155768
rect 280488 155728 280494 155740
rect 333054 155728 333060 155740
rect 333112 155728 333118 155780
rect 336642 155728 336648 155780
rect 336700 155768 336706 155780
rect 361942 155768 361948 155780
rect 336700 155740 361948 155768
rect 336700 155728 336706 155740
rect 361942 155728 361948 155740
rect 362000 155728 362006 155780
rect 362126 155728 362132 155780
rect 362184 155768 362190 155780
rect 367646 155768 367652 155780
rect 362184 155740 367652 155768
rect 362184 155728 362190 155740
rect 367646 155728 367652 155740
rect 367704 155728 367710 155780
rect 370406 155728 370412 155780
rect 370464 155768 370470 155780
rect 401686 155768 401692 155780
rect 370464 155740 401692 155768
rect 370464 155728 370470 155740
rect 401686 155728 401692 155740
rect 401744 155728 401750 155780
rect 41598 155660 41604 155712
rect 41656 155700 41662 155712
rect 150618 155700 150624 155712
rect 41656 155672 150624 155700
rect 41656 155660 41662 155672
rect 150618 155660 150624 155672
rect 150676 155660 150682 155712
rect 192938 155660 192944 155712
rect 192996 155700 193002 155712
rect 265158 155700 265164 155712
rect 192996 155672 265164 155700
rect 192996 155660 193002 155672
rect 265158 155660 265164 155672
rect 265216 155660 265222 155712
rect 277118 155660 277124 155712
rect 277176 155700 277182 155712
rect 330018 155700 330024 155712
rect 277176 155672 330024 155700
rect 277176 155660 277182 155672
rect 330018 155660 330024 155672
rect 330076 155660 330082 155712
rect 334250 155660 334256 155712
rect 334308 155700 334314 155712
rect 374086 155700 374092 155712
rect 334308 155672 374092 155700
rect 334308 155660 334314 155672
rect 374086 155660 374092 155672
rect 374144 155660 374150 155712
rect 23934 155592 23940 155644
rect 23992 155632 23998 155644
rect 136726 155632 136732 155644
rect 23992 155604 136732 155632
rect 23992 155592 23998 155604
rect 136726 155592 136732 155604
rect 136784 155592 136790 155644
rect 160278 155592 160284 155644
rect 160336 155632 160342 155644
rect 185026 155632 185032 155644
rect 160336 155604 185032 155632
rect 160336 155592 160342 155604
rect 185026 155592 185032 155604
rect 185084 155592 185090 155644
rect 186222 155592 186228 155644
rect 186280 155632 186286 155644
rect 261110 155632 261116 155644
rect 186280 155604 261116 155632
rect 186280 155592 186286 155604
rect 261110 155592 261116 155604
rect 261168 155592 261174 155644
rect 273714 155592 273720 155644
rect 273772 155632 273778 155644
rect 327902 155632 327908 155644
rect 273772 155604 327908 155632
rect 273772 155592 273778 155604
rect 327902 155592 327908 155604
rect 327960 155592 327966 155644
rect 328362 155592 328368 155644
rect 328420 155632 328426 155644
rect 368934 155632 368940 155644
rect 328420 155604 368940 155632
rect 328420 155592 328426 155604
rect 368934 155592 368940 155604
rect 368992 155592 368998 155644
rect 369578 155592 369584 155644
rect 369636 155632 369642 155644
rect 400214 155632 400220 155644
rect 369636 155604 400220 155632
rect 369636 155592 369642 155604
rect 400214 155592 400220 155604
rect 400272 155592 400278 155644
rect 22186 155524 22192 155576
rect 22244 155564 22250 155576
rect 135806 155564 135812 155576
rect 22244 155536 135812 155564
rect 22244 155524 22250 155536
rect 135806 155524 135812 155536
rect 135864 155524 135870 155576
rect 150434 155524 150440 155576
rect 150492 155564 150498 155576
rect 229186 155564 229192 155576
rect 150492 155536 229192 155564
rect 150492 155524 150498 155536
rect 229186 155524 229192 155536
rect 229244 155524 229250 155576
rect 230014 155524 230020 155576
rect 230072 155564 230078 155576
rect 294506 155564 294512 155576
rect 230072 155536 294512 155564
rect 230072 155524 230078 155536
rect 294506 155524 294512 155536
rect 294564 155524 294570 155576
rect 297266 155524 297272 155576
rect 297324 155564 297330 155576
rect 345842 155564 345848 155576
rect 297324 155536 345848 155564
rect 297324 155524 297330 155536
rect 345842 155524 345848 155536
rect 345900 155524 345906 155576
rect 364518 155524 364524 155576
rect 364576 155564 364582 155576
rect 396166 155564 396172 155576
rect 364576 155536 396172 155564
rect 364576 155524 364582 155536
rect 396166 155524 396172 155536
rect 396224 155524 396230 155576
rect 15470 155456 15476 155508
rect 15528 155496 15534 155508
rect 130286 155496 130292 155508
rect 15528 155468 130292 155496
rect 15528 155456 15534 155468
rect 130286 155456 130292 155468
rect 130344 155456 130350 155508
rect 156782 155456 156788 155508
rect 156840 155496 156846 155508
rect 238570 155496 238576 155508
rect 156840 155468 238576 155496
rect 156840 155456 156846 155468
rect 238570 155456 238576 155468
rect 238628 155456 238634 155508
rect 238662 155456 238668 155508
rect 238720 155496 238726 155508
rect 294046 155496 294052 155508
rect 238720 155468 294052 155496
rect 238720 155456 238726 155468
rect 294046 155456 294052 155468
rect 294104 155456 294110 155508
rect 294782 155456 294788 155508
rect 294840 155496 294846 155508
rect 343910 155496 343916 155508
rect 294840 155468 343916 155496
rect 294840 155456 294846 155468
rect 343910 155456 343916 155468
rect 343968 155456 343974 155508
rect 353662 155456 353668 155508
rect 353720 155496 353726 155508
rect 388346 155496 388352 155508
rect 353720 155468 388352 155496
rect 353720 155456 353726 155468
rect 388346 155456 388352 155468
rect 388404 155456 388410 155508
rect 408310 155456 408316 155508
rect 408368 155496 408374 155508
rect 430574 155496 430580 155508
rect 408368 155468 430580 155496
rect 408368 155456 408374 155468
rect 430574 155456 430580 155468
rect 430632 155456 430638 155508
rect 433242 155456 433248 155508
rect 433300 155496 433306 155508
rect 444742 155496 444748 155508
rect 433300 155468 444748 155496
rect 433300 155456 433306 155468
rect 444742 155456 444748 155468
rect 444800 155456 444806 155508
rect 8754 155388 8760 155440
rect 8812 155428 8818 155440
rect 125594 155428 125600 155440
rect 8812 155400 125600 155428
rect 8812 155388 8818 155400
rect 125594 155388 125600 155400
rect 125652 155388 125658 155440
rect 138290 155388 138296 155440
rect 138348 155428 138354 155440
rect 222010 155428 222016 155440
rect 138348 155400 222016 155428
rect 138348 155388 138354 155400
rect 222010 155388 222016 155400
rect 222068 155388 222074 155440
rect 225782 155388 225788 155440
rect 225840 155428 225846 155440
rect 291286 155428 291292 155440
rect 225840 155400 291292 155428
rect 225840 155388 225846 155400
rect 291286 155388 291292 155400
rect 291344 155388 291350 155440
rect 293862 155388 293868 155440
rect 293920 155428 293926 155440
rect 343266 155428 343272 155440
rect 293920 155400 343272 155428
rect 293920 155388 293926 155400
rect 343266 155388 343272 155400
rect 343324 155388 343330 155440
rect 344370 155388 344376 155440
rect 344428 155428 344434 155440
rect 380894 155428 380900 155440
rect 344428 155400 380900 155428
rect 344428 155388 344434 155400
rect 380894 155388 380900 155400
rect 380952 155388 380958 155440
rect 394878 155388 394884 155440
rect 394936 155428 394942 155440
rect 420362 155428 420368 155440
rect 394936 155400 420368 155428
rect 394936 155388 394942 155400
rect 420362 155388 420368 155400
rect 420420 155388 420426 155440
rect 429286 155388 429292 155440
rect 429344 155428 429350 155440
rect 446674 155428 446680 155440
rect 429344 155400 446680 155428
rect 429344 155388 429350 155400
rect 446674 155388 446680 155400
rect 446732 155388 446738 155440
rect 2866 155320 2872 155372
rect 2924 155360 2930 155372
rect 121086 155360 121092 155372
rect 2924 155332 121092 155360
rect 2924 155320 2930 155332
rect 121086 155320 121092 155332
rect 121144 155320 121150 155372
rect 146662 155320 146668 155372
rect 146720 155360 146726 155372
rect 230934 155360 230940 155372
rect 146720 155332 230940 155360
rect 146720 155320 146726 155332
rect 230934 155320 230940 155332
rect 230992 155320 230998 155372
rect 232498 155320 232504 155372
rect 232556 155360 232562 155372
rect 296438 155360 296444 155372
rect 232556 155332 296444 155360
rect 232556 155320 232562 155332
rect 296438 155320 296444 155332
rect 296496 155320 296502 155372
rect 300670 155320 300676 155372
rect 300728 155360 300734 155372
rect 348418 155360 348424 155372
rect 300728 155332 348424 155360
rect 300728 155320 300734 155332
rect 348418 155320 348424 155332
rect 348476 155320 348482 155372
rect 354490 155320 354496 155372
rect 354548 155360 354554 155372
rect 389542 155360 389548 155372
rect 354548 155332 389548 155360
rect 354548 155320 354554 155332
rect 389542 155320 389548 155332
rect 389600 155320 389606 155372
rect 397362 155320 397368 155372
rect 397420 155360 397426 155372
rect 422294 155360 422300 155372
rect 397420 155332 422300 155360
rect 397420 155320 397426 155332
rect 422294 155320 422300 155332
rect 422352 155320 422358 155372
rect 424318 155320 424324 155372
rect 424376 155360 424382 155372
rect 441706 155360 441712 155372
rect 424376 155332 441712 155360
rect 424376 155320 424382 155332
rect 441706 155320 441712 155332
rect 441764 155320 441770 155372
rect 444466 155320 444472 155372
rect 444524 155360 444530 155372
rect 458174 155360 458180 155372
rect 444524 155332 458180 155360
rect 444524 155320 444530 155332
rect 458174 155320 458180 155332
rect 458232 155320 458238 155372
rect 5350 155252 5356 155304
rect 5408 155292 5414 155304
rect 123018 155292 123024 155304
rect 5408 155264 123024 155292
rect 5408 155252 5414 155264
rect 123018 155252 123024 155264
rect 123076 155252 123082 155304
rect 136082 155252 136088 155304
rect 136140 155292 136146 155304
rect 219526 155292 219532 155304
rect 136140 155264 219532 155292
rect 136140 155252 136146 155264
rect 219526 155252 219532 155264
rect 219584 155252 219590 155304
rect 223206 155252 223212 155304
rect 223264 155292 223270 155304
rect 289354 155292 289360 155304
rect 223264 155264 289360 155292
rect 223264 155252 223270 155264
rect 289354 155252 289360 155264
rect 289412 155252 289418 155304
rect 290550 155252 290556 155304
rect 290608 155292 290614 155304
rect 339586 155292 339592 155304
rect 290608 155264 339592 155292
rect 290608 155252 290614 155264
rect 339586 155252 339592 155264
rect 339644 155252 339650 155304
rect 345198 155252 345204 155304
rect 345256 155292 345262 155304
rect 382458 155292 382464 155304
rect 345256 155264 382464 155292
rect 345256 155252 345262 155264
rect 382458 155252 382464 155264
rect 382516 155252 382522 155304
rect 383930 155252 383936 155304
rect 383988 155292 383994 155304
rect 411990 155292 411996 155304
rect 383988 155264 411996 155292
rect 383988 155252 383994 155264
rect 411990 155252 411996 155264
rect 412048 155252 412054 155304
rect 421742 155252 421748 155304
rect 421800 155292 421806 155304
rect 440878 155292 440884 155304
rect 421800 155264 440884 155292
rect 421800 155252 421806 155264
rect 440878 155252 440884 155264
rect 440936 155252 440942 155304
rect 441982 155252 441988 155304
rect 442040 155292 442046 155304
rect 455966 155292 455972 155304
rect 442040 155264 455972 155292
rect 442040 155252 442046 155264
rect 455966 155252 455972 155264
rect 456024 155252 456030 155304
rect 1210 155184 1216 155236
rect 1268 155224 1274 155236
rect 118786 155224 118792 155236
rect 1268 155196 118792 155224
rect 1268 155184 1274 155196
rect 118786 155184 118792 155196
rect 118844 155184 118850 155236
rect 125778 155184 125784 155236
rect 125836 155224 125842 155236
rect 214834 155224 214840 155236
rect 125836 155196 214840 155224
rect 125836 155184 125842 155196
rect 214834 155184 214840 155196
rect 214892 155184 214898 155236
rect 216490 155184 216496 155236
rect 216548 155224 216554 155236
rect 283098 155224 283104 155236
rect 216548 155196 283104 155224
rect 216548 155184 216554 155196
rect 283098 155184 283104 155196
rect 283156 155184 283162 155236
rect 283834 155184 283840 155236
rect 283892 155224 283898 155236
rect 335538 155224 335544 155236
rect 283892 155196 335544 155224
rect 283892 155184 283898 155196
rect 335538 155184 335544 155196
rect 335596 155184 335602 155236
rect 343542 155184 343548 155236
rect 343600 155224 343606 155236
rect 381170 155224 381176 155236
rect 343600 155196 381176 155224
rect 343600 155184 343606 155196
rect 381170 155184 381176 155196
rect 381228 155184 381234 155236
rect 381354 155184 381360 155236
rect 381412 155224 381418 155236
rect 410058 155224 410064 155236
rect 381412 155196 410064 155224
rect 381412 155184 381418 155196
rect 410058 155184 410064 155196
rect 410116 155184 410122 155236
rect 410794 155184 410800 155236
rect 410852 155224 410858 155236
rect 432046 155224 432052 155236
rect 410852 155196 432052 155224
rect 410852 155184 410858 155196
rect 432046 155184 432052 155196
rect 432104 155184 432110 155236
rect 442810 155184 442816 155236
rect 442868 155224 442874 155236
rect 456978 155224 456984 155236
rect 442868 155196 456984 155224
rect 442868 155184 442874 155196
rect 456978 155184 456984 155196
rect 457036 155184 457042 155236
rect 89530 155116 89536 155168
rect 89588 155156 89594 155168
rect 187234 155156 187240 155168
rect 89588 155128 187240 155156
rect 89588 155116 89594 155128
rect 187234 155116 187240 155128
rect 187292 155116 187298 155168
rect 219066 155116 219072 155168
rect 219124 155156 219130 155168
rect 286134 155156 286140 155168
rect 219124 155128 286140 155156
rect 219124 155116 219130 155128
rect 286134 155116 286140 155128
rect 286192 155116 286198 155168
rect 291470 155116 291476 155168
rect 291528 155156 291534 155168
rect 331122 155156 331128 155168
rect 291528 155128 331128 155156
rect 291528 155116 291534 155128
rect 331122 155116 331128 155128
rect 331180 155116 331186 155168
rect 356790 155156 356796 155168
rect 335326 155128 356796 155156
rect 118694 155048 118700 155100
rect 118752 155088 118758 155100
rect 201586 155088 201592 155100
rect 118752 155060 201592 155088
rect 118752 155048 118758 155060
rect 201586 155048 201592 155060
rect 201644 155048 201650 155100
rect 226610 155048 226616 155100
rect 226668 155088 226674 155100
rect 291194 155088 291200 155100
rect 226668 155060 291200 155088
rect 226668 155048 226674 155060
rect 291194 155048 291200 155060
rect 291252 155048 291258 155100
rect 330202 155048 330208 155100
rect 330260 155088 330266 155100
rect 335326 155088 335354 155128
rect 356790 155116 356796 155128
rect 356848 155116 356854 155168
rect 330260 155060 335354 155088
rect 330260 155048 330266 155060
rect 128170 154980 128176 155032
rect 128228 155020 128234 155032
rect 197446 155020 197452 155032
rect 128228 154992 197452 155020
rect 128228 154980 128234 154992
rect 197446 154980 197452 154992
rect 197504 154980 197510 155032
rect 269022 154980 269028 155032
rect 269080 155020 269086 155032
rect 317966 155020 317972 155032
rect 269080 154992 317972 155020
rect 269080 154980 269086 154992
rect 317966 154980 317972 154992
rect 318024 154980 318030 155032
rect 120166 154912 120172 154964
rect 120224 154952 120230 154964
rect 154206 154952 154212 154964
rect 120224 154924 154212 154952
rect 120224 154912 120230 154924
rect 154206 154912 154212 154924
rect 154264 154912 154270 154964
rect 157334 154912 157340 154964
rect 157392 154952 157398 154964
rect 225138 154952 225144 154964
rect 157392 154924 225144 154952
rect 157392 154912 157398 154924
rect 225138 154912 225144 154924
rect 225196 154912 225202 154964
rect 262122 154912 262128 154964
rect 262180 154952 262186 154964
rect 307938 154952 307944 154964
rect 262180 154924 307944 154952
rect 262180 154912 262186 154924
rect 307938 154912 307944 154924
rect 307996 154912 308002 154964
rect 134886 154844 134892 154896
rect 134944 154884 134950 154896
rect 197354 154884 197360 154896
rect 134944 154856 197360 154884
rect 134944 154844 134950 154856
rect 197354 154844 197360 154856
rect 197412 154844 197418 154896
rect 118142 154776 118148 154828
rect 118200 154816 118206 154828
rect 144822 154816 144828 154828
rect 118200 154788 144828 154816
rect 118200 154776 118206 154788
rect 144822 154776 144828 154788
rect 144880 154776 144886 154828
rect 183278 154776 183284 154828
rect 183336 154816 183342 154828
rect 209958 154816 209964 154828
rect 183336 154788 209964 154816
rect 183336 154776 183342 154788
rect 209958 154776 209964 154788
rect 210016 154776 210022 154828
rect 103422 154504 103428 154556
rect 103480 154544 103486 154556
rect 197538 154544 197544 154556
rect 103480 154516 197544 154544
rect 103480 154504 103486 154516
rect 197538 154504 197544 154516
rect 197596 154504 197602 154556
rect 215662 154504 215668 154556
rect 215720 154544 215726 154556
rect 283558 154544 283564 154556
rect 215720 154516 283564 154544
rect 215720 154504 215726 154516
rect 283558 154504 283564 154516
rect 283616 154504 283622 154556
rect 284294 154504 284300 154556
rect 284352 154544 284358 154556
rect 320910 154544 320916 154556
rect 284352 154516 320916 154544
rect 284352 154504 284358 154516
rect 320910 154504 320916 154516
rect 320968 154504 320974 154556
rect 338758 154504 338764 154556
rect 338816 154544 338822 154556
rect 341978 154544 341984 154556
rect 338816 154516 341984 154544
rect 338816 154504 338822 154516
rect 341978 154504 341984 154516
rect 342036 154504 342042 154556
rect 92842 154436 92848 154488
rect 92900 154476 92906 154488
rect 189810 154476 189816 154488
rect 92900 154448 189816 154476
rect 92900 154436 92906 154448
rect 189810 154436 189816 154448
rect 189868 154436 189874 154488
rect 198734 154436 198740 154488
rect 198792 154476 198798 154488
rect 268838 154476 268844 154488
rect 198792 154448 268844 154476
rect 198792 154436 198798 154448
rect 268838 154436 268844 154448
rect 268896 154436 268902 154488
rect 274634 154436 274640 154488
rect 274692 154476 274698 154488
rect 310514 154476 310520 154488
rect 274692 154448 310520 154476
rect 274692 154436 274698 154448
rect 310514 154436 310520 154448
rect 310572 154436 310578 154488
rect 319990 154436 319996 154488
rect 320048 154476 320054 154488
rect 363230 154476 363236 154488
rect 320048 154448 363236 154476
rect 320048 154436 320054 154448
rect 363230 154436 363236 154448
rect 363288 154436 363294 154488
rect 366818 154436 366824 154488
rect 366876 154476 366882 154488
rect 395338 154476 395344 154488
rect 366876 154448 395344 154476
rect 366876 154436 366882 154448
rect 395338 154436 395344 154448
rect 395396 154436 395402 154488
rect 58342 154368 58348 154420
rect 58400 154408 58406 154420
rect 156598 154408 156604 154420
rect 58400 154380 156604 154408
rect 58400 154368 58406 154380
rect 156598 154368 156604 154380
rect 156656 154368 156662 154420
rect 192110 154368 192116 154420
rect 192168 154408 192174 154420
rect 265710 154408 265716 154420
rect 192168 154380 265716 154408
rect 192168 154368 192174 154380
rect 265710 154368 265716 154380
rect 265768 154368 265774 154420
rect 266998 154368 267004 154420
rect 267056 154408 267062 154420
rect 322842 154408 322848 154420
rect 267056 154380 322848 154408
rect 267056 154368 267062 154380
rect 322842 154368 322848 154380
rect 322900 154368 322906 154420
rect 335078 154368 335084 154420
rect 335136 154408 335142 154420
rect 338758 154408 338764 154420
rect 335136 154380 338764 154408
rect 335136 154368 335142 154380
rect 338758 154368 338764 154380
rect 338816 154368 338822 154420
rect 340966 154368 340972 154420
rect 341024 154408 341030 154420
rect 379238 154408 379244 154420
rect 341024 154380 379244 154408
rect 341024 154368 341030 154380
rect 379238 154368 379244 154380
rect 379296 154368 379302 154420
rect 51626 154300 51632 154352
rect 51684 154340 51690 154352
rect 158346 154340 158352 154352
rect 51684 154312 158352 154340
rect 51684 154300 51690 154312
rect 158346 154300 158352 154312
rect 158404 154300 158410 154352
rect 158438 154300 158444 154352
rect 158496 154340 158502 154352
rect 180242 154340 180248 154352
rect 158496 154312 180248 154340
rect 158496 154300 158502 154312
rect 180242 154300 180248 154312
rect 180300 154300 180306 154352
rect 185394 154300 185400 154352
rect 185452 154340 185458 154352
rect 260466 154340 260472 154352
rect 185452 154312 260472 154340
rect 185452 154300 185458 154312
rect 260466 154300 260472 154312
rect 260524 154300 260530 154352
rect 270310 154300 270316 154352
rect 270368 154340 270374 154352
rect 325326 154340 325332 154352
rect 270368 154312 325332 154340
rect 270368 154300 270374 154312
rect 325326 154300 325332 154312
rect 325384 154300 325390 154352
rect 326982 154300 326988 154352
rect 327040 154340 327046 154352
rect 368382 154340 368388 154352
rect 327040 154312 368388 154340
rect 327040 154300 327046 154312
rect 368382 154300 368388 154312
rect 368440 154300 368446 154352
rect 44910 154232 44916 154284
rect 44968 154272 44974 154284
rect 153194 154272 153200 154284
rect 44968 154244 153200 154272
rect 44968 154232 44974 154244
rect 153194 154232 153200 154244
rect 153252 154232 153258 154284
rect 154298 154232 154304 154284
rect 154356 154272 154362 154284
rect 183278 154272 183284 154284
rect 154356 154244 183284 154272
rect 154356 154232 154362 154244
rect 183278 154232 183284 154244
rect 183336 154232 183342 154284
rect 188798 154232 188804 154284
rect 188856 154272 188862 154284
rect 263042 154272 263048 154284
rect 188856 154244 263048 154272
rect 188856 154232 188862 154244
rect 263042 154232 263048 154244
rect 263100 154232 263106 154284
rect 263594 154232 263600 154284
rect 263652 154272 263658 154284
rect 320174 154272 320180 154284
rect 263652 154244 320180 154272
rect 263652 154232 263658 154244
rect 320174 154232 320180 154244
rect 320232 154232 320238 154284
rect 323302 154232 323308 154284
rect 323360 154272 323366 154284
rect 365714 154272 365720 154284
rect 323360 154244 365720 154272
rect 323360 154232 323366 154244
rect 365714 154232 365720 154244
rect 365772 154232 365778 154284
rect 371326 154232 371332 154284
rect 371384 154272 371390 154284
rect 402330 154272 402336 154284
rect 371384 154244 402336 154272
rect 371384 154232 371390 154244
rect 402330 154232 402336 154244
rect 402388 154232 402394 154284
rect 34790 154164 34796 154216
rect 34848 154204 34854 154216
rect 145558 154204 145564 154216
rect 34848 154176 145564 154204
rect 34848 154164 34854 154176
rect 145558 154164 145564 154176
rect 145616 154164 145622 154216
rect 147766 154164 147772 154216
rect 147824 154204 147830 154216
rect 177666 154204 177672 154216
rect 147824 154176 177672 154204
rect 147824 154164 147830 154176
rect 177666 154164 177672 154176
rect 177724 154164 177730 154216
rect 181990 154164 181996 154216
rect 182048 154204 182054 154216
rect 257890 154204 257896 154216
rect 182048 154176 257896 154204
rect 182048 154164 182054 154176
rect 257890 154164 257896 154176
rect 257948 154164 257954 154216
rect 257982 154164 257988 154216
rect 258040 154204 258046 154216
rect 315022 154204 315028 154216
rect 258040 154176 315028 154204
rect 258040 154164 258046 154176
rect 315022 154164 315028 154176
rect 315080 154164 315086 154216
rect 316586 154164 316592 154216
rect 316644 154204 316650 154216
rect 360654 154204 360660 154216
rect 316644 154176 360660 154204
rect 316644 154164 316650 154176
rect 360654 154164 360660 154176
rect 360712 154164 360718 154216
rect 368290 154164 368296 154216
rect 368348 154204 368354 154216
rect 399754 154204 399760 154216
rect 368348 154176 399760 154204
rect 368348 154164 368354 154176
rect 399754 154164 399760 154176
rect 399812 154164 399818 154216
rect 422570 154164 422576 154216
rect 422628 154204 422634 154216
rect 422628 154176 430068 154204
rect 422628 154164 422634 154176
rect 25590 154096 25596 154148
rect 25648 154136 25654 154148
rect 138474 154136 138480 154148
rect 25648 154108 138480 154136
rect 25648 154096 25654 154108
rect 138474 154096 138480 154108
rect 138532 154096 138538 154148
rect 156598 154096 156604 154148
rect 156656 154136 156662 154148
rect 163498 154136 163504 154148
rect 156656 154108 163504 154136
rect 156656 154096 156662 154108
rect 163498 154096 163504 154108
rect 163556 154096 163562 154148
rect 172422 154096 172428 154148
rect 172480 154136 172486 154148
rect 250162 154136 250168 154148
rect 172480 154108 250168 154136
rect 172480 154096 172486 154108
rect 250162 154096 250168 154108
rect 250220 154096 250226 154148
rect 250254 154096 250260 154148
rect 250312 154136 250318 154148
rect 309870 154136 309876 154148
rect 250312 154108 309876 154136
rect 250312 154096 250318 154108
rect 309870 154096 309876 154108
rect 309928 154096 309934 154148
rect 313274 154096 313280 154148
rect 313332 154136 313338 154148
rect 358078 154136 358084 154148
rect 313332 154108 358084 154136
rect 313332 154096 313338 154108
rect 358078 154096 358084 154108
rect 358136 154096 358142 154148
rect 360378 154096 360384 154148
rect 360436 154136 360442 154148
rect 394050 154136 394056 154148
rect 360436 154108 394056 154136
rect 360436 154096 360442 154108
rect 394050 154096 394056 154108
rect 394108 154096 394114 154148
rect 407482 154096 407488 154148
rect 407540 154136 407546 154148
rect 429930 154136 429936 154148
rect 407540 154108 429936 154136
rect 407540 154096 407546 154108
rect 429930 154096 429936 154108
rect 429988 154096 429994 154148
rect 13814 154028 13820 154080
rect 13872 154068 13878 154080
rect 129458 154068 129464 154080
rect 13872 154040 129464 154068
rect 13872 154028 13878 154040
rect 129458 154028 129464 154040
rect 129516 154028 129522 154080
rect 131114 154028 131120 154080
rect 131172 154068 131178 154080
rect 217410 154068 217416 154080
rect 131172 154040 217416 154068
rect 131172 154028 131178 154040
rect 217410 154028 217416 154040
rect 217468 154028 217474 154080
rect 219894 154028 219900 154080
rect 219952 154068 219958 154080
rect 286778 154068 286784 154080
rect 219952 154040 286784 154068
rect 219952 154028 219958 154040
rect 286778 154028 286784 154040
rect 286836 154028 286842 154080
rect 286870 154028 286876 154080
rect 286928 154068 286934 154080
rect 337470 154068 337476 154080
rect 286928 154040 337476 154068
rect 286928 154028 286934 154040
rect 337470 154028 337476 154040
rect 337528 154028 337534 154080
rect 338022 154028 338028 154080
rect 338080 154068 338086 154080
rect 376570 154068 376576 154080
rect 338080 154040 376576 154068
rect 338080 154028 338086 154040
rect 376570 154028 376576 154040
rect 376628 154028 376634 154080
rect 398190 154028 398196 154080
rect 398248 154068 398254 154080
rect 422938 154068 422944 154080
rect 398248 154040 422944 154068
rect 398248 154028 398254 154040
rect 422938 154028 422944 154040
rect 422996 154028 423002 154080
rect 430040 154068 430068 154176
rect 438854 154164 438860 154216
rect 438912 154204 438918 154216
rect 451826 154204 451832 154216
rect 438912 154176 451832 154204
rect 438912 154164 438918 154176
rect 451826 154164 451832 154176
rect 451884 154164 451890 154216
rect 431034 154096 431040 154148
rect 431092 154136 431098 154148
rect 447962 154136 447968 154148
rect 431092 154108 447968 154136
rect 431092 154096 431098 154108
rect 447962 154096 447968 154108
rect 448020 154096 448026 154148
rect 441430 154068 441436 154080
rect 430040 154040 441436 154068
rect 441430 154028 441436 154040
rect 441488 154028 441494 154080
rect 20530 153960 20536 154012
rect 20588 154000 20594 154012
rect 134610 154000 134616 154012
rect 20588 153972 134616 154000
rect 20588 153960 20594 153972
rect 134610 153960 134616 153972
rect 134668 153960 134674 154012
rect 143350 153960 143356 154012
rect 143408 154000 143414 154012
rect 228358 154000 228364 154012
rect 143408 153972 228364 154000
rect 143408 153960 143414 153972
rect 228358 153960 228364 153972
rect 228416 153960 228422 154012
rect 243446 153960 243452 154012
rect 243504 154000 243510 154012
rect 304718 154000 304724 154012
rect 243504 153972 304724 154000
rect 243504 153960 243510 153972
rect 304718 153960 304724 153972
rect 304776 153960 304782 154012
rect 304810 153960 304816 154012
rect 304868 154000 304874 154012
rect 349062 154000 349068 154012
rect 304868 153972 349068 154000
rect 304868 153960 304874 153972
rect 349062 153960 349068 153972
rect 349120 153960 349126 154012
rect 355318 153960 355324 154012
rect 355376 154000 355382 154012
rect 355376 153972 355640 154000
rect 355376 153960 355382 153972
rect 17126 153892 17132 153944
rect 17184 153932 17190 153944
rect 132034 153932 132040 153944
rect 17184 153904 132040 153932
rect 17184 153892 17190 153904
rect 132034 153892 132040 153904
rect 132092 153892 132098 153944
rect 135898 153892 135904 153944
rect 135956 153932 135962 153944
rect 222562 153932 222568 153944
rect 135956 153904 222568 153932
rect 135956 153892 135962 153904
rect 222562 153892 222568 153904
rect 222620 153892 222626 153944
rect 233326 153892 233332 153944
rect 233384 153932 233390 153944
rect 297082 153932 297088 153944
rect 233384 153904 297088 153932
rect 233384 153892 233390 153904
rect 297082 153892 297088 153904
rect 297140 153892 297146 153944
rect 309962 153892 309968 153944
rect 310020 153932 310026 153944
rect 355502 153932 355508 153944
rect 310020 153904 355508 153932
rect 310020 153892 310026 153904
rect 355502 153892 355508 153904
rect 355560 153892 355566 153944
rect 355612 153932 355640 153972
rect 357342 153960 357348 154012
rect 357400 154000 357406 154012
rect 391474 154000 391480 154012
rect 357400 153972 391480 154000
rect 357400 153960 357406 153972
rect 391474 153960 391480 153972
rect 391532 153960 391538 154012
rect 391842 153960 391848 154012
rect 391900 154000 391906 154012
rect 417786 154000 417792 154012
rect 391900 153972 417792 154000
rect 391900 153960 391906 153972
rect 417786 153960 417792 153972
rect 417844 153960 417850 154012
rect 425238 153960 425244 154012
rect 425296 154000 425302 154012
rect 443454 154000 443460 154012
rect 425296 153972 443460 154000
rect 425296 153960 425302 153972
rect 443454 153960 443460 153972
rect 443512 153960 443518 154012
rect 390186 153932 390192 153944
rect 355612 153904 390192 153932
rect 390186 153892 390192 153904
rect 390244 153892 390250 153944
rect 390646 153892 390652 153944
rect 390704 153932 390710 153944
rect 417142 153932 417148 153944
rect 390704 153904 417148 153932
rect 390704 153892 390710 153904
rect 417142 153892 417148 153904
rect 417200 153892 417206 153944
rect 418430 153892 418436 153944
rect 418488 153932 418494 153944
rect 438302 153932 438308 153944
rect 418488 153904 438308 153932
rect 418488 153892 418494 153904
rect 438302 153892 438308 153904
rect 438360 153892 438366 153944
rect 440234 153892 440240 153944
rect 440292 153932 440298 153944
rect 455046 153932 455052 153944
rect 440292 153904 455052 153932
rect 440292 153892 440298 153904
rect 455046 153892 455052 153904
rect 455104 153892 455110 153944
rect 4062 153824 4068 153876
rect 4120 153864 4126 153876
rect 121730 153864 121736 153876
rect 4120 153836 121736 153864
rect 4120 153824 4126 153836
rect 121730 153824 121736 153836
rect 121788 153824 121794 153876
rect 122650 153824 122656 153876
rect 122708 153864 122714 153876
rect 212258 153864 212264 153876
rect 122708 153836 212264 153864
rect 122708 153824 122714 153836
rect 212258 153824 212264 153836
rect 212316 153824 212322 153876
rect 213178 153824 213184 153876
rect 213236 153864 213242 153876
rect 281626 153864 281632 153876
rect 213236 153836 281632 153864
rect 213236 153824 213242 153836
rect 281626 153824 281632 153836
rect 281684 153824 281690 153876
rect 282546 153824 282552 153876
rect 282604 153864 282610 153876
rect 333698 153864 333704 153876
rect 282604 153836 333704 153864
rect 282604 153824 282610 153836
rect 333698 153824 333704 153836
rect 333756 153824 333762 153876
rect 373442 153864 373448 153876
rect 335326 153836 373448 153864
rect 105446 153756 105452 153808
rect 105504 153796 105510 153808
rect 199470 153796 199476 153808
rect 105504 153768 199476 153796
rect 105504 153756 105510 153768
rect 199470 153756 199476 153768
rect 199528 153756 199534 153808
rect 208486 153756 208492 153808
rect 208544 153796 208550 153808
rect 273898 153796 273904 153808
rect 208544 153768 273904 153796
rect 208544 153756 208550 153768
rect 273898 153756 273904 153768
rect 273956 153756 273962 153808
rect 280062 153756 280068 153808
rect 280120 153796 280126 153808
rect 315666 153796 315672 153808
rect 280120 153768 315672 153796
rect 280120 153756 280126 153768
rect 315666 153756 315672 153768
rect 315724 153756 315730 153808
rect 333422 153756 333428 153808
rect 333480 153796 333486 153808
rect 335326 153796 335354 153836
rect 373442 153824 373448 153836
rect 373500 153824 373506 153876
rect 380802 153824 380808 153876
rect 380860 153864 380866 153876
rect 409414 153864 409420 153876
rect 380860 153836 409420 153864
rect 380860 153824 380866 153836
rect 409414 153824 409420 153836
rect 409472 153824 409478 153876
rect 417510 153824 417516 153876
rect 417568 153864 417574 153876
rect 437658 153864 437664 153876
rect 417568 153836 437664 153864
rect 417568 153824 417574 153836
rect 437658 153824 437664 153836
rect 437716 153824 437722 153876
rect 438578 153824 438584 153876
rect 438636 153864 438642 153876
rect 453758 153864 453764 153876
rect 438636 153836 453764 153864
rect 438636 153824 438642 153836
rect 453758 153824 453764 153836
rect 453816 153824 453822 153876
rect 333480 153768 335354 153796
rect 333480 153756 333486 153768
rect 63402 153688 63408 153740
rect 63460 153728 63466 153740
rect 118694 153728 118700 153740
rect 63460 153700 118700 153728
rect 63460 153688 63466 153700
rect 118694 153688 118700 153700
rect 118752 153688 118758 153740
rect 119798 153688 119804 153740
rect 119856 153728 119862 153740
rect 208394 153728 208400 153740
rect 119856 153700 208400 153728
rect 119856 153688 119862 153700
rect 208394 153688 208400 153700
rect 208452 153688 208458 153740
rect 244274 153688 244280 153740
rect 244332 153728 244338 153740
rect 305362 153728 305368 153740
rect 244332 153700 305368 153728
rect 244332 153688 244338 153700
rect 305362 153688 305368 153700
rect 305420 153688 305426 153740
rect 305454 153688 305460 153740
rect 305512 153728 305518 153740
rect 336182 153728 336188 153740
rect 305512 153700 336188 153728
rect 305512 153688 305518 153700
rect 336182 153688 336188 153700
rect 336240 153688 336246 153740
rect 128354 153620 128360 153672
rect 128412 153660 128418 153672
rect 159634 153660 159640 153672
rect 128412 153632 159640 153660
rect 128412 153620 128418 153632
rect 159634 153620 159640 153632
rect 159692 153620 159698 153672
rect 168558 153620 168564 153672
rect 168616 153660 168622 153672
rect 215294 153660 215300 153672
rect 168616 153632 215300 153660
rect 168616 153620 168622 153632
rect 215294 153620 215300 153632
rect 215352 153620 215358 153672
rect 263594 153620 263600 153672
rect 263652 153660 263658 153672
rect 263778 153660 263784 153672
rect 263652 153632 263784 153660
rect 263652 153620 263658 153632
rect 263778 153620 263784 153632
rect 263836 153620 263842 153672
rect 296806 153620 296812 153672
rect 296864 153660 296870 153672
rect 325970 153660 325976 153672
rect 296864 153632 325976 153660
rect 296864 153620 296870 153632
rect 325970 153620 325976 153632
rect 326028 153620 326034 153672
rect 197630 153552 197636 153604
rect 197688 153592 197694 153604
rect 238018 153592 238024 153604
rect 197688 153564 238024 153592
rect 197688 153552 197694 153564
rect 238018 153552 238024 153564
rect 238076 153552 238082 153604
rect 109034 153144 109040 153196
rect 109092 153184 109098 153196
rect 198182 153184 198188 153196
rect 109092 153156 198188 153184
rect 109092 153144 109098 153156
rect 198182 153144 198188 153156
rect 198240 153144 198246 153196
rect 202966 153144 202972 153196
rect 203024 153184 203030 153196
rect 252094 153184 252100 153196
rect 203024 153156 252100 153184
rect 203024 153144 203030 153156
rect 252094 153144 252100 153156
rect 252152 153144 252158 153196
rect 259638 153144 259644 153196
rect 259696 153184 259702 153196
rect 270126 153184 270132 153196
rect 259696 153156 270132 153184
rect 259696 153144 259702 153156
rect 270126 153144 270132 153156
rect 270184 153144 270190 153196
rect 272518 153144 272524 153196
rect 272576 153184 272582 153196
rect 285490 153184 285496 153196
rect 272576 153156 285496 153184
rect 272576 153144 272582 153156
rect 285490 153144 285496 153156
rect 285548 153144 285554 153196
rect 292298 153144 292304 153196
rect 292356 153184 292362 153196
rect 339402 153184 339408 153196
rect 292356 153156 339408 153184
rect 292356 153144 292362 153156
rect 339402 153144 339408 153156
rect 339460 153144 339466 153196
rect 355226 153144 355232 153196
rect 355284 153184 355290 153196
rect 357434 153184 357440 153196
rect 355284 153156 357440 153184
rect 355284 153144 355290 153156
rect 357434 153144 357440 153156
rect 357492 153144 357498 153196
rect 368474 153144 368480 153196
rect 368532 153184 368538 153196
rect 372798 153184 372804 153196
rect 368532 153156 372804 153184
rect 368532 153144 368538 153156
rect 372798 153144 372804 153156
rect 372856 153144 372862 153196
rect 385954 153144 385960 153196
rect 386012 153184 386018 153196
rect 388254 153184 388260 153196
rect 386012 153156 388260 153184
rect 386012 153144 386018 153156
rect 388254 153144 388260 153156
rect 388312 153144 388318 153196
rect 408494 153144 408500 153196
rect 408552 153184 408558 153196
rect 410702 153184 410708 153196
rect 408552 153156 410708 153184
rect 408552 153144 408558 153156
rect 410702 153144 410708 153156
rect 410760 153144 410766 153196
rect 435818 153144 435824 153196
rect 435876 153184 435882 153196
rect 439590 153184 439596 153196
rect 435876 153156 439596 153184
rect 435876 153144 435882 153156
rect 439590 153144 439596 153156
rect 439648 153144 439654 153196
rect 447134 153144 447140 153196
rect 447192 153184 447198 153196
rect 449250 153184 449256 153196
rect 447192 153156 449256 153184
rect 447192 153144 447198 153156
rect 449250 153144 449256 153156
rect 449308 153144 449314 153196
rect 461578 153144 461584 153196
rect 461636 153184 461642 153196
rect 465902 153184 465908 153196
rect 461636 153156 465908 153184
rect 461636 153144 461642 153156
rect 465902 153144 465908 153156
rect 465960 153144 465966 153196
rect 466454 153144 466460 153196
rect 466512 153184 466518 153196
rect 469766 153184 469772 153196
rect 466512 153156 469772 153184
rect 466512 153144 466518 153156
rect 469766 153144 469772 153156
rect 469824 153144 469830 153196
rect 471606 153144 471612 153196
rect 471664 153184 471670 153196
rect 473630 153184 473636 153196
rect 471664 153156 473636 153184
rect 471664 153144 471670 153156
rect 473630 153144 473636 153156
rect 473688 153144 473694 153196
rect 474826 153144 474832 153196
rect 474884 153184 474890 153196
rect 476942 153184 476948 153196
rect 474884 153156 476948 153184
rect 474884 153144 474890 153156
rect 476942 153144 476948 153156
rect 477000 153144 477006 153196
rect 485682 153144 485688 153196
rect 485740 153184 485746 153196
rect 489638 153184 489644 153196
rect 485740 153156 489644 153184
rect 485740 153144 485746 153156
rect 489638 153144 489644 153156
rect 489696 153144 489702 153196
rect 490742 153144 490748 153196
rect 490800 153184 490806 153196
rect 493502 153184 493508 153196
rect 490800 153156 493508 153184
rect 490800 153144 490806 153156
rect 493502 153144 493508 153156
rect 493560 153144 493566 153196
rect 494054 153144 494060 153196
rect 494112 153184 494118 153196
rect 496078 153184 496084 153196
rect 494112 153156 496084 153184
rect 494112 153144 494118 153156
rect 496078 153144 496084 153156
rect 496136 153144 496142 153196
rect 496630 153144 496636 153196
rect 496688 153184 496694 153196
rect 498010 153184 498016 153196
rect 496688 153156 498016 153184
rect 496688 153144 496694 153156
rect 498010 153144 498016 153156
rect 498068 153144 498074 153196
rect 498286 153144 498292 153196
rect 498344 153184 498350 153196
rect 499298 153184 499304 153196
rect 498344 153156 499304 153184
rect 498344 153144 498350 153156
rect 499298 153144 499304 153156
rect 499356 153144 499362 153196
rect 500954 153144 500960 153196
rect 501012 153184 501018 153196
rect 501874 153184 501880 153196
rect 501012 153156 501880 153184
rect 501012 153144 501018 153156
rect 501874 153144 501880 153156
rect 501932 153144 501938 153196
rect 510982 153144 510988 153196
rect 511040 153184 511046 153196
rect 513466 153184 513472 153196
rect 511040 153156 513472 153184
rect 511040 153144 511046 153156
rect 513466 153144 513472 153156
rect 513524 153144 513530 153196
rect 514202 153144 514208 153196
rect 514260 153184 514266 153196
rect 517422 153184 517428 153196
rect 514260 153156 517428 153184
rect 514260 153144 514266 153156
rect 517422 153144 517428 153156
rect 517480 153144 517486 153196
rect 117222 153076 117228 153128
rect 117280 153116 117286 153128
rect 208486 153116 208492 153128
rect 117280 153088 208492 153116
rect 117280 153076 117286 153088
rect 208486 153076 208492 153088
rect 208544 153076 208550 153128
rect 215294 153076 215300 153128
rect 215352 153116 215358 153128
rect 247586 153116 247592 153128
rect 215352 153088 247592 153116
rect 215352 153076 215358 153088
rect 247586 153076 247592 153088
rect 247644 153076 247650 153128
rect 252002 153076 252008 153128
rect 252060 153116 252066 153128
rect 301590 153116 301596 153128
rect 252060 153088 301596 153116
rect 252060 153076 252066 153088
rect 301590 153076 301596 153088
rect 301648 153076 301654 153128
rect 301682 153076 301688 153128
rect 301740 153116 301746 153128
rect 311158 153116 311164 153128
rect 301740 153088 311164 153116
rect 301740 153076 301746 153088
rect 311158 153076 311164 153088
rect 311216 153076 311222 153128
rect 321462 153116 321468 153128
rect 311866 153088 321468 153116
rect 113910 153008 113916 153060
rect 113968 153048 113974 153060
rect 205910 153048 205916 153060
rect 113968 153020 205916 153048
rect 113968 153008 113974 153020
rect 205910 153008 205916 153020
rect 205968 153008 205974 153060
rect 216766 153008 216772 153060
rect 216824 153048 216830 153060
rect 239306 153048 239312 153060
rect 216824 153020 239312 153048
rect 216824 153008 216830 153020
rect 239306 153008 239312 153020
rect 239364 153008 239370 153060
rect 239950 153008 239956 153060
rect 240008 153048 240014 153060
rect 293218 153048 293224 153060
rect 240008 153020 293224 153048
rect 240008 153008 240014 153020
rect 293218 153008 293224 153020
rect 293276 153008 293282 153060
rect 298738 153008 298744 153060
rect 298796 153048 298802 153060
rect 306006 153048 306012 153060
rect 298796 153020 306012 153048
rect 298796 153008 298802 153020
rect 306006 153008 306012 153020
rect 306064 153008 306070 153060
rect 311066 153008 311072 153060
rect 311124 153048 311130 153060
rect 311866 153048 311894 153088
rect 321462 153076 321468 153088
rect 321520 153076 321526 153128
rect 338758 153076 338764 153128
rect 338816 153116 338822 153128
rect 374730 153116 374736 153128
rect 338816 153088 374736 153116
rect 338816 153076 338822 153088
rect 374730 153076 374736 153088
rect 374788 153076 374794 153128
rect 463142 153076 463148 153128
rect 463200 153116 463206 153128
rect 467190 153116 467196 153128
rect 463200 153088 467196 153116
rect 463200 153076 463206 153088
rect 467190 153076 467196 153088
rect 467248 153076 467254 153128
rect 471974 153076 471980 153128
rect 472032 153116 472038 153128
rect 474274 153116 474280 153128
rect 472032 153088 474280 153116
rect 472032 153076 472038 153088
rect 474274 153076 474280 153088
rect 474332 153076 474338 153128
rect 476114 153076 476120 153128
rect 476172 153116 476178 153128
rect 478138 153116 478144 153128
rect 476172 153088 478144 153116
rect 476172 153076 476178 153088
rect 478138 153076 478144 153088
rect 478196 153076 478202 153128
rect 484854 153076 484860 153128
rect 484912 153116 484918 153128
rect 488994 153116 489000 153128
rect 484912 153088 489000 153116
rect 484912 153076 484918 153088
rect 488994 153076 489000 153088
rect 489052 153076 489058 153128
rect 489914 153076 489920 153128
rect 489972 153116 489978 153128
rect 492858 153116 492864 153128
rect 489972 153088 492864 153116
rect 489972 153076 489978 153088
rect 492858 153076 492864 153088
rect 492916 153076 492922 153128
rect 493226 153076 493232 153128
rect 493284 153116 493290 153128
rect 495434 153116 495440 153128
rect 493284 153088 495440 153116
rect 493284 153076 493290 153088
rect 495434 153076 495440 153088
rect 495492 153076 495498 153128
rect 495802 153076 495808 153128
rect 495860 153116 495866 153128
rect 497366 153116 497372 153128
rect 495860 153088 497372 153116
rect 495860 153076 495866 153088
rect 497366 153076 497372 153088
rect 497424 153076 497430 153128
rect 497458 153076 497464 153128
rect 497516 153116 497522 153128
rect 498654 153116 498660 153128
rect 497516 153088 498660 153116
rect 497516 153076 497522 153088
rect 498654 153076 498660 153088
rect 498712 153076 498718 153128
rect 512914 153076 512920 153128
rect 512972 153116 512978 153128
rect 515306 153116 515312 153128
rect 512972 153088 515312 153116
rect 512972 153076 512978 153088
rect 515306 153076 515312 153088
rect 515364 153076 515370 153128
rect 311124 153020 311894 153048
rect 311124 153008 311130 153020
rect 318702 153008 318708 153060
rect 318760 153048 318766 153060
rect 360010 153048 360016 153060
rect 318760 153020 360016 153048
rect 318760 153008 318766 153020
rect 360010 153008 360016 153020
rect 360068 153008 360074 153060
rect 399018 153008 399024 153060
rect 399076 153048 399082 153060
rect 423582 153048 423588 153060
rect 399076 153020 423588 153048
rect 399076 153008 399082 153020
rect 423582 153008 423588 153020
rect 423640 153008 423646 153060
rect 462958 153008 462964 153060
rect 463016 153048 463022 153060
rect 466546 153048 466552 153060
rect 463016 153020 466552 153048
rect 463016 153008 463022 153020
rect 466546 153008 466552 153020
rect 466604 153008 466610 153060
rect 466638 153008 466644 153060
rect 466696 153048 466702 153060
rect 470410 153048 470416 153060
rect 466696 153020 470416 153048
rect 466696 153008 466702 153020
rect 470410 153008 470416 153020
rect 470468 153008 470474 153060
rect 472802 153008 472808 153060
rect 472860 153048 472866 153060
rect 474918 153048 474924 153060
rect 472860 153020 474924 153048
rect 472860 153008 472866 153020
rect 474918 153008 474924 153020
rect 474976 153008 474982 153060
rect 484302 153008 484308 153060
rect 484360 153048 484366 153060
rect 488258 153048 488264 153060
rect 484360 153020 488264 153048
rect 484360 153008 484366 153020
rect 488258 153008 488264 153020
rect 488316 153008 488322 153060
rect 492398 153008 492404 153060
rect 492456 153048 492462 153060
rect 494790 153048 494796 153060
rect 492456 153020 494796 153048
rect 492456 153008 492462 153020
rect 494790 153008 494796 153020
rect 494848 153008 494854 153060
rect 495250 153008 495256 153060
rect 495308 153048 495314 153060
rect 496722 153048 496728 153060
rect 495308 153020 496728 153048
rect 495308 153008 495314 153020
rect 496722 153008 496728 153020
rect 496780 153008 496786 153060
rect 107470 152940 107476 152992
rect 107528 152980 107534 152992
rect 200758 152980 200764 152992
rect 107528 152952 200764 152980
rect 107528 152940 107534 152952
rect 200758 152940 200764 152952
rect 200816 152940 200822 152992
rect 205634 152940 205640 152992
rect 205692 152980 205698 152992
rect 212902 152980 212908 152992
rect 205692 152952 212908 152980
rect 205692 152940 205698 152952
rect 212902 152940 212908 152952
rect 212960 152940 212966 152992
rect 213638 152940 213644 152992
rect 213696 152980 213702 152992
rect 267550 152980 267556 152992
rect 213696 152952 267556 152980
rect 213696 152940 213702 152952
rect 267550 152940 267556 152952
rect 267608 152940 267614 152992
rect 271690 152940 271696 152992
rect 271748 152980 271754 152992
rect 324038 152980 324044 152992
rect 271748 152952 324044 152980
rect 271748 152940 271754 152952
rect 324038 152940 324044 152952
rect 324096 152940 324102 152992
rect 337930 152940 337936 152992
rect 337988 152980 337994 152992
rect 375374 152980 375380 152992
rect 337988 152952 375380 152980
rect 337988 152940 337994 152952
rect 375374 152940 375380 152952
rect 375432 152940 375438 152992
rect 389082 152940 389088 152992
rect 389140 152980 389146 152992
rect 413278 152980 413284 152992
rect 389140 152952 413284 152980
rect 389140 152940 389146 152952
rect 413278 152940 413284 152952
rect 413336 152940 413342 152992
rect 415854 152940 415860 152992
rect 415912 152980 415918 152992
rect 436370 152980 436376 152992
rect 415912 152952 436376 152980
rect 415912 152940 415918 152952
rect 436370 152940 436376 152952
rect 436428 152940 436434 152992
rect 465074 152940 465080 152992
rect 465132 152980 465138 152992
rect 469122 152980 469128 152992
rect 465132 152952 469128 152980
rect 465132 152940 465138 152952
rect 469122 152940 469128 152952
rect 469180 152940 469186 152992
rect 471790 152940 471796 152992
rect 471848 152980 471854 152992
rect 472986 152980 472992 152992
rect 471848 152952 472992 152980
rect 471848 152940 471854 152952
rect 472986 152940 472992 152952
rect 473044 152940 473050 152992
rect 473354 152940 473360 152992
rect 473412 152980 473418 152992
rect 475562 152980 475568 152992
rect 473412 152952 475568 152980
rect 473412 152940 473418 152952
rect 475562 152940 475568 152952
rect 475620 152940 475626 152992
rect 483198 152940 483204 152992
rect 483256 152980 483262 152992
rect 487798 152980 487804 152992
rect 483256 152952 487804 152980
rect 483256 152940 483262 152952
rect 487798 152940 487804 152952
rect 487856 152940 487862 152992
rect 491570 152940 491576 152992
rect 491628 152980 491634 152992
rect 494146 152980 494152 152992
rect 491628 152952 494152 152980
rect 491628 152940 491634 152952
rect 494146 152940 494152 152952
rect 494204 152940 494210 152992
rect 512270 152940 512276 152992
rect 512328 152980 512334 152992
rect 514754 152980 514760 152992
rect 512328 152952 514760 152980
rect 512328 152940 512334 152952
rect 514754 152940 514760 152952
rect 514812 152940 514818 152992
rect 97074 152872 97080 152924
rect 97132 152912 97138 152924
rect 193030 152912 193036 152924
rect 97132 152884 193036 152912
rect 97132 152872 97138 152884
rect 193030 152872 193036 152884
rect 193088 152872 193094 152924
rect 210142 152872 210148 152924
rect 210200 152912 210206 152924
rect 262398 152912 262404 152924
rect 210200 152884 262404 152912
rect 210200 152872 210206 152884
rect 262398 152872 262404 152884
rect 262456 152872 262462 152924
rect 263410 152872 263416 152924
rect 263468 152912 263474 152924
rect 318886 152912 318892 152924
rect 263468 152884 318892 152912
rect 263468 152872 263474 152884
rect 318886 152872 318892 152884
rect 318944 152872 318950 152924
rect 328270 152872 328276 152924
rect 328328 152912 328334 152924
rect 369578 152912 369584 152924
rect 328328 152884 369584 152912
rect 328328 152872 328334 152884
rect 369578 152872 369584 152884
rect 369636 152872 369642 152924
rect 372614 152872 372620 152924
rect 372672 152912 372678 152924
rect 380526 152912 380532 152924
rect 372672 152884 380532 152912
rect 372672 152872 372678 152884
rect 380526 152872 380532 152884
rect 380584 152872 380590 152924
rect 380986 152872 380992 152924
rect 381044 152912 381050 152924
rect 408126 152912 408132 152924
rect 381044 152884 408132 152912
rect 381044 152872 381050 152884
rect 408126 152872 408132 152884
rect 408184 152872 408190 152924
rect 409966 152872 409972 152924
rect 410024 152912 410030 152924
rect 431862 152912 431868 152924
rect 410024 152884 431868 152912
rect 410024 152872 410030 152884
rect 431862 152872 431868 152884
rect 431920 152872 431926 152924
rect 464706 152872 464712 152924
rect 464764 152912 464770 152924
rect 468386 152912 468392 152924
rect 464764 152884 468392 152912
rect 464764 152872 464770 152884
rect 468386 152872 468392 152884
rect 468444 152872 468450 152924
rect 90358 152804 90364 152856
rect 90416 152844 90422 152856
rect 187878 152844 187884 152856
rect 90416 152816 187884 152844
rect 90416 152804 90422 152816
rect 187878 152804 187884 152816
rect 187936 152804 187942 152856
rect 192570 152804 192576 152856
rect 192628 152844 192634 152856
rect 229002 152844 229008 152856
rect 192628 152816 229008 152844
rect 192628 152804 192634 152816
rect 229002 152804 229008 152816
rect 229060 152804 229066 152856
rect 244642 152804 244648 152856
rect 244700 152844 244706 152856
rect 303522 152844 303528 152856
rect 244700 152816 303528 152844
rect 244700 152804 244706 152816
rect 303522 152804 303528 152816
rect 303580 152804 303586 152856
rect 304994 152804 305000 152856
rect 305052 152844 305058 152856
rect 316310 152844 316316 152856
rect 305052 152816 316316 152844
rect 305052 152804 305058 152816
rect 316310 152804 316316 152816
rect 316368 152804 316374 152856
rect 322750 152804 322756 152856
rect 322808 152844 322814 152856
rect 365162 152844 365168 152856
rect 322808 152816 365168 152844
rect 322808 152804 322814 152816
rect 365162 152804 365168 152816
rect 365220 152804 365226 152856
rect 374270 152804 374276 152856
rect 374328 152844 374334 152856
rect 402974 152844 402980 152856
rect 374328 152816 402980 152844
rect 374328 152804 374334 152816
rect 402974 152804 402980 152816
rect 403032 152804 403038 152856
rect 412542 152804 412548 152856
rect 412600 152844 412606 152856
rect 433794 152844 433800 152856
rect 412600 152816 433800 152844
rect 412600 152804 412606 152816
rect 433794 152804 433800 152816
rect 433852 152804 433858 152856
rect 510338 152804 510344 152856
rect 510396 152844 510402 152856
rect 511994 152844 512000 152856
rect 510396 152816 512000 152844
rect 510396 152804 510402 152816
rect 511994 152804 512000 152816
rect 512052 152804 512058 152856
rect 84102 152736 84108 152788
rect 84160 152776 84166 152788
rect 182726 152776 182732 152788
rect 84160 152748 182732 152776
rect 84160 152736 84166 152748
rect 182726 152736 182732 152748
rect 182784 152736 182790 152788
rect 187694 152736 187700 152788
rect 187752 152776 187758 152788
rect 213546 152776 213552 152788
rect 187752 152748 213552 152776
rect 187752 152736 187758 152748
rect 213546 152736 213552 152748
rect 213604 152736 213610 152788
rect 222010 152736 222016 152788
rect 222068 152776 222074 152788
rect 224494 152776 224500 152788
rect 222068 152748 224500 152776
rect 222068 152736 222074 152748
rect 224494 152736 224500 152748
rect 224552 152736 224558 152788
rect 224586 152736 224592 152788
rect 224644 152776 224650 152788
rect 282914 152776 282920 152788
rect 224644 152748 282920 152776
rect 224644 152736 224650 152748
rect 282914 152736 282920 152748
rect 282972 152736 282978 152788
rect 284386 152736 284392 152788
rect 284444 152776 284450 152788
rect 295794 152776 295800 152788
rect 284444 152748 295800 152776
rect 284444 152736 284450 152748
rect 295794 152736 295800 152748
rect 295852 152736 295858 152788
rect 295886 152736 295892 152788
rect 295944 152776 295950 152788
rect 344554 152776 344560 152788
rect 295944 152748 344560 152776
rect 295944 152736 295950 152748
rect 344554 152736 344560 152748
rect 344612 152736 344618 152788
rect 358814 152736 358820 152788
rect 358872 152776 358878 152788
rect 390830 152776 390836 152788
rect 358872 152748 390836 152776
rect 358872 152736 358878 152748
rect 390830 152736 390836 152748
rect 390888 152736 390894 152788
rect 391566 152736 391572 152788
rect 391624 152776 391630 152788
rect 416498 152776 416504 152788
rect 391624 152748 416504 152776
rect 391624 152736 391630 152748
rect 416498 152736 416504 152748
rect 416556 152736 416562 152788
rect 416682 152736 416688 152788
rect 416740 152776 416746 152788
rect 437014 152776 437020 152788
rect 416740 152748 437020 152776
rect 416740 152736 416746 152748
rect 437014 152736 437020 152748
rect 437072 152736 437078 152788
rect 73522 152668 73528 152720
rect 73580 152708 73586 152720
rect 175090 152708 175096 152720
rect 73580 152680 175096 152708
rect 73580 152668 73586 152680
rect 175090 152668 175096 152680
rect 175148 152668 175154 152720
rect 179414 152668 179420 152720
rect 179472 152708 179478 152720
rect 195606 152708 195612 152720
rect 179472 152680 195612 152708
rect 179472 152668 179478 152680
rect 195606 152668 195612 152680
rect 195664 152668 195670 152720
rect 211890 152668 211896 152720
rect 211948 152708 211954 152720
rect 272702 152708 272708 152720
rect 211948 152680 272708 152708
rect 211948 152668 211954 152680
rect 272702 152668 272708 152680
rect 272760 152668 272766 152720
rect 278314 152668 278320 152720
rect 278372 152708 278378 152720
rect 329190 152708 329196 152720
rect 278372 152680 329196 152708
rect 278372 152668 278378 152680
rect 329190 152668 329196 152680
rect 329248 152668 329254 152720
rect 329282 152668 329288 152720
rect 329340 152708 329346 152720
rect 370222 152708 370228 152720
rect 329340 152680 370228 152708
rect 329340 152668 329346 152680
rect 370222 152668 370228 152680
rect 370280 152668 370286 152720
rect 376662 152668 376668 152720
rect 376720 152708 376726 152720
rect 406194 152708 406200 152720
rect 376720 152680 406200 152708
rect 376720 152668 376726 152680
rect 406194 152668 406200 152680
rect 406252 152668 406258 152720
rect 407022 152668 407028 152720
rect 407080 152708 407086 152720
rect 428642 152708 428648 152720
rect 407080 152680 428648 152708
rect 407080 152668 407086 152680
rect 428642 152668 428648 152680
rect 428700 152668 428706 152720
rect 444282 152668 444288 152720
rect 444340 152708 444346 152720
rect 453114 152708 453120 152720
rect 444340 152680 453120 152708
rect 444340 152668 444346 152680
rect 453114 152668 453120 152680
rect 453172 152668 453178 152720
rect 34422 152600 34428 152652
rect 34480 152640 34486 152652
rect 144914 152640 144920 152652
rect 34480 152612 144920 152640
rect 34480 152600 34486 152612
rect 144914 152600 144920 152612
rect 144972 152600 144978 152652
rect 167730 152600 167736 152652
rect 167788 152640 167794 152652
rect 246942 152640 246948 152652
rect 167788 152612 246948 152640
rect 167788 152600 167794 152612
rect 246942 152600 246948 152612
rect 247000 152600 247006 152652
rect 255222 152600 255228 152652
rect 255280 152640 255286 152652
rect 313734 152640 313740 152652
rect 255280 152612 313740 152640
rect 255280 152600 255286 152612
rect 313734 152600 313740 152612
rect 313792 152600 313798 152652
rect 314930 152600 314936 152652
rect 314988 152640 314994 152652
rect 359366 152640 359372 152652
rect 314988 152612 359372 152640
rect 314988 152600 314994 152612
rect 359366 152600 359372 152612
rect 359424 152600 359430 152652
rect 362954 152600 362960 152652
rect 363012 152640 363018 152652
rect 395982 152640 395988 152652
rect 363012 152612 395988 152640
rect 363012 152600 363018 152612
rect 395982 152600 395988 152612
rect 396040 152600 396046 152652
rect 396626 152600 396632 152652
rect 396684 152640 396690 152652
rect 421650 152640 421656 152652
rect 396684 152612 421656 152640
rect 396684 152600 396690 152612
rect 421650 152600 421656 152612
rect 421708 152600 421714 152652
rect 445662 152600 445668 152652
rect 445720 152640 445726 152652
rect 455690 152640 455696 152652
rect 445720 152612 455696 152640
rect 445720 152600 445726 152612
rect 455690 152600 455696 152612
rect 455748 152600 455754 152652
rect 23382 152532 23388 152584
rect 23440 152572 23446 152584
rect 136542 152572 136548 152584
rect 23440 152544 136548 152572
rect 23440 152532 23446 152544
rect 136542 152532 136548 152544
rect 136600 152532 136606 152584
rect 147582 152532 147588 152584
rect 147640 152572 147646 152584
rect 231578 152572 231584 152584
rect 147640 152544 231584 152572
rect 147640 152532 147646 152544
rect 231578 152532 231584 152544
rect 231636 152532 231642 152584
rect 248506 152532 248512 152584
rect 248564 152572 248570 152584
rect 308582 152572 308588 152584
rect 248564 152544 308588 152572
rect 248564 152532 248570 152544
rect 308582 152532 308588 152544
rect 308640 152532 308646 152584
rect 309042 152532 309048 152584
rect 309100 152572 309106 152584
rect 354858 152572 354864 152584
rect 309100 152544 354864 152572
rect 309100 152532 309106 152544
rect 354858 152532 354864 152544
rect 354916 152532 354922 152584
rect 365438 152532 365444 152584
rect 365496 152572 365502 152584
rect 397822 152572 397828 152584
rect 365496 152544 397828 152572
rect 365496 152532 365502 152544
rect 397822 152532 397828 152544
rect 397880 152532 397886 152584
rect 403250 152532 403256 152584
rect 403308 152572 403314 152584
rect 426802 152572 426808 152584
rect 403308 152544 426808 152572
rect 403308 152532 403314 152544
rect 426802 152532 426808 152544
rect 426860 152532 426866 152584
rect 446950 152532 446956 152584
rect 447008 152572 447014 152584
rect 460014 152572 460020 152584
rect 447008 152544 460020 152572
rect 447008 152532 447014 152544
rect 460014 152532 460020 152544
rect 460072 152532 460078 152584
rect 460106 152532 460112 152584
rect 460164 152572 460170 152584
rect 464614 152572 464620 152584
rect 460164 152544 464620 152572
rect 460164 152532 460170 152544
rect 464614 152532 464620 152544
rect 464672 152532 464678 152584
rect 6270 152464 6276 152516
rect 6328 152504 6334 152516
rect 123662 152504 123668 152516
rect 6328 152476 123668 152504
rect 6328 152464 6334 152476
rect 123662 152464 123668 152476
rect 123720 152464 123726 152516
rect 125686 152464 125692 152516
rect 125744 152504 125750 152516
rect 127526 152504 127532 152516
rect 125744 152476 127532 152504
rect 125744 152464 125750 152476
rect 127526 152464 127532 152476
rect 127584 152464 127590 152516
rect 134058 152464 134064 152516
rect 134116 152504 134122 152516
rect 221274 152504 221280 152516
rect 134116 152476 221280 152504
rect 134116 152464 134122 152476
rect 221274 152464 221280 152476
rect 221332 152464 221338 152516
rect 234982 152464 234988 152516
rect 235040 152504 235046 152516
rect 298370 152504 298376 152516
rect 235040 152476 298376 152504
rect 235040 152464 235046 152476
rect 298370 152464 298376 152476
rect 298428 152464 298434 152516
rect 302326 152464 302332 152516
rect 302384 152504 302390 152516
rect 349706 152504 349712 152516
rect 302384 152476 349712 152504
rect 302384 152464 302390 152476
rect 349706 152464 349712 152476
rect 349764 152464 349770 152516
rect 385586 152504 385592 152516
rect 354646 152476 385592 152504
rect 109126 152396 109132 152448
rect 109184 152436 109190 152448
rect 122374 152436 122380 152448
rect 109184 152408 122380 152436
rect 109184 152396 109190 152408
rect 122374 152396 122380 152408
rect 122432 152396 122438 152448
rect 123938 152396 123944 152448
rect 123996 152436 124002 152448
rect 128814 152436 128820 152448
rect 123996 152408 128820 152436
rect 123996 152396 124002 152408
rect 128814 152396 128820 152408
rect 128872 152396 128878 152448
rect 129826 152396 129832 152448
rect 129884 152436 129890 152448
rect 139118 152436 139124 152448
rect 129884 152408 139124 152436
rect 129884 152396 129890 152408
rect 139118 152396 139124 152408
rect 139176 152396 139182 152448
rect 144822 152396 144828 152448
rect 144880 152436 144886 152448
rect 209130 152436 209136 152448
rect 144880 152408 209136 152436
rect 144880 152396 144886 152408
rect 209130 152396 209136 152408
rect 209188 152396 209194 152448
rect 221918 152396 221924 152448
rect 221976 152436 221982 152448
rect 244366 152436 244372 152448
rect 221976 152408 244372 152436
rect 221976 152396 221982 152408
rect 244366 152396 244372 152408
rect 244424 152396 244430 152448
rect 245654 152396 245660 152448
rect 245712 152436 245718 152448
rect 288066 152436 288072 152448
rect 245712 152408 288072 152436
rect 245712 152396 245718 152408
rect 288066 152396 288072 152408
rect 288124 152396 288130 152448
rect 289906 152396 289912 152448
rect 289964 152436 289970 152448
rect 334342 152436 334348 152448
rect 289964 152408 334348 152436
rect 289964 152396 289970 152408
rect 334342 152396 334348 152408
rect 334400 152396 334406 152448
rect 349430 152396 349436 152448
rect 349488 152436 349494 152448
rect 354646 152436 354674 152476
rect 385586 152464 385592 152476
rect 385644 152464 385650 152516
rect 392302 152464 392308 152516
rect 392360 152504 392366 152516
rect 418430 152504 418436 152516
rect 392360 152476 418436 152504
rect 392360 152464 392366 152476
rect 418430 152464 418436 152476
rect 418488 152464 418494 152516
rect 437382 152464 437388 152516
rect 437440 152504 437446 152516
rect 452470 152504 452476 152516
rect 437440 152476 452476 152504
rect 437440 152464 437446 152476
rect 452470 152464 452476 152476
rect 452528 152464 452534 152516
rect 349488 152408 354674 152436
rect 349488 152396 349494 152408
rect 414290 152396 414296 152448
rect 414348 152436 414354 152448
rect 415854 152436 415860 152448
rect 414348 152408 415860 152436
rect 414348 152396 414354 152408
rect 415854 152396 415860 152408
rect 415912 152396 415918 152448
rect 118694 152328 118700 152380
rect 118752 152368 118758 152380
rect 167362 152368 167368 152380
rect 118752 152340 167368 152368
rect 118752 152328 118758 152340
rect 167362 152328 167368 152340
rect 167420 152328 167426 152380
rect 183278 152328 183284 152380
rect 183336 152368 183342 152380
rect 236730 152368 236736 152380
rect 183336 152340 236736 152368
rect 183336 152328 183342 152340
rect 236730 152328 236736 152340
rect 236788 152328 236794 152380
rect 247218 152328 247224 152380
rect 247276 152368 247282 152380
rect 259822 152368 259828 152380
rect 247276 152340 259828 152368
rect 247276 152328 247282 152340
rect 259822 152328 259828 152340
rect 259880 152328 259886 152380
rect 268930 152328 268936 152380
rect 268988 152368 268994 152380
rect 280338 152368 280344 152380
rect 268988 152340 280344 152368
rect 268988 152328 268994 152340
rect 280338 152328 280344 152340
rect 280396 152328 280402 152380
rect 288342 152328 288348 152380
rect 288400 152368 288406 152380
rect 300946 152368 300952 152380
rect 288400 152340 300952 152368
rect 288400 152328 288406 152340
rect 300946 152328 300952 152340
rect 301004 152328 301010 152380
rect 511626 152328 511632 152380
rect 511684 152368 511690 152380
rect 513558 152368 513564 152380
rect 511684 152340 513564 152368
rect 511684 152328 511690 152340
rect 513558 152328 513564 152340
rect 513616 152328 513622 152380
rect 173986 152260 173992 152312
rect 174044 152300 174050 152312
rect 226426 152300 226432 152312
rect 174044 152272 226432 152300
rect 174044 152260 174050 152272
rect 226426 152260 226432 152272
rect 226484 152260 226490 152312
rect 230658 152260 230664 152312
rect 230716 152300 230722 152312
rect 257246 152300 257252 152312
rect 230716 152272 257252 152300
rect 230716 152260 230722 152272
rect 257246 152260 257252 152272
rect 257304 152260 257310 152312
rect 257338 152260 257344 152312
rect 257396 152300 257402 152312
rect 264974 152300 264980 152312
rect 257396 152272 264980 152300
rect 257396 152260 257402 152272
rect 264974 152260 264980 152272
rect 265032 152260 265038 152312
rect 265066 152260 265072 152312
rect 265124 152300 265130 152312
rect 275094 152300 275100 152312
rect 265124 152272 275100 152300
rect 265124 152260 265130 152272
rect 275094 152260 275100 152272
rect 275152 152260 275158 152312
rect 281442 152260 281448 152312
rect 281500 152300 281506 152312
rect 290642 152300 290648 152312
rect 281500 152272 290648 152300
rect 281500 152260 281506 152272
rect 290642 152260 290648 152272
rect 290700 152260 290706 152312
rect 146110 152192 146116 152244
rect 146168 152232 146174 152244
rect 179598 152232 179604 152244
rect 146168 152204 179604 152232
rect 146168 152192 146174 152204
rect 179598 152192 179604 152204
rect 179656 152192 179662 152244
rect 197354 152192 197360 152244
rect 197412 152232 197418 152244
rect 221918 152232 221924 152244
rect 197412 152204 221924 152232
rect 197412 152192 197418 152204
rect 221918 152192 221924 152204
rect 221976 152192 221982 152244
rect 230382 152192 230388 152244
rect 230440 152232 230446 152244
rect 249518 152232 249524 152244
rect 230440 152204 249524 152232
rect 230440 152192 230446 152204
rect 249518 152192 249524 152204
rect 249576 152192 249582 152244
rect 513558 152192 513564 152244
rect 513616 152232 513622 152244
rect 516134 152232 516140 152244
rect 513616 152204 516140 152232
rect 513616 152192 513622 152204
rect 516134 152192 516140 152204
rect 516192 152192 516198 152244
rect 26694 152124 26700 152176
rect 26752 152164 26758 152176
rect 110138 152164 110144 152176
rect 26752 152136 110144 152164
rect 26752 152124 26758 152136
rect 110138 152124 110144 152136
rect 110196 152124 110202 152176
rect 197446 152124 197452 152176
rect 197504 152164 197510 152176
rect 216766 152164 216772 152176
rect 197504 152136 216772 152164
rect 197504 152124 197510 152136
rect 216766 152124 216772 152136
rect 216824 152124 216830 152176
rect 241698 152124 241704 152176
rect 241756 152164 241762 152176
rect 254670 152164 254676 152176
rect 241756 152136 254676 152164
rect 241756 152124 241762 152136
rect 254670 152124 254676 152136
rect 254728 152124 254734 152176
rect 516686 152124 516692 152176
rect 516744 152164 516750 152176
rect 520274 152164 520280 152176
rect 516744 152136 520280 152164
rect 516744 152124 516750 152136
rect 520274 152124 520280 152136
rect 520332 152124 520338 152176
rect 102318 152056 102324 152108
rect 102376 152096 102382 152108
rect 109954 152096 109960 152108
rect 102376 152068 109960 152096
rect 102376 152056 102382 152068
rect 109954 152056 109960 152068
rect 110012 152056 110018 152108
rect 515490 152056 515496 152108
rect 515548 152096 515554 152108
rect 518894 152096 518900 152108
rect 515548 152068 518900 152096
rect 515548 152056 515554 152068
rect 518894 152056 518900 152068
rect 518952 152056 518958 152108
rect 40494 151988 40500 152040
rect 40552 152028 40558 152040
rect 89162 152028 89168 152040
rect 40552 152000 89168 152028
rect 40552 151988 40558 152000
rect 89162 151988 89168 152000
rect 89220 151988 89226 152040
rect 95510 151988 95516 152040
rect 95568 152028 95574 152040
rect 114370 152028 114376 152040
rect 95568 152000 114376 152028
rect 95568 151988 95574 152000
rect 114370 151988 114376 152000
rect 114428 151988 114434 152040
rect 467834 151988 467840 152040
rect 467892 152028 467898 152040
rect 471698 152028 471704 152040
rect 467892 152000 471704 152028
rect 467892 151988 467898 152000
rect 471698 151988 471704 152000
rect 471756 151988 471762 152040
rect 488166 151988 488172 152040
rect 488224 152028 488230 152040
rect 491570 152028 491576 152040
rect 488224 152000 491576 152028
rect 488224 151988 488230 152000
rect 491570 151988 491576 152000
rect 491628 151988 491634 152040
rect 515950 151988 515956 152040
rect 516008 152028 516014 152040
rect 519446 152028 519452 152040
rect 516008 152000 519452 152028
rect 516008 151988 516014 152000
rect 519446 151988 519452 152000
rect 519504 151988 519510 152040
rect 88610 151920 88616 151972
rect 88668 151960 88674 151972
rect 110322 151960 110328 151972
rect 88668 151932 110328 151960
rect 88668 151920 88674 151932
rect 110322 151920 110328 151932
rect 110380 151920 110386 151972
rect 136358 151920 136364 151972
rect 136416 151960 136422 151972
rect 144270 151960 144276 151972
rect 136416 151932 144276 151960
rect 136416 151920 136422 151932
rect 144270 151920 144276 151932
rect 144328 151920 144334 151972
rect 469214 151920 469220 151972
rect 469272 151960 469278 151972
rect 472342 151960 472348 151972
rect 469272 151932 472348 151960
rect 469272 151920 469278 151932
rect 472342 151920 472348 151932
rect 472400 151920 472406 151972
rect 487338 151920 487344 151972
rect 487396 151960 487402 151972
rect 490926 151960 490932 151972
rect 487396 151932 490932 151960
rect 487396 151920 487402 151932
rect 490926 151920 490932 151932
rect 490984 151920 490990 151972
rect 507670 151920 507676 151972
rect 507728 151960 507734 151972
rect 509234 151960 509240 151972
rect 507728 151932 509240 151960
rect 507728 151920 507734 151932
rect 509234 151920 509240 151932
rect 509292 151920 509298 151972
rect 517422 151920 517428 151972
rect 517480 151960 517486 151972
rect 521562 151960 521568 151972
rect 517480 151932 521568 151960
rect 517480 151920 517486 151932
rect 521562 151920 521568 151932
rect 521620 151920 521626 151972
rect 33594 151852 33600 151904
rect 33652 151892 33658 151904
rect 110230 151892 110236 151904
rect 33652 151864 110236 151892
rect 33652 151852 33658 151864
rect 110230 151852 110236 151864
rect 110288 151852 110294 151904
rect 127618 151852 127624 151904
rect 127676 151892 127682 151904
rect 133966 151892 133972 151904
rect 127676 151864 133972 151892
rect 127676 151852 127682 151864
rect 133966 151852 133972 151864
rect 134024 151852 134030 151904
rect 139486 151852 139492 151904
rect 139544 151892 139550 151904
rect 142982 151892 142988 151904
rect 139544 151864 142988 151892
rect 139544 151852 139550 151864
rect 142982 151852 142988 151864
rect 143040 151852 143046 151904
rect 235994 151852 236000 151904
rect 236052 151892 236058 151904
rect 240594 151892 240600 151904
rect 236052 151864 240600 151892
rect 236052 151852 236058 151864
rect 240594 151852 240600 151864
rect 240652 151852 240658 151904
rect 320726 151852 320732 151904
rect 320784 151892 320790 151904
rect 326614 151892 326620 151904
rect 320784 151864 326620 151892
rect 320784 151852 320790 151864
rect 326614 151852 326620 151864
rect 326672 151852 326678 151904
rect 332594 151852 332600 151904
rect 332652 151892 332658 151904
rect 336826 151892 336832 151904
rect 332652 151864 336832 151892
rect 332652 151852 332658 151864
rect 336826 151852 336832 151864
rect 336884 151852 336890 151904
rect 343634 151852 343640 151904
rect 343692 151892 343698 151904
rect 347130 151892 347136 151904
rect 343692 151864 347136 151892
rect 343692 151852 343698 151864
rect 347130 151852 347136 151864
rect 347188 151852 347194 151904
rect 359458 151852 359464 151904
rect 359516 151892 359522 151904
rect 364518 151892 364524 151904
rect 359516 151864 364524 151892
rect 359516 151852 359522 151864
rect 364518 151852 364524 151864
rect 364576 151852 364582 151904
rect 456058 151852 456064 151904
rect 456116 151892 456122 151904
rect 462682 151892 462688 151904
rect 456116 151864 462688 151892
rect 456116 151852 456122 151864
rect 462682 151852 462688 151864
rect 462740 151852 462746 151904
rect 464338 151852 464344 151904
rect 464396 151892 464402 151904
rect 467834 151892 467840 151904
rect 464396 151864 467840 151892
rect 464396 151852 464402 151864
rect 467834 151852 467840 151864
rect 467892 151852 467898 151904
rect 467926 151852 467932 151904
rect 467984 151892 467990 151904
rect 471054 151892 471060 151904
rect 467984 151864 471060 151892
rect 467984 151852 467990 151864
rect 471054 151852 471060 151864
rect 471112 151852 471118 151904
rect 486510 151852 486516 151904
rect 486568 151852 486574 151904
rect 489086 151852 489092 151904
rect 489144 151892 489150 151904
rect 492214 151892 492220 151904
rect 489144 151864 492220 151892
rect 489144 151852 489150 151864
rect 492214 151852 492220 151864
rect 492272 151852 492278 151904
rect 499482 151852 499488 151904
rect 499540 151892 499546 151904
rect 499942 151892 499948 151904
rect 499540 151864 499948 151892
rect 499540 151852 499546 151864
rect 499942 151852 499948 151864
rect 500000 151852 500006 151904
rect 81710 151784 81716 151836
rect 81768 151824 81774 151836
rect 97718 151824 97724 151836
rect 81768 151796 97724 151824
rect 81768 151784 81774 151796
rect 97718 151784 97724 151796
rect 97776 151784 97782 151836
rect 105814 151784 105820 151836
rect 105872 151824 105878 151836
rect 106918 151824 106924 151836
rect 105872 151796 106924 151824
rect 105872 151784 105878 151796
rect 106918 151784 106924 151796
rect 106976 151784 106982 151836
rect 208394 151784 208400 151836
rect 208452 151824 208458 151836
rect 210418 151824 210424 151836
rect 208452 151796 210424 151824
rect 208452 151784 208458 151796
rect 210418 151784 210424 151796
rect 210476 151784 210482 151836
rect 486528 151824 486556 151852
rect 490282 151824 490288 151836
rect 486528 151796 490288 151824
rect 490282 151784 490288 151796
rect 490340 151784 490346 151836
rect 509050 151784 509056 151836
rect 509108 151824 509114 151836
rect 510890 151824 510896 151836
rect 509108 151796 510896 151824
rect 509108 151784 509114 151796
rect 510890 151784 510896 151796
rect 510948 151784 510954 151836
rect 132402 151716 132408 151768
rect 132460 151756 132466 151768
rect 219342 151756 219348 151768
rect 132460 151728 219348 151756
rect 132460 151716 132466 151728
rect 219342 151716 219348 151728
rect 219400 151716 219406 151768
rect 122742 151648 122748 151700
rect 122800 151688 122806 151700
rect 211614 151688 211620 151700
rect 122800 151660 211620 151688
rect 122800 151648 122806 151660
rect 211614 151648 211620 151660
rect 211672 151648 211678 151700
rect 111702 151580 111708 151632
rect 111760 151620 111766 151632
rect 203978 151620 203984 151632
rect 111760 151592 203984 151620
rect 111760 151580 111766 151592
rect 203978 151580 203984 151592
rect 204036 151580 204042 151632
rect 104802 151512 104808 151564
rect 104860 151552 104866 151564
rect 198826 151552 198832 151564
rect 104860 151524 198832 151552
rect 104860 151512 104866 151524
rect 198826 151512 198832 151524
rect 198884 151512 198890 151564
rect 212442 151512 212448 151564
rect 212500 151552 212506 151564
rect 280982 151552 280988 151564
rect 212500 151524 280988 151552
rect 212500 151512 212506 151524
rect 280982 151512 280988 151524
rect 281040 151512 281046 151564
rect 97902 151444 97908 151496
rect 97960 151484 97966 151496
rect 193674 151484 193680 151496
rect 97960 151456 193680 151484
rect 97960 151444 97966 151456
rect 193674 151444 193680 151456
rect 193732 151444 193738 151496
rect 202782 151444 202788 151496
rect 202840 151484 202846 151496
rect 273254 151484 273260 151496
rect 202840 151456 273260 151484
rect 202840 151444 202846 151456
rect 273254 151444 273260 151456
rect 273312 151444 273318 151496
rect 92382 151376 92388 151428
rect 92440 151416 92446 151428
rect 188522 151416 188528 151428
rect 92440 151388 188528 151416
rect 92440 151376 92446 151388
rect 188522 151376 188528 151388
rect 188580 151376 188586 151428
rect 195882 151376 195888 151428
rect 195940 151416 195946 151428
rect 268194 151416 268200 151428
rect 195940 151388 268200 151416
rect 195940 151376 195946 151388
rect 268194 151376 268200 151388
rect 268252 151376 268258 151428
rect 78582 151308 78588 151360
rect 78640 151348 78646 151360
rect 178310 151348 178316 151360
rect 78640 151320 178316 151348
rect 78640 151308 78646 151320
rect 178310 151308 178316 151320
rect 178368 151308 178374 151360
rect 180702 151308 180708 151360
rect 180760 151348 180766 151360
rect 256602 151348 256608 151360
rect 180760 151320 256608 151348
rect 180760 151308 180766 151320
rect 256602 151308 256608 151320
rect 256660 151308 256666 151360
rect 64782 151240 64788 151292
rect 64840 151280 64846 151292
rect 64840 151252 167592 151280
rect 64840 151240 64846 151252
rect 57882 151172 57888 151224
rect 57940 151212 57946 151224
rect 162854 151212 162860 151224
rect 57940 151184 162860 151212
rect 57940 151172 57946 151184
rect 162854 151172 162860 151184
rect 162912 151172 162918 151224
rect 167564 151212 167592 151252
rect 167638 151240 167644 151292
rect 167696 151280 167702 151292
rect 245010 151280 245016 151292
rect 167696 151252 245016 151280
rect 167696 151240 167702 151252
rect 245010 151240 245016 151252
rect 245068 151240 245074 151292
rect 168006 151212 168012 151224
rect 167564 151184 168012 151212
rect 168006 151172 168012 151184
rect 168064 151172 168070 151224
rect 168098 151172 168104 151224
rect 168156 151212 168162 151224
rect 246298 151212 246304 151224
rect 168156 151184 246304 151212
rect 168156 151172 168162 151184
rect 246298 151172 246304 151184
rect 246356 151172 246362 151224
rect 50982 151104 50988 151156
rect 51040 151144 51046 151156
rect 157702 151144 157708 151156
rect 51040 151116 157708 151144
rect 51040 151104 51046 151116
rect 157702 151104 157708 151116
rect 157760 151104 157766 151156
rect 158622 151104 158628 151156
rect 158680 151144 158686 151156
rect 239950 151144 239956 151156
rect 158680 151116 239956 151144
rect 158680 151104 158686 151116
rect 239950 151104 239956 151116
rect 240008 151104 240014 151156
rect 38562 151036 38568 151088
rect 38620 151076 38626 151088
rect 147490 151076 147496 151088
rect 38620 151048 147496 151076
rect 38620 151036 38626 151048
rect 147490 151036 147496 151048
rect 147548 151036 147554 151088
rect 151722 151036 151728 151088
rect 151780 151076 151786 151088
rect 234798 151076 234804 151088
rect 151780 151048 234804 151076
rect 151780 151036 151786 151048
rect 234798 151036 234804 151048
rect 234856 151036 234862 151088
rect 146202 150968 146208 151020
rect 146260 151008 146266 151020
rect 229646 151008 229652 151020
rect 146260 150980 229652 151008
rect 146260 150968 146266 150980
rect 229646 150968 229652 150980
rect 229704 150968 229710 151020
rect 153102 150900 153108 150952
rect 153160 150940 153166 150952
rect 235442 150940 235448 150952
rect 153160 150912 235448 150940
rect 153160 150900 153166 150912
rect 235442 150900 235448 150912
rect 235500 150900 235506 150952
rect 166902 150832 166908 150884
rect 166960 150872 166966 150884
rect 168098 150872 168104 150884
rect 166960 150844 168104 150872
rect 166960 150832 166966 150844
rect 168098 150832 168104 150844
rect 168156 150832 168162 150884
rect 98914 150560 98920 150612
rect 98972 150600 98978 150612
rect 114462 150600 114468 150612
rect 98972 150572 114468 150600
rect 98972 150560 98978 150572
rect 114462 150560 114468 150572
rect 114520 150560 114526 150612
rect 92014 150492 92020 150544
rect 92072 150532 92078 150544
rect 114094 150532 114100 150544
rect 92072 150504 114100 150532
rect 92072 150492 92078 150504
rect 114094 150492 114100 150504
rect 114152 150492 114158 150544
rect 85206 150424 85212 150476
rect 85264 150464 85270 150476
rect 116302 150464 116308 150476
rect 85264 150436 116308 150464
rect 85264 150424 85270 150436
rect 116302 150424 116308 150436
rect 116360 150424 116366 150476
rect 127066 150152 127072 150204
rect 127124 150192 127130 150204
rect 128216 150192 128222 150204
rect 127124 150164 128222 150192
rect 127124 150152 127130 150164
rect 128216 150152 128222 150164
rect 128274 150152 128280 150204
rect 132494 150152 132500 150204
rect 132552 150192 132558 150204
rect 133368 150192 133374 150204
rect 132552 150164 133374 150192
rect 132552 150152 132558 150164
rect 133368 150152 133374 150164
rect 133426 150152 133432 150204
rect 139394 150152 139400 150204
rect 139452 150192 139458 150204
rect 140452 150192 140458 150204
rect 139452 150164 140458 150192
rect 139452 150152 139458 150164
rect 140452 150152 140458 150164
rect 140510 150152 140516 150204
rect 145098 150152 145104 150204
rect 145156 150192 145162 150204
rect 146248 150192 146254 150204
rect 145156 150164 146254 150192
rect 145156 150152 145162 150164
rect 146248 150152 146254 150164
rect 146306 150152 146312 150204
rect 147674 150152 147680 150204
rect 147732 150192 147738 150204
rect 148824 150192 148830 150204
rect 147732 150164 148830 150192
rect 147732 150152 147738 150164
rect 148824 150152 148830 150164
rect 148882 150152 148888 150204
rect 149146 150152 149152 150204
rect 149204 150192 149210 150204
rect 150020 150192 150026 150204
rect 149204 150164 150026 150192
rect 149204 150152 149210 150164
rect 150020 150152 150026 150164
rect 150078 150152 150084 150204
rect 150526 150152 150532 150204
rect 150584 150192 150590 150204
rect 151308 150192 151314 150204
rect 150584 150164 151314 150192
rect 150584 150152 150590 150164
rect 151308 150152 151314 150164
rect 151366 150152 151372 150204
rect 154666 150152 154672 150204
rect 154724 150192 154730 150204
rect 155816 150192 155822 150204
rect 154724 150164 155822 150192
rect 154724 150152 154730 150164
rect 155816 150152 155822 150164
rect 155874 150152 155880 150204
rect 160094 150152 160100 150204
rect 160152 150192 160158 150204
rect 160968 150192 160974 150204
rect 160152 150164 160974 150192
rect 160152 150152 160158 150164
rect 160968 150152 160974 150164
rect 161026 150152 161032 150204
rect 161474 150152 161480 150204
rect 161532 150192 161538 150204
rect 162256 150192 162262 150204
rect 161532 150164 162262 150192
rect 161532 150152 161538 150164
rect 162256 150152 162262 150164
rect 162314 150152 162320 150204
rect 163038 150152 163044 150204
rect 163096 150192 163102 150204
rect 164188 150192 164194 150204
rect 163096 150164 164194 150192
rect 163096 150152 163102 150164
rect 164188 150152 164194 150164
rect 164246 150152 164252 150204
rect 168374 150152 168380 150204
rect 168432 150192 168438 150204
rect 169340 150192 169346 150204
rect 168432 150164 169346 150192
rect 168432 150152 168438 150164
rect 169340 150152 169346 150164
rect 169398 150152 169404 150204
rect 169754 150152 169760 150204
rect 169812 150192 169818 150204
rect 170628 150192 170634 150204
rect 169812 150164 170634 150192
rect 169812 150152 169818 150164
rect 170628 150152 170634 150164
rect 170686 150152 170692 150204
rect 171134 150152 171140 150204
rect 171192 150192 171198 150204
rect 171916 150192 171922 150204
rect 171192 150164 171922 150192
rect 171192 150152 171198 150164
rect 171916 150152 171922 150164
rect 171974 150152 171980 150204
rect 172698 150152 172704 150204
rect 172756 150192 172762 150204
rect 173848 150192 173854 150204
rect 172756 150164 173854 150192
rect 172756 150152 172762 150164
rect 173848 150152 173854 150164
rect 173906 150152 173912 150204
rect 180978 150152 180984 150204
rect 181036 150192 181042 150204
rect 182128 150192 182134 150204
rect 181036 150164 182134 150192
rect 181036 150152 181042 150164
rect 182128 150152 182134 150164
rect 182186 150152 182192 150204
rect 183554 150152 183560 150204
rect 183612 150192 183618 150204
rect 184704 150192 184710 150204
rect 183612 150164 184710 150192
rect 183612 150152 183618 150164
rect 184704 150152 184710 150164
rect 184762 150152 184768 150204
rect 190730 150152 190736 150204
rect 190788 150192 190794 150204
rect 191788 150192 191794 150204
rect 190788 150164 191794 150192
rect 190788 150152 190794 150164
rect 191788 150152 191794 150164
rect 191846 150152 191852 150204
rect 200298 150152 200304 150204
rect 200356 150192 200362 150204
rect 201448 150192 201454 150204
rect 200356 150164 201454 150192
rect 200356 150152 200362 150164
rect 201448 150152 201454 150164
rect 201506 150152 201512 150204
rect 201586 150152 201592 150204
rect 201644 150192 201650 150204
rect 202736 150192 202742 150204
rect 201644 150164 202742 150192
rect 201644 150152 201650 150164
rect 202736 150152 202742 150164
rect 202794 150152 202800 150204
rect 207014 150152 207020 150204
rect 207072 150192 207078 150204
rect 207888 150192 207894 150204
rect 207072 150164 207894 150192
rect 207072 150152 207078 150164
rect 207888 150152 207894 150164
rect 207946 150152 207952 150204
rect 209958 150152 209964 150204
rect 210016 150192 210022 150204
rect 211108 150192 211114 150204
rect 210016 150164 211114 150192
rect 210016 150152 210022 150164
rect 211108 150152 211114 150164
rect 211166 150152 211172 150204
rect 215386 150152 215392 150204
rect 215444 150192 215450 150204
rect 216168 150192 216174 150204
rect 215444 150164 216174 150192
rect 215444 150152 215450 150164
rect 216168 150152 216174 150164
rect 216226 150152 216232 150204
rect 224954 150152 224960 150204
rect 225012 150192 225018 150204
rect 225828 150192 225834 150204
rect 225012 150164 225834 150192
rect 225012 150152 225018 150164
rect 225828 150152 225834 150164
rect 225886 150152 225892 150204
rect 229186 150152 229192 150204
rect 229244 150192 229250 150204
rect 230336 150192 230342 150204
rect 229244 150164 230342 150192
rect 229244 150152 229250 150164
rect 230336 150152 230342 150164
rect 230394 150152 230400 150204
rect 231946 150152 231952 150204
rect 232004 150192 232010 150204
rect 232912 150192 232918 150204
rect 232004 150164 232918 150192
rect 232004 150152 232010 150164
rect 232912 150152 232918 150164
rect 232970 150152 232976 150204
rect 233234 150152 233240 150204
rect 233292 150192 233298 150204
rect 234200 150192 234206 150204
rect 233292 150164 234206 150192
rect 233292 150152 233298 150164
rect 234200 150152 234206 150164
rect 234258 150152 234264 150204
rect 242894 150152 242900 150204
rect 242952 150192 242958 150204
rect 243768 150192 243774 150204
rect 242952 150164 243774 150192
rect 242952 150152 242958 150164
rect 243768 150152 243774 150164
rect 243826 150152 243832 150204
rect 247126 150152 247132 150204
rect 247184 150192 247190 150204
rect 248276 150192 248282 150204
rect 247184 150164 248282 150192
rect 247184 150152 247190 150164
rect 248276 150152 248282 150164
rect 248334 150152 248340 150204
rect 252554 150152 252560 150204
rect 252612 150192 252618 150204
rect 253428 150192 253434 150204
rect 252612 150164 253434 150192
rect 252612 150152 252618 150164
rect 253428 150152 253434 150164
rect 253486 150152 253492 150204
rect 258074 150152 258080 150204
rect 258132 150192 258138 150204
rect 259224 150192 259230 150204
rect 258132 150164 259230 150192
rect 258132 150152 258138 150164
rect 259224 150152 259230 150164
rect 259282 150152 259288 150204
rect 260834 150152 260840 150204
rect 260892 150192 260898 150204
rect 261800 150192 261806 150204
rect 260892 150164 261806 150192
rect 260892 150152 260898 150164
rect 261800 150152 261806 150164
rect 261858 150152 261864 150204
rect 263594 150152 263600 150204
rect 263652 150192 263658 150204
rect 264376 150192 264382 150204
rect 263652 150164 264382 150192
rect 263652 150152 263658 150164
rect 264376 150152 264382 150164
rect 264434 150152 264440 150204
rect 265158 150152 265164 150204
rect 265216 150192 265222 150204
rect 266308 150192 266314 150204
rect 265216 150164 266314 150192
rect 265216 150152 265222 150164
rect 266308 150152 266314 150164
rect 266366 150152 266372 150204
rect 273438 150152 273444 150204
rect 273496 150192 273502 150204
rect 274588 150192 274594 150204
rect 273496 150164 274594 150192
rect 273496 150152 273502 150164
rect 274588 150152 274594 150164
rect 274646 150152 274652 150204
rect 276014 150152 276020 150204
rect 276072 150192 276078 150204
rect 277164 150192 277170 150204
rect 276072 150164 277170 150192
rect 276072 150152 276078 150164
rect 277164 150152 277170 150164
rect 277222 150152 277228 150204
rect 278774 150152 278780 150204
rect 278832 150192 278838 150204
rect 279740 150192 279746 150204
rect 278832 150164 279746 150192
rect 278832 150152 278838 150164
rect 279740 150152 279746 150164
rect 279798 150152 279804 150204
rect 283098 150152 283104 150204
rect 283156 150192 283162 150204
rect 284248 150192 284254 150204
rect 283156 150164 284254 150192
rect 283156 150152 283162 150164
rect 284248 150152 284254 150164
rect 284306 150152 284312 150204
rect 291194 150152 291200 150204
rect 291252 150192 291258 150204
rect 291976 150192 291982 150204
rect 291252 150164 291982 150192
rect 291252 150152 291258 150164
rect 291976 150152 291982 150164
rect 292034 150152 292040 150204
rect 292758 150152 292764 150204
rect 292816 150192 292822 150204
rect 293908 150192 293914 150204
rect 292816 150164 293914 150192
rect 292816 150152 292822 150164
rect 293908 150152 293914 150164
rect 293966 150152 293972 150204
rect 294046 150152 294052 150204
rect 294104 150192 294110 150204
rect 295196 150192 295202 150204
rect 294104 150164 295202 150192
rect 294104 150152 294110 150164
rect 295196 150152 295202 150164
rect 295254 150152 295260 150204
rect 310606 150152 310612 150204
rect 310664 150192 310670 150204
rect 311848 150192 311854 150204
rect 310664 150164 311854 150192
rect 310664 150152 310670 150164
rect 311848 150152 311854 150164
rect 311906 150152 311912 150204
rect 311986 150152 311992 150204
rect 312044 150192 312050 150204
rect 313136 150192 313142 150204
rect 312044 150164 313142 150192
rect 312044 150152 312050 150164
rect 313136 150152 313142 150164
rect 313194 150152 313200 150204
rect 331306 150152 331312 150204
rect 331364 150192 331370 150204
rect 332456 150192 332462 150204
rect 331364 150164 332462 150192
rect 331364 150152 331370 150164
rect 332456 150152 332462 150164
rect 332514 150152 332520 150204
rect 339586 150152 339592 150204
rect 339644 150192 339650 150204
rect 340736 150192 340742 150204
rect 339644 150164 340742 150192
rect 339644 150152 339650 150164
rect 340736 150152 340742 150164
rect 340794 150152 340800 150204
rect 349246 150152 349252 150204
rect 349304 150192 349310 150204
rect 350396 150192 350402 150204
rect 349304 150164 350402 150192
rect 349304 150152 349310 150164
rect 350396 150152 350402 150164
rect 350454 150152 350460 150204
rect 350534 150152 350540 150204
rect 350592 150192 350598 150204
rect 351684 150192 351690 150204
rect 350592 150164 351690 150192
rect 350592 150152 350598 150164
rect 351684 150152 351690 150164
rect 351742 150152 351748 150204
rect 351914 150152 351920 150204
rect 351972 150192 351978 150204
rect 352972 150192 352978 150204
rect 351972 150164 352978 150192
rect 351972 150152 351978 150164
rect 352972 150152 352978 150164
rect 353030 150152 353036 150204
rect 357618 150152 357624 150204
rect 357676 150192 357682 150204
rect 358768 150192 358774 150204
rect 357676 150164 358774 150192
rect 357676 150152 357682 150164
rect 358768 150152 358774 150164
rect 358826 150152 358832 150204
rect 360194 150152 360200 150204
rect 360252 150192 360258 150204
rect 361344 150192 361350 150204
rect 360252 150164 361350 150192
rect 360252 150152 360258 150164
rect 361344 150152 361350 150164
rect 361402 150152 361408 150204
rect 361574 150152 361580 150204
rect 361632 150192 361638 150204
rect 362632 150192 362638 150204
rect 361632 150164 362638 150192
rect 361632 150152 361638 150164
rect 362632 150152 362638 150164
rect 362690 150152 362696 150204
rect 365898 150152 365904 150204
rect 365956 150192 365962 150204
rect 367048 150192 367054 150204
rect 365956 150164 367054 150192
rect 365956 150152 365962 150164
rect 367048 150152 367054 150164
rect 367106 150152 367112 150204
rect 380894 150152 380900 150204
rect 380952 150192 380958 150204
rect 381860 150192 381866 150204
rect 380952 150164 381866 150192
rect 380952 150152 380958 150164
rect 381860 150152 381866 150164
rect 381918 150152 381924 150204
rect 382274 150152 382280 150204
rect 382332 150192 382338 150204
rect 383148 150192 383154 150204
rect 382332 150164 383154 150192
rect 382332 150152 382338 150164
rect 383148 150152 383154 150164
rect 383206 150152 383212 150204
rect 385218 150152 385224 150204
rect 385276 150192 385282 150204
rect 386368 150192 386374 150204
rect 385276 150164 386374 150192
rect 385276 150152 385282 150164
rect 386368 150152 386374 150164
rect 386426 150152 386432 150204
rect 386506 150152 386512 150204
rect 386564 150192 386570 150204
rect 387656 150192 387662 150204
rect 386564 150164 387662 150192
rect 386564 150152 386570 150164
rect 387656 150152 387662 150164
rect 387714 150152 387720 150204
rect 391934 150152 391940 150204
rect 391992 150192 391998 150204
rect 392808 150192 392814 150204
rect 391992 150164 392814 150192
rect 391992 150152 391998 150164
rect 392808 150152 392814 150164
rect 392866 150152 392872 150204
rect 396166 150152 396172 150204
rect 396224 150192 396230 150204
rect 397224 150192 397230 150204
rect 396224 150164 397230 150192
rect 396224 150152 396230 150164
rect 397224 150152 397230 150164
rect 397282 150152 397288 150204
rect 400214 150152 400220 150204
rect 400272 150192 400278 150204
rect 401088 150192 401094 150204
rect 400272 150164 401094 150192
rect 400272 150152 400278 150164
rect 401088 150152 401094 150164
rect 401146 150152 401152 150204
rect 412818 150152 412824 150204
rect 412876 150192 412882 150204
rect 413968 150192 413974 150204
rect 412876 150164 413974 150192
rect 412876 150152 412882 150164
rect 413968 150152 413974 150164
rect 414026 150152 414032 150204
rect 423766 150152 423772 150204
rect 423824 150192 423830 150204
rect 424916 150192 424922 150204
rect 423824 150164 424922 150192
rect 423824 150152 423830 150164
rect 424916 150152 424922 150164
rect 424974 150152 424980 150204
rect 434714 150152 434720 150204
rect 434772 150192 434778 150204
rect 435772 150192 435778 150204
rect 434772 150164 435778 150192
rect 434772 150152 434778 150164
rect 435772 150152 435778 150164
rect 435830 150152 435836 150204
rect 441706 150152 441712 150204
rect 441764 150192 441770 150204
rect 442856 150192 442862 150204
rect 441764 150164 442862 150192
rect 441764 150152 441770 150164
rect 442856 150152 442862 150164
rect 442914 150152 442920 150204
rect 442994 150152 443000 150204
rect 443052 150192 443058 150204
rect 444144 150192 444150 150204
rect 443052 150164 444150 150192
rect 443052 150152 443058 150164
rect 444144 150152 444150 150164
rect 444202 150152 444208 150204
rect 444374 150152 444380 150204
rect 444432 150192 444438 150204
rect 445432 150192 445438 150204
rect 444432 150164 445438 150192
rect 444432 150152 444438 150164
rect 445432 150152 445438 150164
rect 445490 150152 445496 150204
rect 456794 150152 456800 150204
rect 456852 150192 456858 150204
rect 457668 150192 457674 150204
rect 456852 150164 457674 150192
rect 456852 150152 456858 150164
rect 457668 150152 457674 150164
rect 457726 150152 457732 150204
rect 458358 150152 458364 150204
rect 458416 150192 458422 150204
rect 459508 150192 459514 150204
rect 458416 150164 459514 150192
rect 458416 150152 458422 150164
rect 459508 150152 459514 150164
rect 459566 150152 459572 150204
rect 477678 150152 477684 150204
rect 477736 150192 477742 150204
rect 478828 150192 478834 150204
rect 477736 150164 478834 150192
rect 477736 150152 477742 150164
rect 478828 150152 478834 150164
rect 478886 150152 478892 150204
rect 478966 150152 478972 150204
rect 479024 150192 479030 150204
rect 480116 150192 480122 150204
rect 479024 150164 480122 150192
rect 479024 150152 479030 150164
rect 480116 150152 480122 150164
rect 480174 150152 480180 150204
rect 480254 150152 480260 150204
rect 480312 150192 480318 150204
rect 481404 150192 481410 150204
rect 480312 150164 481410 150192
rect 480312 150152 480318 150164
rect 481404 150152 481410 150164
rect 481462 150152 481468 150204
rect 481634 150152 481640 150204
rect 481692 150192 481698 150204
rect 482692 150192 482698 150204
rect 481692 150164 482698 150192
rect 481692 150152 481698 150164
rect 482692 150152 482698 150164
rect 482750 150152 482756 150204
rect 97718 149880 97724 149932
rect 97776 149920 97782 149932
rect 117222 149920 117228 149932
rect 97776 149892 117228 149920
rect 97776 149880 97782 149892
rect 117222 149880 117228 149892
rect 117280 149880 117286 149932
rect 89162 149812 89168 149864
rect 89220 149852 89226 149864
rect 117130 149852 117136 149864
rect 89220 149824 117136 149852
rect 89220 149812 89226 149824
rect 117130 149812 117136 149824
rect 117188 149812 117194 149864
rect 78582 149744 78588 149796
rect 78640 149784 78646 149796
rect 112806 149784 112812 149796
rect 78640 149756 112812 149784
rect 78640 149744 78646 149756
rect 112806 149744 112812 149756
rect 112864 149744 112870 149796
rect 71682 149676 71688 149728
rect 71740 149716 71746 149728
rect 109678 149716 109684 149728
rect 71740 149688 109684 149716
rect 71740 149676 71746 149688
rect 109678 149676 109684 149688
rect 109736 149676 109742 149728
rect 75178 149608 75184 149660
rect 75236 149648 75242 149660
rect 114278 149648 114284 149660
rect 75236 149620 114284 149648
rect 75236 149608 75242 149620
rect 114278 149608 114284 149620
rect 114336 149608 114342 149660
rect 68370 149540 68376 149592
rect 68428 149580 68434 149592
rect 112714 149580 112720 149592
rect 68428 149552 112720 149580
rect 68428 149540 68434 149552
rect 112714 149540 112720 149552
rect 112772 149540 112778 149592
rect 64690 149472 64696 149524
rect 64748 149512 64754 149524
rect 111334 149512 111340 149524
rect 64748 149484 111340 149512
rect 64748 149472 64754 149484
rect 111334 149472 111340 149484
rect 111392 149472 111398 149524
rect 61378 149404 61384 149456
rect 61436 149444 61442 149456
rect 112622 149444 112628 149456
rect 61436 149416 112628 149444
rect 61436 149404 61442 149416
rect 112622 149404 112628 149416
rect 112680 149404 112686 149456
rect 57882 149336 57888 149388
rect 57940 149376 57946 149388
rect 112530 149376 112536 149388
rect 57940 149348 112536 149376
rect 57940 149336 57946 149348
rect 112530 149336 112536 149348
rect 112588 149336 112594 149388
rect 44082 149268 44088 149320
rect 44140 149308 44146 149320
rect 44140 149280 45554 149308
rect 44140 149268 44146 149280
rect 45526 149104 45554 149280
rect 47578 149268 47584 149320
rect 47636 149268 47642 149320
rect 50982 149268 50988 149320
rect 51040 149268 51046 149320
rect 54570 149268 54576 149320
rect 54628 149308 54634 149320
rect 111242 149308 111248 149320
rect 54628 149280 111248 149308
rect 54628 149268 54634 149280
rect 111242 149268 111248 149280
rect 111300 149268 111306 149320
rect 47596 149172 47624 149268
rect 51000 149240 51028 149268
rect 112438 149240 112444 149252
rect 51000 149212 112444 149240
rect 112438 149200 112444 149212
rect 112496 149200 112502 149252
rect 111150 149172 111156 149184
rect 47596 149144 111156 149172
rect 111150 149132 111156 149144
rect 111208 149132 111214 149184
rect 111058 149104 111064 149116
rect 45526 149076 111064 149104
rect 111058 149064 111064 149076
rect 111116 149064 111122 149116
rect 109586 148996 109592 149048
rect 109644 149036 109650 149048
rect 116118 149036 116124 149048
rect 109644 149008 116124 149036
rect 109644 148996 109650 149008
rect 116118 148996 116124 149008
rect 116176 148996 116182 149048
rect 111794 147568 111800 147620
rect 111852 147608 111858 147620
rect 116118 147608 116124 147620
rect 111852 147580 116124 147608
rect 111852 147568 111858 147580
rect 116118 147568 116124 147580
rect 116176 147568 116182 147620
rect 109954 147092 109960 147144
rect 110012 147132 110018 147144
rect 116026 147132 116032 147144
rect 110012 147104 116032 147132
rect 110012 147092 110018 147104
rect 116026 147092 116032 147104
rect 116084 147092 116090 147144
rect 110322 147024 110328 147076
rect 110380 147064 110386 147076
rect 116394 147064 116400 147076
rect 110380 147036 116400 147064
rect 110380 147024 110386 147036
rect 116394 147024 116400 147036
rect 116452 147024 116458 147076
rect 110046 146956 110052 147008
rect 110104 146996 110110 147008
rect 116762 146996 116768 147008
rect 110104 146968 116768 146996
rect 110104 146956 110110 146968
rect 116762 146956 116768 146968
rect 116820 146956 116826 147008
rect 110138 146888 110144 146940
rect 110196 146928 110202 146940
rect 116854 146928 116860 146940
rect 110196 146900 116860 146928
rect 110196 146888 110202 146900
rect 116854 146888 116860 146900
rect 116912 146888 116918 146940
rect 110230 145528 110236 145580
rect 110288 145568 110294 145580
rect 117038 145568 117044 145580
rect 110288 145540 117044 145568
rect 110288 145528 110294 145540
rect 117038 145528 117044 145540
rect 117096 145528 117102 145580
rect 113726 143556 113732 143608
rect 113784 143596 113790 143608
rect 115198 143596 115204 143608
rect 113784 143568 115204 143596
rect 113784 143556 113790 143568
rect 115198 143556 115204 143568
rect 115256 143556 115262 143608
rect 114462 143488 114468 143540
rect 114520 143528 114526 143540
rect 116118 143528 116124 143540
rect 114520 143500 116124 143528
rect 114520 143488 114526 143500
rect 116118 143488 116124 143500
rect 116176 143488 116182 143540
rect 114370 141720 114376 141772
rect 114428 141760 114434 141772
rect 116486 141760 116492 141772
rect 114428 141732 116492 141760
rect 114428 141720 114434 141732
rect 116486 141720 116492 141732
rect 116544 141720 116550 141772
rect 114094 140700 114100 140752
rect 114152 140740 114158 140752
rect 116486 140740 116492 140752
rect 114152 140712 116492 140740
rect 114152 140700 114158 140712
rect 116486 140700 116492 140712
rect 116544 140700 116550 140752
rect 112806 132404 112812 132456
rect 112864 132444 112870 132456
rect 116118 132444 116124 132456
rect 112864 132416 116124 132444
rect 112864 132404 112870 132416
rect 116118 132404 116124 132416
rect 116176 132404 116182 132456
rect 114278 131044 114284 131096
rect 114336 131084 114342 131096
rect 115934 131084 115940 131096
rect 114336 131056 115940 131084
rect 114336 131044 114342 131056
rect 115934 131044 115940 131056
rect 115992 131044 115998 131096
rect 109678 128256 109684 128308
rect 109736 128296 109742 128308
rect 116118 128296 116124 128308
rect 109736 128268 116124 128296
rect 109736 128256 109742 128268
rect 116118 128256 116124 128268
rect 116176 128256 116182 128308
rect 112714 126896 112720 126948
rect 112772 126936 112778 126948
rect 116118 126936 116124 126948
rect 112772 126908 116124 126936
rect 112772 126896 112778 126908
rect 116118 126896 116124 126908
rect 116176 126896 116182 126948
rect 111334 124108 111340 124160
rect 111392 124148 111398 124160
rect 116118 124148 116124 124160
rect 111392 124120 116124 124148
rect 111392 124108 111398 124120
rect 116118 124108 116124 124120
rect 116176 124108 116182 124160
rect 112622 122748 112628 122800
rect 112680 122788 112686 122800
rect 115934 122788 115940 122800
rect 112680 122760 115940 122788
rect 112680 122748 112686 122760
rect 115934 122748 115940 122760
rect 115992 122748 115998 122800
rect 112530 121388 112536 121440
rect 112588 121428 112594 121440
rect 116118 121428 116124 121440
rect 112588 121400 116124 121428
rect 112588 121388 112594 121400
rect 116118 121388 116124 121400
rect 116176 121388 116182 121440
rect 114278 118736 114284 118788
rect 114336 118776 114342 118788
rect 115290 118776 115296 118788
rect 114336 118748 115296 118776
rect 114336 118736 114342 118748
rect 115290 118736 115296 118748
rect 115348 118736 115354 118788
rect 111242 118600 111248 118652
rect 111300 118640 111306 118652
rect 116118 118640 116124 118652
rect 111300 118612 116124 118640
rect 111300 118600 111306 118612
rect 116118 118600 116124 118612
rect 116176 118600 116182 118652
rect 112438 117240 112444 117292
rect 112496 117280 112502 117292
rect 116118 117280 116124 117292
rect 112496 117252 116124 117280
rect 112496 117240 112502 117252
rect 116118 117240 116124 117252
rect 116176 117240 116182 117292
rect 111150 114452 111156 114504
rect 111208 114492 111214 114504
rect 116118 114492 116124 114504
rect 111208 114464 116124 114492
rect 111208 114452 111214 114464
rect 116118 114452 116124 114464
rect 116176 114452 116182 114504
rect 111058 113092 111064 113144
rect 111116 113132 111122 113144
rect 116118 113132 116124 113144
rect 111116 113104 116124 113132
rect 111116 113092 111122 113104
rect 116118 113092 116124 113104
rect 116176 113092 116182 113144
rect 113542 109624 113548 109676
rect 113600 109664 113606 109676
rect 115382 109664 115388 109676
rect 113600 109636 115388 109664
rect 113600 109624 113606 109636
rect 115382 109624 115388 109636
rect 115440 109624 115446 109676
rect 114186 104796 114192 104848
rect 114244 104836 114250 104848
rect 115934 104836 115940 104848
rect 114244 104808 115940 104836
rect 114244 104796 114250 104808
rect 115934 104796 115940 104808
rect 115992 104796 115998 104848
rect 114002 99288 114008 99340
rect 114060 99328 114066 99340
rect 116486 99328 116492 99340
rect 114060 99300 116492 99328
rect 114060 99288 114066 99300
rect 116486 99288 116492 99300
rect 116544 99288 116550 99340
rect 114462 96840 114468 96892
rect 114520 96880 114526 96892
rect 116762 96880 116768 96892
rect 114520 96852 116768 96880
rect 114520 96840 114526 96852
rect 116762 96840 116768 96852
rect 116820 96840 116826 96892
rect 113818 93576 113824 93628
rect 113876 93616 113882 93628
rect 116486 93616 116492 93628
rect 113876 93588 116492 93616
rect 113876 93576 113882 93588
rect 116486 93576 116492 93588
rect 116544 93576 116550 93628
rect 113910 92420 113916 92472
rect 113968 92460 113974 92472
rect 116118 92460 116124 92472
rect 113968 92432 116124 92460
rect 113968 92420 113974 92432
rect 116118 92420 116124 92432
rect 116176 92420 116182 92472
rect 115198 91604 115204 91656
rect 115256 91644 115262 91656
rect 116854 91644 116860 91656
rect 115256 91616 116860 91644
rect 115256 91604 115262 91616
rect 116854 91604 116860 91616
rect 116912 91604 116918 91656
rect 114462 87184 114468 87236
rect 114520 87224 114526 87236
rect 116670 87224 116676 87236
rect 114520 87196 116676 87224
rect 114520 87184 114526 87196
rect 116670 87184 116676 87196
rect 116728 87184 116734 87236
rect 114094 86912 114100 86964
rect 114152 86952 114158 86964
rect 116210 86952 116216 86964
rect 114152 86924 116216 86952
rect 114152 86912 114158 86924
rect 116210 86912 116216 86924
rect 116268 86912 116274 86964
rect 113910 71748 113916 71800
rect 113968 71788 113974 71800
rect 116486 71788 116492 71800
rect 113968 71760 116492 71788
rect 113968 71748 113974 71760
rect 116486 71748 116492 71760
rect 116544 71748 116550 71800
rect 114094 69028 114100 69080
rect 114152 69068 114158 69080
rect 116302 69068 116308 69080
rect 114152 69040 116308 69068
rect 114152 69028 114158 69040
rect 116302 69028 116308 69040
rect 116360 69028 116366 69080
rect 114186 67600 114192 67652
rect 114244 67640 114250 67652
rect 116210 67640 116216 67652
rect 114244 67612 116216 67640
rect 114244 67600 114250 67612
rect 116210 67600 116216 67612
rect 116268 67600 116274 67652
rect 113542 64744 113548 64796
rect 113600 64784 113606 64796
rect 116578 64784 116584 64796
rect 113600 64756 116584 64784
rect 113600 64744 113606 64756
rect 116578 64744 116584 64756
rect 116636 64744 116642 64796
rect 112438 62092 112444 62144
rect 112496 62132 112502 62144
rect 116118 62132 116124 62144
rect 112496 62104 116124 62132
rect 112496 62092 112502 62104
rect 116118 62092 116124 62104
rect 116176 62092 116182 62144
rect 113818 52436 113824 52488
rect 113876 52476 113882 52488
rect 116394 52476 116400 52488
rect 113876 52448 116400 52476
rect 113876 52436 113882 52448
rect 116394 52436 116400 52448
rect 116452 52436 116458 52488
rect 113910 48288 113916 48340
rect 113968 48328 113974 48340
rect 115934 48328 115940 48340
rect 113968 48300 115940 48328
rect 113968 48288 113974 48300
rect 115934 48288 115940 48300
rect 115992 48288 115998 48340
rect 111058 46928 111064 46980
rect 111116 46968 111122 46980
rect 116026 46968 116032 46980
rect 111116 46940 116032 46968
rect 111116 46928 111122 46940
rect 116026 46928 116032 46940
rect 116084 46928 116090 46980
rect 113634 44140 113640 44192
rect 113692 44180 113698 44192
rect 117130 44180 117136 44192
rect 113692 44152 117136 44180
rect 113692 44140 113698 44152
rect 117130 44140 117136 44152
rect 117188 44140 117194 44192
rect 114002 41420 114008 41472
rect 114060 41460 114066 41472
rect 115934 41460 115940 41472
rect 114060 41432 115940 41460
rect 114060 41420 114066 41432
rect 115934 41420 115940 41432
rect 115992 41420 115998 41472
rect 114094 38632 114100 38684
rect 114152 38672 114158 38684
rect 115934 38672 115940 38684
rect 114152 38644 115940 38672
rect 114152 38632 114158 38644
rect 115934 38632 115940 38644
rect 115992 38632 115998 38684
rect 114278 37272 114284 37324
rect 114336 37312 114342 37324
rect 116394 37312 116400 37324
rect 114336 37284 116400 37312
rect 114336 37272 114342 37284
rect 116394 37272 116400 37284
rect 116452 37272 116458 37324
rect 114370 34484 114376 34536
rect 114428 34524 114434 34536
rect 115934 34524 115940 34536
rect 114428 34496 115940 34524
rect 114428 34484 114434 34496
rect 115934 34484 115940 34496
rect 115992 34484 115998 34536
rect 113726 33124 113732 33176
rect 113784 33164 113790 33176
rect 116394 33164 116400 33176
rect 113784 33136 116400 33164
rect 113784 33124 113790 33136
rect 116394 33124 116400 33136
rect 116452 33124 116458 33176
rect 114462 31764 114468 31816
rect 114520 31804 114526 31816
rect 115934 31804 115940 31816
rect 114520 31776 115940 31804
rect 114520 31764 114526 31776
rect 115934 31764 115940 31776
rect 115992 31764 115998 31816
rect 111150 28976 111156 29028
rect 111208 29016 111214 29028
rect 116118 29016 116124 29028
rect 111208 28988 116124 29016
rect 111208 28976 111214 28988
rect 116118 28976 116124 28988
rect 116176 28976 116182 29028
rect 111242 27616 111248 27668
rect 111300 27656 111306 27668
rect 116118 27656 116124 27668
rect 111300 27628 116124 27656
rect 111300 27616 111306 27628
rect 116118 27616 116124 27628
rect 116176 27616 116182 27668
rect 112530 24828 112536 24880
rect 112588 24868 112594 24880
rect 116118 24868 116124 24880
rect 112588 24840 116124 24868
rect 112588 24828 112594 24840
rect 116118 24828 116124 24840
rect 116176 24828 116182 24880
rect 114186 22108 114192 22160
rect 114244 22148 114250 22160
rect 115934 22148 115940 22160
rect 114244 22120 115940 22148
rect 114244 22108 114250 22120
rect 115934 22108 115940 22120
rect 115992 22108 115998 22160
rect 111334 19320 111340 19372
rect 111392 19360 111398 19372
rect 116118 19360 116124 19372
rect 111392 19332 116124 19360
rect 111392 19320 111398 19332
rect 116118 19320 116124 19332
rect 116176 19320 116182 19372
rect 113542 13812 113548 13864
rect 113600 13852 113606 13864
rect 116210 13852 116216 13864
rect 113600 13824 116216 13852
rect 113600 13812 113606 13824
rect 116210 13812 116216 13824
rect 116268 13812 116274 13864
rect 113634 8236 113640 8288
rect 113692 8276 113698 8288
rect 115198 8276 115204 8288
rect 113692 8248 115204 8276
rect 113692 8236 113698 8248
rect 115198 8236 115204 8248
rect 115256 8236 115262 8288
rect 109678 4904 109684 4956
rect 109736 4944 109742 4956
rect 116486 4944 116492 4956
rect 109736 4916 116492 4944
rect 109736 4904 109742 4916
rect 116486 4904 116492 4916
rect 116544 4904 116550 4956
rect 109862 4836 109868 4888
rect 109920 4876 109926 4888
rect 116394 4876 116400 4888
rect 109920 4848 116400 4876
rect 109920 4836 109926 4848
rect 116394 4836 116400 4848
rect 116452 4836 116458 4888
rect 109770 4768 109776 4820
rect 109828 4808 109834 4820
rect 117130 4808 117136 4820
rect 109828 4780 117136 4808
rect 109828 4768 109834 4780
rect 117130 4768 117136 4780
rect 117188 4768 117194 4820
rect 109586 4496 109592 4548
rect 109644 4536 109650 4548
rect 112438 4536 112444 4548
rect 109644 4508 112444 4536
rect 109644 4496 109650 4508
rect 112438 4496 112444 4508
rect 112496 4496 112502 4548
rect 109954 4156 109960 4208
rect 110012 4196 110018 4208
rect 116118 4196 116124 4208
rect 110012 4168 116124 4196
rect 110012 4156 110018 4168
rect 116118 4156 116124 4168
rect 116176 4156 116182 4208
rect 110046 2972 110052 2984
rect 84166 2944 110052 2972
rect 84166 2836 84194 2944
rect 110046 2932 110052 2944
rect 110104 2932 110110 2984
rect 110414 2904 110420 2916
rect 32508 2808 84194 2836
rect 98380 2876 110420 2904
rect 32508 2644 32536 2808
rect 32490 2592 32496 2644
rect 32548 2592 32554 2644
rect 98270 2592 98276 2644
rect 98328 2632 98334 2644
rect 98380 2632 98408 2876
rect 110414 2864 110420 2876
rect 110472 2864 110478 2916
rect 98328 2604 98408 2632
rect 98328 2592 98334 2604
rect 106182 2320 106188 2372
rect 106240 2360 106246 2372
rect 116578 2360 116584 2372
rect 106240 2332 116584 2360
rect 106240 2320 106246 2332
rect 116578 2320 116584 2332
rect 116636 2320 116642 2372
rect 102962 2252 102968 2304
rect 103020 2292 103026 2304
rect 116670 2292 116676 2304
rect 103020 2264 116676 2292
rect 103020 2252 103026 2264
rect 116670 2252 116676 2264
rect 116728 2252 116734 2304
rect 99650 2184 99656 2236
rect 99708 2224 99714 2236
rect 116762 2224 116768 2236
rect 99708 2196 116768 2224
rect 99708 2184 99714 2196
rect 116762 2184 116768 2196
rect 116820 2184 116826 2236
rect 96338 2116 96344 2168
rect 96396 2156 96402 2168
rect 116854 2156 116860 2168
rect 96396 2128 116860 2156
rect 96396 2116 96402 2128
rect 116854 2116 116860 2128
rect 116912 2116 116918 2168
rect 89622 2048 89628 2100
rect 89680 2088 89686 2100
rect 116946 2088 116952 2100
rect 89680 2060 116952 2088
rect 89680 2048 89686 2060
rect 116946 2048 116952 2060
rect 117004 2048 117010 2100
rect 82722 1980 82728 2032
rect 82780 2020 82786 2032
rect 111058 2020 111064 2032
rect 82780 1992 111064 2020
rect 82780 1980 82786 1992
rect 111058 1980 111064 1992
rect 111116 1980 111122 2032
rect 76006 1912 76012 1964
rect 76064 1952 76070 1964
rect 109770 1952 109776 1964
rect 76064 1924 109776 1952
rect 76064 1912 76070 1924
rect 109770 1912 109776 1924
rect 109828 1912 109834 1964
rect 62666 1844 62672 1896
rect 62724 1884 62730 1896
rect 114370 1884 114376 1896
rect 62724 1856 114376 1884
rect 62724 1844 62730 1856
rect 114370 1844 114376 1856
rect 114428 1844 114434 1896
rect 491294 1844 491300 1896
rect 491352 1884 491358 1896
rect 493916 1884 493922 1896
rect 491352 1856 493922 1884
rect 491352 1844 491358 1856
rect 493916 1844 493922 1856
rect 493974 1844 493980 1896
rect 59354 1776 59360 1828
rect 59412 1816 59418 1828
rect 113726 1816 113732 1828
rect 59412 1788 113732 1816
rect 59412 1776 59418 1788
rect 113726 1776 113732 1788
rect 113784 1776 113790 1828
rect 49326 1708 49332 1760
rect 49384 1748 49390 1760
rect 111150 1748 111156 1760
rect 49384 1720 111156 1748
rect 49384 1708 49390 1720
rect 111150 1708 111156 1720
rect 111208 1708 111214 1760
rect 46014 1640 46020 1692
rect 46072 1680 46078 1692
rect 111242 1680 111248 1692
rect 46072 1652 111248 1680
rect 46072 1640 46078 1652
rect 111242 1640 111248 1652
rect 111300 1640 111306 1692
rect 35986 1572 35992 1624
rect 36044 1612 36050 1624
rect 114186 1612 114192 1624
rect 36044 1584 114192 1612
rect 36044 1572 36050 1584
rect 114186 1572 114192 1584
rect 114244 1572 114250 1624
rect 39298 1504 39304 1556
rect 39356 1544 39362 1556
rect 117222 1544 117228 1556
rect 39356 1516 117228 1544
rect 39356 1504 39362 1516
rect 117222 1504 117228 1516
rect 117280 1504 117286 1556
rect 15930 1436 15936 1488
rect 15988 1476 15994 1488
rect 98638 1476 98644 1488
rect 15988 1448 98644 1476
rect 15988 1436 15994 1448
rect 98638 1436 98644 1448
rect 98696 1436 98702 1488
rect 110046 1436 110052 1488
rect 110104 1476 110110 1488
rect 143626 1476 143632 1488
rect 110104 1448 143632 1476
rect 110104 1436 110110 1448
rect 143626 1436 143632 1448
rect 143684 1436 143690 1488
rect 12618 1368 12624 1420
rect 12676 1408 12682 1420
rect 100754 1408 100760 1420
rect 12676 1380 100760 1408
rect 12676 1368 12682 1380
rect 100754 1368 100760 1380
rect 100812 1368 100818 1420
rect 110414 1368 110420 1420
rect 110472 1408 110478 1420
rect 193582 1408 193588 1420
rect 110472 1380 193588 1408
rect 110472 1368 110478 1380
rect 193582 1368 193588 1380
rect 193640 1368 193646 1420
rect 92658 1300 92664 1352
rect 92716 1340 92722 1352
rect 113818 1340 113824 1352
rect 92716 1312 113824 1340
rect 92716 1300 92722 1312
rect 113818 1300 113824 1312
rect 113876 1300 113882 1352
rect 22646 1232 22652 1284
rect 22704 1272 22710 1284
rect 113634 1272 113640 1284
rect 22704 1244 113640 1272
rect 22704 1232 22710 1244
rect 113634 1232 113640 1244
rect 113692 1232 113698 1284
rect 42610 1164 42616 1216
rect 42668 1204 42674 1216
rect 112530 1204 112536 1216
rect 42668 1176 112536 1204
rect 42668 1164 42674 1176
rect 112530 1164 112536 1176
rect 112588 1164 112594 1216
rect 52638 1096 52644 1148
rect 52696 1136 52702 1148
rect 114462 1136 114468 1148
rect 52696 1108 114468 1136
rect 52696 1096 52702 1108
rect 114462 1096 114468 1108
rect 114520 1096 114526 1148
rect 65978 1028 65984 1080
rect 66036 1068 66042 1080
rect 114278 1068 114284 1080
rect 66036 1040 114284 1068
rect 66036 1028 66042 1040
rect 114278 1028 114284 1040
rect 114336 1028 114342 1080
rect 69290 960 69296 1012
rect 69348 1000 69354 1012
rect 114094 1000 114100 1012
rect 69348 972 114100 1000
rect 69348 960 69354 972
rect 114094 960 114100 972
rect 114152 960 114158 1012
rect 72694 892 72700 944
rect 72752 932 72758 944
rect 114002 932 114008 944
rect 72752 904 114008 932
rect 72752 892 72758 904
rect 114002 892 114008 904
rect 114060 892 114066 944
rect 79318 824 79324 876
rect 79376 864 79382 876
rect 117038 864 117044 876
rect 79376 836 117044 864
rect 79376 824 79382 836
rect 117038 824 117044 836
rect 117096 824 117102 876
rect 86034 756 86040 808
rect 86092 796 86098 808
rect 113910 796 113916 808
rect 86092 768 113916 796
rect 86092 756 86098 768
rect 113910 756 113916 768
rect 113968 756 113974 808
rect 2682 688 2688 740
rect 2740 728 2746 740
rect 116118 728 116124 740
rect 2740 700 116124 728
rect 2740 688 2746 700
rect 116118 688 116124 700
rect 116176 688 116182 740
<< via1 >>
rect 43260 162596 43312 162648
rect 151912 162596 151964 162648
rect 39856 162528 39908 162580
rect 149428 162528 149480 162580
rect 102140 162460 102192 162512
rect 196900 162460 196952 162512
rect 108856 162392 108908 162444
rect 202052 162392 202104 162444
rect 95424 162324 95476 162376
rect 190736 162324 190788 162376
rect 98736 162256 98788 162308
rect 193404 162256 193456 162308
rect 92020 162188 92072 162240
rect 189172 162188 189224 162240
rect 88708 162120 88760 162172
rect 186320 162120 186372 162172
rect 81900 162052 81952 162104
rect 181076 162052 181128 162104
rect 71872 161984 71924 162036
rect 172704 161984 172756 162036
rect 78588 161916 78640 161968
rect 178224 161916 178276 161968
rect 75184 161848 75236 161900
rect 175556 161848 175608 161900
rect 65156 161780 65208 161832
rect 168472 161780 168524 161832
rect 68468 161712 68520 161764
rect 171324 161712 171376 161764
rect 61752 161644 61804 161696
rect 165620 161644 165672 161696
rect 56692 161576 56744 161628
rect 161480 161576 161532 161628
rect 115572 161508 115624 161560
rect 207204 161508 207256 161560
rect 112260 161440 112312 161492
rect 204260 161440 204312 161492
rect 114744 161372 114796 161424
rect 206192 161372 206244 161424
rect 108028 161304 108080 161356
rect 200304 161304 200356 161356
rect 101312 161236 101364 161288
rect 196256 161236 196308 161288
rect 94596 161168 94648 161220
rect 191104 161168 191156 161220
rect 205548 161168 205600 161220
rect 275192 161168 275244 161220
rect 81072 161100 81124 161152
rect 180892 161100 180944 161152
rect 198832 161100 198884 161152
rect 270500 161100 270552 161152
rect 67640 161032 67692 161084
rect 169760 161032 169812 161084
rect 183744 161032 183796 161084
rect 258080 161032 258132 161084
rect 60924 160964 60976 161016
rect 165436 160964 165488 161016
rect 175280 160964 175332 161016
rect 252744 160964 252796 161016
rect 54208 160896 54260 160948
rect 160376 160896 160428 160948
rect 166080 160896 166132 160948
rect 245752 160896 245804 160948
rect 47492 160828 47544 160880
rect 155040 160828 155092 160880
rect 161848 160828 161900 160880
rect 242072 160828 242124 160880
rect 40684 160760 40736 160812
rect 149152 160760 149204 160812
rect 155132 160760 155184 160812
rect 237380 160760 237432 160812
rect 36544 160692 36596 160744
rect 146852 160692 146904 160744
rect 148416 160692 148468 160744
rect 232228 160692 232280 160744
rect 124864 160624 124916 160676
rect 213920 160624 213972 160676
rect 141700 160556 141752 160608
rect 227076 160556 227128 160608
rect 149244 160488 149296 160540
rect 231952 160488 232004 160540
rect 49976 160012 50028 160064
rect 109224 160012 109276 160064
rect 120632 160012 120684 160064
rect 183284 160012 183336 160064
rect 187884 160012 187936 160064
rect 210148 160012 210200 160064
rect 217324 160012 217376 160064
rect 223488 160012 223540 160064
rect 228272 160012 228324 160064
rect 239956 160012 240008 160064
rect 240876 160012 240928 160064
rect 263876 160012 263928 160064
rect 265348 160012 265400 160064
rect 311072 160012 311124 160064
rect 318340 160012 318392 160064
rect 336648 160012 336700 160064
rect 342720 160012 342772 160064
rect 372620 160012 372672 160064
rect 409144 160012 409196 160064
rect 431224 160012 431276 160064
rect 457076 160012 457128 160064
rect 464344 160012 464396 160064
rect 66812 159944 66864 159996
rect 135628 159944 135680 159996
rect 164332 159944 164384 159996
rect 221924 159944 221976 159996
rect 234160 159944 234212 159996
rect 255504 159944 255556 159996
rect 258540 159944 258592 159996
rect 305000 159944 305052 159996
rect 311532 159944 311584 159996
rect 330208 159944 330260 159996
rect 332600 159944 332652 159996
rect 368480 159944 368532 159996
rect 393136 159944 393188 159996
rect 419080 159944 419132 159996
rect 425980 159944 426032 159996
rect 426440 159944 426492 159996
rect 430212 159944 430264 159996
rect 433064 159944 433116 159996
rect 450360 159944 450412 159996
rect 456064 159944 456116 159996
rect 457904 159944 457956 159996
rect 464712 159944 464764 159996
rect 76932 159876 76984 159928
rect 147772 159876 147824 159928
rect 150900 159876 150952 159928
rect 207020 159876 207072 159928
rect 208952 159876 209004 159928
rect 220176 159876 220228 159928
rect 222384 159876 222436 159928
rect 225696 159876 225748 159928
rect 238392 159876 238444 159928
rect 288348 159876 288400 159928
rect 291384 159876 291436 159928
rect 311900 159876 311952 159928
rect 325884 159876 325936 159928
rect 362132 159876 362184 159928
rect 386420 159876 386472 159928
rect 412824 159876 412876 159928
rect 86960 159808 87012 159860
rect 160284 159808 160336 159860
rect 171140 159808 171192 159860
rect 230388 159808 230440 159860
rect 231676 159808 231728 159860
rect 284392 159808 284444 159860
rect 305644 159808 305696 159860
rect 346308 159808 346360 159860
rect 375472 159808 375524 159860
rect 405556 159808 405608 159860
rect 406660 159808 406712 159860
rect 429384 159808 429436 159860
rect 472256 159808 472308 159860
rect 479432 159808 479484 159860
rect 479800 159808 479852 159860
rect 485228 159808 485280 159860
rect 60096 159740 60148 159792
rect 133512 159740 133564 159792
rect 157616 159740 157668 159792
rect 216772 159740 216824 159792
rect 218244 159740 218296 159792
rect 272524 159740 272576 159792
rect 277952 159740 278004 159792
rect 287060 159740 287112 159792
rect 287980 159740 288032 159792
rect 288624 159740 288676 159792
rect 298928 159740 298980 159792
rect 343640 159740 343692 159792
rect 366272 159740 366324 159792
rect 398472 159740 398524 159792
rect 399852 159740 399904 159792
rect 424232 159740 424284 159792
rect 451188 159740 451240 159792
rect 462872 159740 462924 159792
rect 463792 159740 463844 159792
rect 471796 159740 471848 159792
rect 478972 159740 479024 159792
rect 484584 159740 484636 159792
rect 46572 159672 46624 159724
rect 120172 159672 120224 159724
rect 124036 159672 124088 159724
rect 187700 159672 187752 159724
rect 194692 159672 194744 159724
rect 213644 159672 213696 159724
rect 214840 159672 214892 159724
rect 224592 159672 224644 159724
rect 224960 159672 225012 159724
rect 281448 159672 281500 159724
rect 282092 159672 282144 159724
rect 289912 159672 289964 159724
rect 292212 159672 292264 159724
rect 338764 159672 338816 159724
rect 352748 159672 352800 159724
rect 385960 159672 386012 159724
rect 388996 159672 389048 159724
rect 414296 159672 414348 159724
rect 420092 159672 420144 159724
rect 435824 159672 435876 159724
rect 458732 159672 458784 159724
rect 465080 159672 465132 159724
rect 53380 159604 53432 159656
rect 128360 159604 128412 159656
rect 130752 159604 130804 159656
rect 195244 159604 195296 159656
rect 211436 159604 211488 159656
rect 268936 159604 268988 159656
rect 285496 159604 285548 159656
rect 332600 159604 332652 159656
rect 346032 159604 346084 159656
rect 378140 159604 378192 159656
rect 382188 159604 382240 159656
rect 408500 159604 408552 159656
rect 413376 159604 413428 159656
rect 434444 159604 434496 159656
rect 441068 159604 441120 159656
rect 445668 159604 445720 159656
rect 447876 159604 447928 159656
rect 460204 159604 460256 159656
rect 468024 159604 468076 159656
rect 476028 159604 476080 159656
rect 80244 159536 80296 159588
rect 158444 159536 158496 159588
rect 170220 159536 170272 159588
rect 176660 159536 176712 159588
rect 198004 159536 198056 159588
rect 259644 159536 259696 159588
rect 272064 159536 272116 159588
rect 320732 159536 320784 159588
rect 339316 159536 339368 159588
rect 377956 159536 378008 159588
rect 379704 159536 379756 159588
rect 408776 159536 408828 159588
rect 431868 159536 431920 159588
rect 436376 159536 436428 159588
rect 449532 159536 449584 159588
rect 461492 159536 461544 159588
rect 470508 159536 470560 159588
rect 476120 159536 476172 159588
rect 100484 159468 100536 159520
rect 179420 159468 179472 159520
rect 184572 159468 184624 159520
rect 247224 159468 247276 159520
rect 251824 159468 251876 159520
rect 301688 159468 301740 159520
rect 308220 159468 308272 159520
rect 317788 159468 317840 159520
rect 319168 159468 319220 159520
rect 361580 159468 361632 159520
rect 368756 159468 368808 159520
rect 400404 159468 400456 159520
rect 402428 159468 402480 159520
rect 426164 159468 426216 159520
rect 433524 159468 433576 159520
rect 449808 159468 449860 159520
rect 453764 159468 453816 159520
rect 465264 159468 465316 159520
rect 467196 159468 467248 159520
rect 473360 159468 473412 159520
rect 482284 159468 482336 159520
rect 487252 159468 487304 159520
rect 26424 159400 26476 159452
rect 129832 159400 129884 159452
rect 139124 159400 139176 159452
rect 157340 159400 157392 159452
rect 177856 159400 177908 159452
rect 241704 159400 241756 159452
rect 245108 159400 245160 159452
rect 298744 159400 298796 159452
rect 312452 159400 312504 159452
rect 355232 159400 355284 159452
rect 359556 159400 359608 159452
rect 393412 159400 393464 159452
rect 395712 159400 395764 159452
rect 421104 159400 421156 159452
rect 432696 159400 432748 159452
rect 447140 159400 447192 159452
rect 448704 159400 448756 159452
rect 460940 159400 460992 159452
rect 468852 159400 468904 159452
rect 474832 159400 474884 159452
rect 477316 159400 477368 159452
rect 483296 159400 483348 159452
rect 518072 159400 518124 159452
rect 522672 159400 522724 159452
rect 12992 159332 13044 159384
rect 123944 159332 123996 159384
rect 132408 159332 132460 159384
rect 136088 159332 136140 159384
rect 140780 159332 140832 159384
rect 173992 159332 174044 159384
rect 191288 159332 191340 159384
rect 257344 159332 257396 159384
rect 287060 159332 287112 159384
rect 291476 159332 291528 159384
rect 331772 159332 331824 159384
rect 372068 159332 372120 159384
rect 372988 159332 373040 159384
rect 403164 159332 403216 159384
rect 426808 159332 426860 159384
rect 433248 159332 433300 159384
rect 434352 159332 434404 159384
rect 450084 159332 450136 159384
rect 452016 159332 452068 159384
rect 463976 159332 464028 159384
rect 469680 159332 469732 159384
rect 477408 159332 477460 159384
rect 478144 159332 478196 159384
rect 483940 159332 483992 159384
rect 518716 159332 518768 159384
rect 523500 159332 523552 159384
rect 93676 159264 93728 159316
rect 146024 159264 146076 159316
rect 181168 159264 181220 159316
rect 230664 159264 230716 159316
rect 237564 159264 237616 159316
rect 251732 159264 251784 159316
rect 271236 159264 271288 159316
rect 296812 159264 296864 159316
rect 298100 159264 298152 159316
rect 311992 159264 312044 159316
rect 325056 159264 325108 159316
rect 352012 159264 352064 159316
rect 461308 159264 461360 159316
rect 467932 159264 467984 159316
rect 109684 159196 109736 159248
rect 118700 159196 118752 159248
rect 144184 159196 144236 159248
rect 192576 159196 192628 159248
rect 208124 159196 208176 159248
rect 222108 159196 222160 159248
rect 227444 159196 227496 159248
rect 247040 159196 247092 159248
rect 250996 159196 251048 159248
rect 274640 159196 274692 159248
rect 284668 159196 284720 159248
rect 305460 159196 305512 159248
rect 460480 159196 460532 159248
rect 466644 159196 466696 159248
rect 110512 159128 110564 159180
rect 146116 159128 146168 159180
rect 155960 159128 156012 159180
rect 197636 159128 197688 159180
rect 201408 159128 201460 159180
rect 211896 159128 211948 159180
rect 257712 159128 257764 159180
rect 280068 159128 280120 159180
rect 304816 159128 304868 159180
rect 324320 159128 324372 159180
rect 446128 159128 446180 159180
rect 458364 159128 458416 159180
rect 462964 159128 463016 159180
rect 469220 159128 469272 159180
rect 37372 159060 37424 159112
rect 38568 159060 38620 159112
rect 91192 159060 91244 159112
rect 92388 159060 92440 159112
rect 127348 159060 127400 159112
rect 147680 159060 147732 159112
rect 174452 159060 174504 159112
rect 202972 159060 203024 159112
rect 214012 159060 214064 159112
rect 216680 159060 216732 159112
rect 247684 159060 247736 159112
rect 262128 159060 262180 159112
rect 264428 159060 264480 159112
rect 284300 159060 284352 159112
rect 459652 159060 459704 159112
rect 466460 159060 466512 159112
rect 471428 159060 471480 159112
rect 477684 159060 477736 159112
rect 210608 158992 210660 159044
rect 215024 158992 215076 159044
rect 267832 158992 267884 159044
rect 279516 158992 279568 159044
rect 288900 158992 288952 159044
rect 292304 158992 292356 159044
rect 455420 158992 455472 159044
rect 462964 158992 463016 159044
rect 473912 158992 473964 159044
rect 480720 158992 480772 159044
rect 507124 158992 507176 159044
rect 508412 158992 508464 159044
rect 118976 158924 119028 158976
rect 125508 158924 125560 158976
rect 224132 158924 224184 158976
rect 227720 158924 227772 158976
rect 278780 158924 278832 158976
rect 275376 158856 275428 158908
rect 278320 158856 278372 158908
rect 327540 158924 327592 158976
rect 328368 158924 328420 158976
rect 362040 158924 362092 158976
rect 366824 158924 366876 158976
rect 372160 158924 372212 158976
rect 374276 158924 374328 158976
rect 405740 158924 405792 158976
rect 407028 158924 407080 158976
rect 437756 158924 437808 158976
rect 444288 158924 444340 158976
rect 454592 158924 454644 158976
rect 461584 158924 461636 158976
rect 466368 158924 466420 158976
rect 472808 158924 472860 158976
rect 475568 158924 475620 158976
rect 482008 158924 482060 158976
rect 331772 158856 331824 158908
rect 456248 158856 456300 158908
rect 463148 158856 463200 158908
rect 465540 158856 465592 158908
rect 471980 158856 472032 158908
rect 474740 158856 474792 158908
rect 480260 158856 480312 158908
rect 480628 158856 480680 158908
rect 485964 158856 486016 158908
rect 508412 158856 508464 158908
rect 510068 158856 510120 158908
rect 145840 158788 145892 158840
rect 150440 158788 150492 158840
rect 196348 158788 196400 158840
rect 198740 158788 198792 158840
rect 261944 158788 261996 158840
rect 263416 158788 263468 158840
rect 268660 158788 268712 158840
rect 271696 158788 271748 158840
rect 315764 158788 315816 158840
rect 318708 158788 318760 158840
rect 336004 158788 336056 158840
rect 337936 158788 337988 158840
rect 436100 158788 436152 158840
rect 438860 158788 438912 158840
rect 464620 158788 464672 158840
rect 471612 158788 471664 158840
rect 476396 158788 476448 158840
rect 481640 158788 481692 158840
rect 499948 158788 500000 158840
rect 500592 158788 500644 158840
rect 506388 158788 506440 158840
rect 507584 158788 507636 158840
rect 388 158720 440 158772
rect 2044 158720 2096 158772
rect 64236 158720 64288 158772
rect 64788 158720 64840 158772
rect 71044 158720 71096 158772
rect 71688 158720 71740 158772
rect 77760 158720 77812 158772
rect 78588 158720 78640 158772
rect 84476 158720 84528 158772
rect 85488 158720 85540 158772
rect 103796 158720 103848 158772
rect 109040 158720 109092 158772
rect 121460 158720 121512 158772
rect 122748 158720 122800 158772
rect 129004 158720 129056 158772
rect 131120 158720 131172 158772
rect 131580 158720 131632 158772
rect 132408 158720 132460 158772
rect 145012 158720 145064 158772
rect 146208 158720 146260 158772
rect 152556 158720 152608 158772
rect 153108 158720 153160 158772
rect 165252 158720 165304 158772
rect 167644 158720 167696 158772
rect 202236 158720 202288 158772
rect 202788 158720 202840 158772
rect 203064 158720 203116 158772
rect 208492 158720 208544 158772
rect 220728 158720 220780 158772
rect 227904 158720 227956 158772
rect 230848 158720 230900 158772
rect 238668 158720 238720 158772
rect 241796 158720 241848 158772
rect 244648 158720 244700 158772
rect 256884 158720 256936 158772
rect 257988 158720 258040 158772
rect 261116 158720 261168 158772
rect 269028 158720 269080 158772
rect 281264 158720 281316 158772
rect 282552 158720 282604 158772
rect 286324 158720 286376 158772
rect 286876 158720 286928 158772
rect 301504 158720 301556 158772
rect 304816 158720 304868 158772
rect 378876 158720 378928 158772
rect 380992 158720 381044 158772
rect 385592 158720 385644 158772
rect 389088 158720 389140 158772
rect 389824 158720 389876 158772
rect 391572 158720 391624 158772
rect 452844 158720 452896 158772
rect 460112 158720 460164 158772
rect 462136 158720 462188 158772
rect 467840 158720 467892 158772
rect 473084 158720 473136 158772
rect 478972 158720 479024 158772
rect 481456 158720 481508 158772
rect 486424 158720 486476 158772
rect 504456 158720 504508 158772
rect 505008 158720 505060 158772
rect 505836 158720 505888 158772
rect 506756 158720 506808 158772
rect 509700 158720 509752 158772
rect 511724 158720 511776 158772
rect 514852 158720 514904 158772
rect 518532 158720 518584 158772
rect 99564 158652 99616 158704
rect 194968 158652 195020 158704
rect 220176 158652 220228 158704
rect 277952 158652 278004 158704
rect 279608 158652 279660 158704
rect 331312 158652 331364 158704
rect 86132 158584 86184 158636
rect 183560 158584 183612 158636
rect 200580 158584 200632 158636
rect 272064 158584 272116 158636
rect 274548 158584 274600 158636
rect 328552 158584 328604 158636
rect 351920 158584 351972 158636
rect 386512 158584 386564 158636
rect 62580 158516 62632 158568
rect 166724 158516 166776 158568
rect 197176 158516 197228 158568
rect 269396 158516 269448 158568
rect 272892 158516 272944 158568
rect 327080 158516 327132 158568
rect 350264 158516 350316 158568
rect 385224 158516 385276 158568
rect 65984 158448 66036 158500
rect 168380 158448 168432 158500
rect 190460 158448 190512 158500
rect 263784 158448 263836 158500
rect 266176 158448 266228 158500
rect 322112 158448 322164 158500
rect 338488 158448 338540 158500
rect 376852 158448 376904 158500
rect 377220 158448 377272 158500
rect 406844 158448 406896 158500
rect 59268 158380 59320 158432
rect 163044 158380 163096 158432
rect 187056 158380 187108 158432
rect 260840 158380 260892 158432
rect 262772 158380 262824 158432
rect 319536 158380 319588 158432
rect 330116 158380 330168 158432
rect 370872 158380 370924 158432
rect 52460 158312 52512 158364
rect 158996 158312 159048 158364
rect 177028 158312 177080 158364
rect 254032 158312 254084 158364
rect 256056 158312 256108 158364
rect 314384 158312 314436 158364
rect 317420 158312 317472 158364
rect 360200 158312 360252 158364
rect 378048 158312 378100 158364
rect 407396 158312 407448 158364
rect 45744 158244 45796 158296
rect 153384 158244 153436 158296
rect 173624 158244 173676 158296
rect 251456 158244 251508 158296
rect 252652 158244 252704 158296
rect 310612 158244 310664 158296
rect 320824 158244 320876 158296
rect 363512 158244 363564 158296
rect 367100 158244 367152 158296
rect 399116 158244 399168 158296
rect 31484 158176 31536 158228
rect 139492 158176 139544 158228
rect 163504 158176 163556 158228
rect 242900 158176 242952 158228
rect 245936 158176 245988 158228
rect 306380 158176 306432 158228
rect 314108 158176 314160 158228
rect 357624 158176 357676 158228
rect 361212 158176 361264 158228
rect 394700 158176 394752 158228
rect 404084 158176 404136 158228
rect 427360 158312 427412 158364
rect 439412 158244 439464 158296
rect 454408 158244 454460 158296
rect 426440 158176 426492 158228
rect 443000 158176 443052 158228
rect 35716 158108 35768 158160
rect 145104 158108 145156 158160
rect 153476 158108 153528 158160
rect 236092 158108 236144 158160
rect 242624 158108 242676 158160
rect 304080 158108 304132 158160
rect 307392 158108 307444 158160
rect 353300 158108 353352 158160
rect 358636 158108 358688 158160
rect 391940 158108 391992 158160
rect 404912 158108 404964 158160
rect 428004 158108 428056 158160
rect 428464 158108 428516 158160
rect 445760 158108 445812 158160
rect 18880 158040 18932 158092
rect 132500 158040 132552 158092
rect 139952 158040 140004 158092
rect 224960 158040 225012 158092
rect 229100 158040 229152 158092
rect 292764 158040 292816 158092
rect 293040 158040 293092 158092
rect 342260 158040 342312 158092
rect 351092 158040 351144 158092
rect 386972 158040 387024 158092
rect 393964 158040 394016 158092
rect 419540 158040 419592 158092
rect 420920 158040 420972 158092
rect 440332 158040 440384 158092
rect 443644 158040 443696 158092
rect 456800 158040 456852 158092
rect 2136 157972 2188 158024
rect 120080 157972 120132 158024
rect 133236 157972 133288 158024
rect 220636 157972 220688 158024
rect 225696 157972 225748 158024
rect 288440 157972 288492 158024
rect 289728 157972 289780 158024
rect 340052 157972 340104 158024
rect 340144 157972 340196 158024
rect 378600 157972 378652 158024
rect 388076 157972 388128 158024
rect 414572 157972 414624 158024
rect 415032 157972 415084 158024
rect 434720 157972 434772 158024
rect 435180 157972 435232 158024
rect 451188 157972 451240 158024
rect 106372 157904 106424 157956
rect 200120 157904 200172 157956
rect 207020 157904 207072 157956
rect 233240 157904 233292 157956
rect 239220 157904 239272 157956
rect 252008 157904 252060 157956
rect 259460 157904 259512 157956
rect 316960 157904 317012 157956
rect 321652 157904 321704 157956
rect 359464 157904 359516 157956
rect 123116 157836 123168 157888
rect 205640 157836 205692 157888
rect 221556 157836 221608 157888
rect 245660 157836 245712 157888
rect 269488 157836 269540 157888
rect 79416 157768 79468 157820
rect 146116 157768 146168 157820
rect 147680 157768 147732 157820
rect 215392 157768 215444 157820
rect 311900 157768 311952 157820
rect 324320 157836 324372 157888
rect 350540 157836 350592 157888
rect 146024 157700 146076 157752
rect 190460 157700 190512 157752
rect 201316 157700 201368 157752
rect 223856 157700 223908 157752
rect 324688 157768 324740 157820
rect 341340 157768 341392 157820
rect 76012 157292 76064 157344
rect 177028 157292 177080 157344
rect 193772 157292 193824 157344
rect 266912 157292 266964 157344
rect 296444 157292 296496 157344
rect 345020 157292 345072 157344
rect 356152 157292 356204 157344
rect 358820 157292 358872 157344
rect 69296 157224 69348 157276
rect 171140 157224 171192 157276
rect 179512 157224 179564 157276
rect 255872 157224 255924 157276
rect 276204 157224 276256 157276
rect 329840 157224 329892 157276
rect 352012 157224 352064 157276
rect 365904 157224 365956 157276
rect 4528 157156 4580 157208
rect 109132 157156 109184 157208
rect 113088 157156 113140 157208
rect 205272 157156 205324 157208
rect 209780 157156 209832 157208
rect 279056 157156 279108 157208
rect 288624 157156 288676 157208
rect 338672 157156 338724 157208
rect 347780 157156 347832 157208
rect 384396 157156 384448 157208
rect 55864 157088 55916 157140
rect 161572 157088 161624 157140
rect 172796 157088 172848 157140
rect 250812 157088 250864 157140
rect 260288 157088 260340 157140
rect 317420 157088 317472 157140
rect 346860 157088 346912 157140
rect 383752 157088 383804 157140
rect 49148 157020 49200 157072
rect 156420 157020 156472 157072
rect 176108 157020 176160 157072
rect 252560 157020 252612 157072
rect 254400 157020 254452 157072
rect 311900 157020 311952 157072
rect 336832 157020 336884 157072
rect 376024 157020 376076 157072
rect 383108 157020 383160 157072
rect 411352 157020 411404 157072
rect 39028 156952 39080 157004
rect 147680 156952 147732 157004
rect 169392 156952 169444 157004
rect 247132 156952 247184 157004
rect 253572 156952 253624 157004
rect 307024 156952 307076 157004
rect 330944 156952 330996 157004
rect 371240 156952 371292 157004
rect 373816 156952 373868 157004
rect 404084 156952 404136 157004
rect 423404 156952 423456 157004
rect 442172 156952 442224 157004
rect 24768 156884 24820 156936
rect 137836 156884 137888 156936
rect 160192 156884 160244 156936
rect 241244 156884 241296 156936
rect 249340 156884 249392 156936
rect 306380 156884 306432 156936
rect 21364 156816 21416 156868
rect 135260 156816 135312 156868
rect 150072 156816 150124 156868
rect 233516 156816 233568 156868
rect 246764 156816 246816 156868
rect 307300 156884 307352 156936
rect 310704 156884 310756 156936
rect 356152 156884 356204 156936
rect 374644 156884 374696 156936
rect 404452 156884 404504 156936
rect 411628 156884 411680 156936
rect 433156 156884 433208 156936
rect 306656 156816 306708 156868
rect 351920 156816 351972 156868
rect 363696 156816 363748 156868
rect 396540 156816 396592 156868
rect 401600 156816 401652 156868
rect 425152 156816 425204 156868
rect 433064 156816 433116 156868
rect 447324 156816 447376 156868
rect 18052 156748 18104 156800
rect 132684 156748 132736 156800
rect 136640 156748 136692 156800
rect 222752 156748 222804 156800
rect 236736 156748 236788 156800
rect 299480 156748 299532 156800
rect 299756 156748 299808 156800
rect 347780 156748 347832 156800
rect 348608 156748 348660 156800
rect 385040 156748 385092 156800
rect 387248 156748 387300 156800
rect 414112 156748 414164 156800
rect 414204 156748 414256 156800
rect 435088 156748 435140 156800
rect 436376 156748 436428 156800
rect 448612 156748 448664 156800
rect 11244 156680 11296 156732
rect 125692 156680 125744 156732
rect 126520 156680 126572 156732
rect 215484 156680 215536 156732
rect 216680 156680 216732 156732
rect 282092 156680 282144 156732
rect 283012 156680 283064 156732
rect 334900 156680 334952 156732
rect 341892 156680 341944 156732
rect 379888 156680 379940 156732
rect 384764 156680 384816 156732
rect 412640 156680 412692 156732
rect 419264 156680 419316 156732
rect 438952 156680 439004 156732
rect 14648 156612 14700 156664
rect 129740 156612 129792 156664
rect 129924 156612 129976 156664
rect 218060 156612 218112 156664
rect 240048 156612 240100 156664
rect 302240 156612 302292 156664
rect 303988 156612 304040 156664
rect 351000 156612 351052 156664
rect 357808 156612 357860 156664
rect 392124 156612 392176 156664
rect 400772 156612 400824 156664
rect 423772 156612 423824 156664
rect 427636 156612 427688 156664
rect 444380 156612 444432 156664
rect 445300 156612 445352 156664
rect 458824 156612 458876 156664
rect 96252 156544 96304 156596
rect 192392 156544 192444 156596
rect 215024 156544 215076 156596
rect 278780 156544 278832 156596
rect 303160 156544 303212 156596
rect 349252 156544 349304 156596
rect 116400 156476 116452 156528
rect 207020 156476 207072 156528
rect 227720 156476 227772 156528
rect 290004 156476 290056 156528
rect 307024 156476 307076 156528
rect 312452 156476 312504 156528
rect 317788 156476 317840 156528
rect 354220 156476 354272 156528
rect 135628 156408 135680 156460
rect 169944 156408 169996 156460
rect 176660 156408 176712 156460
rect 248880 156408 248932 156460
rect 251732 156408 251784 156460
rect 300308 156408 300360 156460
rect 306380 156408 306432 156460
rect 309232 156408 309284 156460
rect 311992 156408 312044 156460
rect 346492 156408 346544 156460
rect 133512 156340 133564 156392
rect 164424 156340 164476 156392
rect 279516 156340 279568 156392
rect 323400 156340 323452 156392
rect 72700 155864 72752 155916
rect 174452 155864 174504 155916
rect 203892 155864 203944 155916
rect 273444 155864 273496 155916
rect 324228 155864 324280 155916
rect 366272 155864 366324 155916
rect 378140 155864 378192 155916
rect 382280 155864 382332 155916
rect 55036 155796 55088 155848
rect 160100 155796 160152 155848
rect 206468 155796 206520 155848
rect 276480 155796 276532 155848
rect 287152 155796 287204 155848
rect 338120 155796 338172 155848
rect 346308 155796 346360 155848
rect 352288 155796 352340 155848
rect 48320 155728 48372 155780
rect 154672 155728 154724 155780
rect 199660 155728 199712 155780
rect 271052 155728 271104 155780
rect 280436 155728 280488 155780
rect 333060 155728 333112 155780
rect 336648 155728 336700 155780
rect 361948 155728 362000 155780
rect 362132 155728 362184 155780
rect 367652 155728 367704 155780
rect 370412 155728 370464 155780
rect 401692 155728 401744 155780
rect 41604 155660 41656 155712
rect 150624 155660 150676 155712
rect 192944 155660 192996 155712
rect 265164 155660 265216 155712
rect 277124 155660 277176 155712
rect 330024 155660 330076 155712
rect 334256 155660 334308 155712
rect 374092 155660 374144 155712
rect 23940 155592 23992 155644
rect 136732 155592 136784 155644
rect 160284 155592 160336 155644
rect 185032 155592 185084 155644
rect 186228 155592 186280 155644
rect 261116 155592 261168 155644
rect 273720 155592 273772 155644
rect 327908 155592 327960 155644
rect 328368 155592 328420 155644
rect 368940 155592 368992 155644
rect 369584 155592 369636 155644
rect 400220 155592 400272 155644
rect 22192 155524 22244 155576
rect 135812 155524 135864 155576
rect 150440 155524 150492 155576
rect 229192 155524 229244 155576
rect 230020 155524 230072 155576
rect 294512 155524 294564 155576
rect 297272 155524 297324 155576
rect 345848 155524 345900 155576
rect 364524 155524 364576 155576
rect 396172 155524 396224 155576
rect 15476 155456 15528 155508
rect 130292 155456 130344 155508
rect 156788 155456 156840 155508
rect 238576 155456 238628 155508
rect 238668 155456 238720 155508
rect 294052 155456 294104 155508
rect 294788 155456 294840 155508
rect 343916 155456 343968 155508
rect 353668 155456 353720 155508
rect 388352 155456 388404 155508
rect 408316 155456 408368 155508
rect 430580 155456 430632 155508
rect 433248 155456 433300 155508
rect 444748 155456 444800 155508
rect 8760 155388 8812 155440
rect 125600 155388 125652 155440
rect 138296 155388 138348 155440
rect 222016 155388 222068 155440
rect 225788 155388 225840 155440
rect 291292 155388 291344 155440
rect 293868 155388 293920 155440
rect 343272 155388 343324 155440
rect 344376 155388 344428 155440
rect 380900 155388 380952 155440
rect 394884 155388 394936 155440
rect 420368 155388 420420 155440
rect 429292 155388 429344 155440
rect 446680 155388 446732 155440
rect 2872 155320 2924 155372
rect 121092 155320 121144 155372
rect 146668 155320 146720 155372
rect 230940 155320 230992 155372
rect 232504 155320 232556 155372
rect 296444 155320 296496 155372
rect 300676 155320 300728 155372
rect 348424 155320 348476 155372
rect 354496 155320 354548 155372
rect 389548 155320 389600 155372
rect 397368 155320 397420 155372
rect 422300 155320 422352 155372
rect 424324 155320 424376 155372
rect 441712 155320 441764 155372
rect 444472 155320 444524 155372
rect 458180 155320 458232 155372
rect 5356 155252 5408 155304
rect 123024 155252 123076 155304
rect 136088 155252 136140 155304
rect 219532 155252 219584 155304
rect 223212 155252 223264 155304
rect 289360 155252 289412 155304
rect 290556 155252 290608 155304
rect 339592 155252 339644 155304
rect 345204 155252 345256 155304
rect 382464 155252 382516 155304
rect 383936 155252 383988 155304
rect 411996 155252 412048 155304
rect 421748 155252 421800 155304
rect 440884 155252 440936 155304
rect 441988 155252 442040 155304
rect 455972 155252 456024 155304
rect 1216 155184 1268 155236
rect 118792 155184 118844 155236
rect 125784 155184 125836 155236
rect 214840 155184 214892 155236
rect 216496 155184 216548 155236
rect 283104 155184 283156 155236
rect 283840 155184 283892 155236
rect 335544 155184 335596 155236
rect 343548 155184 343600 155236
rect 381176 155184 381228 155236
rect 381360 155184 381412 155236
rect 410064 155184 410116 155236
rect 410800 155184 410852 155236
rect 432052 155184 432104 155236
rect 442816 155184 442868 155236
rect 456984 155184 457036 155236
rect 89536 155116 89588 155168
rect 187240 155116 187292 155168
rect 219072 155116 219124 155168
rect 286140 155116 286192 155168
rect 291476 155116 291528 155168
rect 331128 155116 331180 155168
rect 118700 155048 118752 155100
rect 201592 155048 201644 155100
rect 226616 155048 226668 155100
rect 291200 155048 291252 155100
rect 330208 155048 330260 155100
rect 356796 155116 356848 155168
rect 128176 154980 128228 155032
rect 197452 154980 197504 155032
rect 269028 154980 269080 155032
rect 317972 154980 318024 155032
rect 120172 154912 120224 154964
rect 154212 154912 154264 154964
rect 157340 154912 157392 154964
rect 225144 154912 225196 154964
rect 262128 154912 262180 154964
rect 307944 154912 307996 154964
rect 134892 154844 134944 154896
rect 197360 154844 197412 154896
rect 118148 154776 118200 154828
rect 144828 154776 144880 154828
rect 183284 154776 183336 154828
rect 209964 154776 210016 154828
rect 103428 154504 103480 154556
rect 197544 154504 197596 154556
rect 215668 154504 215720 154556
rect 283564 154504 283616 154556
rect 284300 154504 284352 154556
rect 320916 154504 320968 154556
rect 338764 154504 338816 154556
rect 341984 154504 342036 154556
rect 92848 154436 92900 154488
rect 189816 154436 189868 154488
rect 198740 154436 198792 154488
rect 268844 154436 268896 154488
rect 274640 154436 274692 154488
rect 310520 154436 310572 154488
rect 319996 154436 320048 154488
rect 363236 154436 363288 154488
rect 366824 154436 366876 154488
rect 395344 154436 395396 154488
rect 58348 154368 58400 154420
rect 156604 154368 156656 154420
rect 192116 154368 192168 154420
rect 265716 154368 265768 154420
rect 267004 154368 267056 154420
rect 322848 154368 322900 154420
rect 335084 154368 335136 154420
rect 338764 154368 338816 154420
rect 340972 154368 341024 154420
rect 379244 154368 379296 154420
rect 51632 154300 51684 154352
rect 158352 154300 158404 154352
rect 158444 154300 158496 154352
rect 180248 154300 180300 154352
rect 185400 154300 185452 154352
rect 260472 154300 260524 154352
rect 270316 154300 270368 154352
rect 325332 154300 325384 154352
rect 326988 154300 327040 154352
rect 368388 154300 368440 154352
rect 44916 154232 44968 154284
rect 153200 154232 153252 154284
rect 154304 154232 154356 154284
rect 183284 154232 183336 154284
rect 188804 154232 188856 154284
rect 263048 154232 263100 154284
rect 263600 154232 263652 154284
rect 320180 154232 320232 154284
rect 323308 154232 323360 154284
rect 365720 154232 365772 154284
rect 371332 154232 371384 154284
rect 402336 154232 402388 154284
rect 34796 154164 34848 154216
rect 145564 154164 145616 154216
rect 147772 154164 147824 154216
rect 177672 154164 177724 154216
rect 181996 154164 182048 154216
rect 257896 154164 257948 154216
rect 257988 154164 258040 154216
rect 315028 154164 315080 154216
rect 316592 154164 316644 154216
rect 360660 154164 360712 154216
rect 368296 154164 368348 154216
rect 399760 154164 399812 154216
rect 422576 154164 422628 154216
rect 25596 154096 25648 154148
rect 138480 154096 138532 154148
rect 156604 154096 156656 154148
rect 163504 154096 163556 154148
rect 172428 154096 172480 154148
rect 250168 154096 250220 154148
rect 250260 154096 250312 154148
rect 309876 154096 309928 154148
rect 313280 154096 313332 154148
rect 358084 154096 358136 154148
rect 360384 154096 360436 154148
rect 394056 154096 394108 154148
rect 407488 154096 407540 154148
rect 429936 154096 429988 154148
rect 13820 154028 13872 154080
rect 129464 154028 129516 154080
rect 131120 154028 131172 154080
rect 217416 154028 217468 154080
rect 219900 154028 219952 154080
rect 286784 154028 286836 154080
rect 286876 154028 286928 154080
rect 337476 154028 337528 154080
rect 338028 154028 338080 154080
rect 376576 154028 376628 154080
rect 398196 154028 398248 154080
rect 422944 154028 422996 154080
rect 438860 154164 438912 154216
rect 451832 154164 451884 154216
rect 431040 154096 431092 154148
rect 447968 154096 448020 154148
rect 441436 154028 441488 154080
rect 20536 153960 20588 154012
rect 134616 153960 134668 154012
rect 143356 153960 143408 154012
rect 228364 153960 228416 154012
rect 243452 153960 243504 154012
rect 304724 153960 304776 154012
rect 304816 153960 304868 154012
rect 349068 153960 349120 154012
rect 355324 153960 355376 154012
rect 17132 153892 17184 153944
rect 132040 153892 132092 153944
rect 135904 153892 135956 153944
rect 222568 153892 222620 153944
rect 233332 153892 233384 153944
rect 297088 153892 297140 153944
rect 309968 153892 310020 153944
rect 355508 153892 355560 153944
rect 357348 153960 357400 154012
rect 391480 153960 391532 154012
rect 391848 153960 391900 154012
rect 417792 153960 417844 154012
rect 425244 153960 425296 154012
rect 443460 153960 443512 154012
rect 390192 153892 390244 153944
rect 390652 153892 390704 153944
rect 417148 153892 417200 153944
rect 418436 153892 418488 153944
rect 438308 153892 438360 153944
rect 440240 153892 440292 153944
rect 455052 153892 455104 153944
rect 4068 153824 4120 153876
rect 121736 153824 121788 153876
rect 122656 153824 122708 153876
rect 212264 153824 212316 153876
rect 213184 153824 213236 153876
rect 281632 153824 281684 153876
rect 282552 153824 282604 153876
rect 333704 153824 333756 153876
rect 105452 153756 105504 153808
rect 199476 153756 199528 153808
rect 208492 153756 208544 153808
rect 273904 153756 273956 153808
rect 280068 153756 280120 153808
rect 315672 153756 315724 153808
rect 333428 153756 333480 153808
rect 373448 153824 373500 153876
rect 380808 153824 380860 153876
rect 409420 153824 409472 153876
rect 417516 153824 417568 153876
rect 437664 153824 437716 153876
rect 438584 153824 438636 153876
rect 453764 153824 453816 153876
rect 63408 153688 63460 153740
rect 118700 153688 118752 153740
rect 119804 153688 119856 153740
rect 208400 153688 208452 153740
rect 244280 153688 244332 153740
rect 305368 153688 305420 153740
rect 305460 153688 305512 153740
rect 336188 153688 336240 153740
rect 128360 153620 128412 153672
rect 159640 153620 159692 153672
rect 168564 153620 168616 153672
rect 215300 153620 215352 153672
rect 263600 153620 263652 153672
rect 263784 153620 263836 153672
rect 296812 153620 296864 153672
rect 325976 153620 326028 153672
rect 197636 153552 197688 153604
rect 238024 153552 238076 153604
rect 109040 153144 109092 153196
rect 198188 153144 198240 153196
rect 202972 153144 203024 153196
rect 252100 153144 252152 153196
rect 259644 153144 259696 153196
rect 270132 153144 270184 153196
rect 272524 153144 272576 153196
rect 285496 153144 285548 153196
rect 292304 153144 292356 153196
rect 339408 153144 339460 153196
rect 355232 153144 355284 153196
rect 357440 153144 357492 153196
rect 368480 153144 368532 153196
rect 372804 153144 372856 153196
rect 385960 153144 386012 153196
rect 388260 153144 388312 153196
rect 408500 153144 408552 153196
rect 410708 153144 410760 153196
rect 435824 153144 435876 153196
rect 439596 153144 439648 153196
rect 447140 153144 447192 153196
rect 449256 153144 449308 153196
rect 461584 153144 461636 153196
rect 465908 153144 465960 153196
rect 466460 153144 466512 153196
rect 469772 153144 469824 153196
rect 471612 153144 471664 153196
rect 473636 153144 473688 153196
rect 474832 153144 474884 153196
rect 476948 153144 477000 153196
rect 485688 153144 485740 153196
rect 489644 153144 489696 153196
rect 490748 153144 490800 153196
rect 493508 153144 493560 153196
rect 494060 153144 494112 153196
rect 496084 153144 496136 153196
rect 496636 153144 496688 153196
rect 498016 153144 498068 153196
rect 498292 153144 498344 153196
rect 499304 153144 499356 153196
rect 500960 153144 501012 153196
rect 501880 153144 501932 153196
rect 510988 153144 511040 153196
rect 513472 153144 513524 153196
rect 514208 153144 514260 153196
rect 517428 153144 517480 153196
rect 117228 153076 117280 153128
rect 208492 153076 208544 153128
rect 215300 153076 215352 153128
rect 247592 153076 247644 153128
rect 252008 153076 252060 153128
rect 301596 153076 301648 153128
rect 301688 153076 301740 153128
rect 311164 153076 311216 153128
rect 113916 153008 113968 153060
rect 205916 153008 205968 153060
rect 216772 153008 216824 153060
rect 239312 153008 239364 153060
rect 239956 153008 240008 153060
rect 293224 153008 293276 153060
rect 298744 153008 298796 153060
rect 306012 153008 306064 153060
rect 311072 153008 311124 153060
rect 321468 153076 321520 153128
rect 338764 153076 338816 153128
rect 374736 153076 374788 153128
rect 463148 153076 463200 153128
rect 467196 153076 467248 153128
rect 471980 153076 472032 153128
rect 474280 153076 474332 153128
rect 476120 153076 476172 153128
rect 478144 153076 478196 153128
rect 484860 153076 484912 153128
rect 489000 153076 489052 153128
rect 489920 153076 489972 153128
rect 492864 153076 492916 153128
rect 493232 153076 493284 153128
rect 495440 153076 495492 153128
rect 495808 153076 495860 153128
rect 497372 153076 497424 153128
rect 497464 153076 497516 153128
rect 498660 153076 498712 153128
rect 512920 153076 512972 153128
rect 515312 153076 515364 153128
rect 318708 153008 318760 153060
rect 360016 153008 360068 153060
rect 399024 153008 399076 153060
rect 423588 153008 423640 153060
rect 462964 153008 463016 153060
rect 466552 153008 466604 153060
rect 466644 153008 466696 153060
rect 470416 153008 470468 153060
rect 472808 153008 472860 153060
rect 474924 153008 474976 153060
rect 484308 153008 484360 153060
rect 488264 153008 488316 153060
rect 492404 153008 492456 153060
rect 494796 153008 494848 153060
rect 495256 153008 495308 153060
rect 496728 153008 496780 153060
rect 107476 152940 107528 152992
rect 200764 152940 200816 152992
rect 205640 152940 205692 152992
rect 212908 152940 212960 152992
rect 213644 152940 213696 152992
rect 267556 152940 267608 152992
rect 271696 152940 271748 152992
rect 324044 152940 324096 152992
rect 337936 152940 337988 152992
rect 375380 152940 375432 152992
rect 389088 152940 389140 152992
rect 413284 152940 413336 152992
rect 415860 152940 415912 152992
rect 436376 152940 436428 152992
rect 465080 152940 465132 152992
rect 469128 152940 469180 152992
rect 471796 152940 471848 152992
rect 472992 152940 473044 152992
rect 473360 152940 473412 152992
rect 475568 152940 475620 152992
rect 483204 152940 483256 152992
rect 487804 152940 487856 152992
rect 491576 152940 491628 152992
rect 494152 152940 494204 152992
rect 512276 152940 512328 152992
rect 514760 152940 514812 152992
rect 97080 152872 97132 152924
rect 193036 152872 193088 152924
rect 210148 152872 210200 152924
rect 262404 152872 262456 152924
rect 263416 152872 263468 152924
rect 318892 152872 318944 152924
rect 328276 152872 328328 152924
rect 369584 152872 369636 152924
rect 372620 152872 372672 152924
rect 380532 152872 380584 152924
rect 380992 152872 381044 152924
rect 408132 152872 408184 152924
rect 409972 152872 410024 152924
rect 431868 152872 431920 152924
rect 464712 152872 464764 152924
rect 468392 152872 468444 152924
rect 90364 152804 90416 152856
rect 187884 152804 187936 152856
rect 192576 152804 192628 152856
rect 229008 152804 229060 152856
rect 244648 152804 244700 152856
rect 303528 152804 303580 152856
rect 305000 152804 305052 152856
rect 316316 152804 316368 152856
rect 322756 152804 322808 152856
rect 365168 152804 365220 152856
rect 374276 152804 374328 152856
rect 402980 152804 403032 152856
rect 412548 152804 412600 152856
rect 433800 152804 433852 152856
rect 510344 152804 510396 152856
rect 512000 152804 512052 152856
rect 84108 152736 84160 152788
rect 182732 152736 182784 152788
rect 187700 152736 187752 152788
rect 213552 152736 213604 152788
rect 222016 152736 222068 152788
rect 224500 152736 224552 152788
rect 224592 152736 224644 152788
rect 282920 152736 282972 152788
rect 284392 152736 284444 152788
rect 295800 152736 295852 152788
rect 295892 152736 295944 152788
rect 344560 152736 344612 152788
rect 358820 152736 358872 152788
rect 390836 152736 390888 152788
rect 391572 152736 391624 152788
rect 416504 152736 416556 152788
rect 416688 152736 416740 152788
rect 437020 152736 437072 152788
rect 73528 152668 73580 152720
rect 175096 152668 175148 152720
rect 179420 152668 179472 152720
rect 195612 152668 195664 152720
rect 211896 152668 211948 152720
rect 272708 152668 272760 152720
rect 278320 152668 278372 152720
rect 329196 152668 329248 152720
rect 329288 152668 329340 152720
rect 370228 152668 370280 152720
rect 376668 152668 376720 152720
rect 406200 152668 406252 152720
rect 407028 152668 407080 152720
rect 428648 152668 428700 152720
rect 444288 152668 444340 152720
rect 453120 152668 453172 152720
rect 34428 152600 34480 152652
rect 144920 152600 144972 152652
rect 167736 152600 167788 152652
rect 246948 152600 247000 152652
rect 255228 152600 255280 152652
rect 313740 152600 313792 152652
rect 314936 152600 314988 152652
rect 359372 152600 359424 152652
rect 362960 152600 363012 152652
rect 395988 152600 396040 152652
rect 396632 152600 396684 152652
rect 421656 152600 421708 152652
rect 445668 152600 445720 152652
rect 455696 152600 455748 152652
rect 23388 152532 23440 152584
rect 136548 152532 136600 152584
rect 147588 152532 147640 152584
rect 231584 152532 231636 152584
rect 248512 152532 248564 152584
rect 308588 152532 308640 152584
rect 309048 152532 309100 152584
rect 354864 152532 354916 152584
rect 365444 152532 365496 152584
rect 397828 152532 397880 152584
rect 403256 152532 403308 152584
rect 426808 152532 426860 152584
rect 446956 152532 447008 152584
rect 460020 152532 460072 152584
rect 460112 152532 460164 152584
rect 464620 152532 464672 152584
rect 6276 152464 6328 152516
rect 123668 152464 123720 152516
rect 125692 152464 125744 152516
rect 127532 152464 127584 152516
rect 134064 152464 134116 152516
rect 221280 152464 221332 152516
rect 234988 152464 235040 152516
rect 298376 152464 298428 152516
rect 302332 152464 302384 152516
rect 349712 152464 349764 152516
rect 109132 152396 109184 152448
rect 122380 152396 122432 152448
rect 123944 152396 123996 152448
rect 128820 152396 128872 152448
rect 129832 152396 129884 152448
rect 139124 152396 139176 152448
rect 144828 152396 144880 152448
rect 209136 152396 209188 152448
rect 221924 152396 221976 152448
rect 244372 152396 244424 152448
rect 245660 152396 245712 152448
rect 288072 152396 288124 152448
rect 289912 152396 289964 152448
rect 334348 152396 334400 152448
rect 349436 152396 349488 152448
rect 385592 152464 385644 152516
rect 392308 152464 392360 152516
rect 418436 152464 418488 152516
rect 437388 152464 437440 152516
rect 452476 152464 452528 152516
rect 414296 152396 414348 152448
rect 415860 152396 415912 152448
rect 118700 152328 118752 152380
rect 167368 152328 167420 152380
rect 183284 152328 183336 152380
rect 236736 152328 236788 152380
rect 247224 152328 247276 152380
rect 259828 152328 259880 152380
rect 268936 152328 268988 152380
rect 280344 152328 280396 152380
rect 288348 152328 288400 152380
rect 300952 152328 301004 152380
rect 511632 152328 511684 152380
rect 513564 152328 513616 152380
rect 173992 152260 174044 152312
rect 226432 152260 226484 152312
rect 230664 152260 230716 152312
rect 257252 152260 257304 152312
rect 257344 152260 257396 152312
rect 264980 152260 265032 152312
rect 265072 152260 265124 152312
rect 275100 152260 275152 152312
rect 281448 152260 281500 152312
rect 290648 152260 290700 152312
rect 146116 152192 146168 152244
rect 179604 152192 179656 152244
rect 197360 152192 197412 152244
rect 221924 152192 221976 152244
rect 230388 152192 230440 152244
rect 249524 152192 249576 152244
rect 513564 152192 513616 152244
rect 516140 152192 516192 152244
rect 26700 152124 26752 152176
rect 110144 152124 110196 152176
rect 197452 152124 197504 152176
rect 216772 152124 216824 152176
rect 241704 152124 241756 152176
rect 254676 152124 254728 152176
rect 516692 152124 516744 152176
rect 520280 152124 520332 152176
rect 102324 152056 102376 152108
rect 109960 152056 110012 152108
rect 515496 152056 515548 152108
rect 518900 152056 518952 152108
rect 40500 151988 40552 152040
rect 89168 151988 89220 152040
rect 95516 151988 95568 152040
rect 114376 151988 114428 152040
rect 467840 151988 467892 152040
rect 471704 151988 471756 152040
rect 488172 151988 488224 152040
rect 491576 151988 491628 152040
rect 515956 151988 516008 152040
rect 519452 151988 519504 152040
rect 88616 151920 88668 151972
rect 110328 151920 110380 151972
rect 136364 151920 136416 151972
rect 144276 151920 144328 151972
rect 469220 151920 469272 151972
rect 472348 151920 472400 151972
rect 487344 151920 487396 151972
rect 490932 151920 490984 151972
rect 507676 151920 507728 151972
rect 509240 151920 509292 151972
rect 517428 151920 517480 151972
rect 521568 151920 521620 151972
rect 33600 151852 33652 151904
rect 110236 151852 110288 151904
rect 127624 151852 127676 151904
rect 133972 151852 134024 151904
rect 139492 151852 139544 151904
rect 142988 151852 143040 151904
rect 236000 151852 236052 151904
rect 240600 151852 240652 151904
rect 320732 151852 320784 151904
rect 326620 151852 326672 151904
rect 332600 151852 332652 151904
rect 336832 151852 336884 151904
rect 343640 151852 343692 151904
rect 347136 151852 347188 151904
rect 359464 151852 359516 151904
rect 364524 151852 364576 151904
rect 456064 151852 456116 151904
rect 462688 151852 462740 151904
rect 464344 151852 464396 151904
rect 467840 151852 467892 151904
rect 467932 151852 467984 151904
rect 471060 151852 471112 151904
rect 486516 151852 486568 151904
rect 489092 151852 489144 151904
rect 492220 151852 492272 151904
rect 499488 151852 499540 151904
rect 499948 151852 500000 151904
rect 81716 151784 81768 151836
rect 97724 151784 97776 151836
rect 105820 151784 105872 151836
rect 106924 151784 106976 151836
rect 208400 151784 208452 151836
rect 210424 151784 210476 151836
rect 490288 151784 490340 151836
rect 509056 151784 509108 151836
rect 510896 151784 510948 151836
rect 132408 151716 132460 151768
rect 219348 151716 219400 151768
rect 122748 151648 122800 151700
rect 211620 151648 211672 151700
rect 111708 151580 111760 151632
rect 203984 151580 204036 151632
rect 104808 151512 104860 151564
rect 198832 151512 198884 151564
rect 212448 151512 212500 151564
rect 280988 151512 281040 151564
rect 97908 151444 97960 151496
rect 193680 151444 193732 151496
rect 202788 151444 202840 151496
rect 273260 151444 273312 151496
rect 92388 151376 92440 151428
rect 188528 151376 188580 151428
rect 195888 151376 195940 151428
rect 268200 151376 268252 151428
rect 78588 151308 78640 151360
rect 178316 151308 178368 151360
rect 180708 151308 180760 151360
rect 256608 151308 256660 151360
rect 64788 151240 64840 151292
rect 57888 151172 57940 151224
rect 162860 151172 162912 151224
rect 167644 151240 167696 151292
rect 245016 151240 245068 151292
rect 168012 151172 168064 151224
rect 168104 151172 168156 151224
rect 246304 151172 246356 151224
rect 50988 151104 51040 151156
rect 157708 151104 157760 151156
rect 158628 151104 158680 151156
rect 239956 151104 240008 151156
rect 38568 151036 38620 151088
rect 147496 151036 147548 151088
rect 151728 151036 151780 151088
rect 234804 151036 234856 151088
rect 146208 150968 146260 151020
rect 229652 150968 229704 151020
rect 153108 150900 153160 150952
rect 235448 150900 235500 150952
rect 166908 150832 166960 150884
rect 168104 150832 168156 150884
rect 98920 150560 98972 150612
rect 114468 150560 114520 150612
rect 92020 150492 92072 150544
rect 114100 150492 114152 150544
rect 85212 150424 85264 150476
rect 116308 150424 116360 150476
rect 127072 150152 127124 150204
rect 128222 150152 128274 150204
rect 132500 150152 132552 150204
rect 133374 150152 133426 150204
rect 139400 150152 139452 150204
rect 140458 150152 140510 150204
rect 145104 150152 145156 150204
rect 146254 150152 146306 150204
rect 147680 150152 147732 150204
rect 148830 150152 148882 150204
rect 149152 150152 149204 150204
rect 150026 150152 150078 150204
rect 150532 150152 150584 150204
rect 151314 150152 151366 150204
rect 154672 150152 154724 150204
rect 155822 150152 155874 150204
rect 160100 150152 160152 150204
rect 160974 150152 161026 150204
rect 161480 150152 161532 150204
rect 162262 150152 162314 150204
rect 163044 150152 163096 150204
rect 164194 150152 164246 150204
rect 168380 150152 168432 150204
rect 169346 150152 169398 150204
rect 169760 150152 169812 150204
rect 170634 150152 170686 150204
rect 171140 150152 171192 150204
rect 171922 150152 171974 150204
rect 172704 150152 172756 150204
rect 173854 150152 173906 150204
rect 180984 150152 181036 150204
rect 182134 150152 182186 150204
rect 183560 150152 183612 150204
rect 184710 150152 184762 150204
rect 190736 150152 190788 150204
rect 191794 150152 191846 150204
rect 200304 150152 200356 150204
rect 201454 150152 201506 150204
rect 201592 150152 201644 150204
rect 202742 150152 202794 150204
rect 207020 150152 207072 150204
rect 207894 150152 207946 150204
rect 209964 150152 210016 150204
rect 211114 150152 211166 150204
rect 215392 150152 215444 150204
rect 216174 150152 216226 150204
rect 224960 150152 225012 150204
rect 225834 150152 225886 150204
rect 229192 150152 229244 150204
rect 230342 150152 230394 150204
rect 231952 150152 232004 150204
rect 232918 150152 232970 150204
rect 233240 150152 233292 150204
rect 234206 150152 234258 150204
rect 242900 150152 242952 150204
rect 243774 150152 243826 150204
rect 247132 150152 247184 150204
rect 248282 150152 248334 150204
rect 252560 150152 252612 150204
rect 253434 150152 253486 150204
rect 258080 150152 258132 150204
rect 259230 150152 259282 150204
rect 260840 150152 260892 150204
rect 261806 150152 261858 150204
rect 263600 150152 263652 150204
rect 264382 150152 264434 150204
rect 265164 150152 265216 150204
rect 266314 150152 266366 150204
rect 273444 150152 273496 150204
rect 274594 150152 274646 150204
rect 276020 150152 276072 150204
rect 277170 150152 277222 150204
rect 278780 150152 278832 150204
rect 279746 150152 279798 150204
rect 283104 150152 283156 150204
rect 284254 150152 284306 150204
rect 291200 150152 291252 150204
rect 291982 150152 292034 150204
rect 292764 150152 292816 150204
rect 293914 150152 293966 150204
rect 294052 150152 294104 150204
rect 295202 150152 295254 150204
rect 310612 150152 310664 150204
rect 311854 150152 311906 150204
rect 311992 150152 312044 150204
rect 313142 150152 313194 150204
rect 331312 150152 331364 150204
rect 332462 150152 332514 150204
rect 339592 150152 339644 150204
rect 340742 150152 340794 150204
rect 349252 150152 349304 150204
rect 350402 150152 350454 150204
rect 350540 150152 350592 150204
rect 351690 150152 351742 150204
rect 351920 150152 351972 150204
rect 352978 150152 353030 150204
rect 357624 150152 357676 150204
rect 358774 150152 358826 150204
rect 360200 150152 360252 150204
rect 361350 150152 361402 150204
rect 361580 150152 361632 150204
rect 362638 150152 362690 150204
rect 365904 150152 365956 150204
rect 367054 150152 367106 150204
rect 380900 150152 380952 150204
rect 381866 150152 381918 150204
rect 382280 150152 382332 150204
rect 383154 150152 383206 150204
rect 385224 150152 385276 150204
rect 386374 150152 386426 150204
rect 386512 150152 386564 150204
rect 387662 150152 387714 150204
rect 391940 150152 391992 150204
rect 392814 150152 392866 150204
rect 396172 150152 396224 150204
rect 397230 150152 397282 150204
rect 400220 150152 400272 150204
rect 401094 150152 401146 150204
rect 412824 150152 412876 150204
rect 413974 150152 414026 150204
rect 423772 150152 423824 150204
rect 424922 150152 424974 150204
rect 434720 150152 434772 150204
rect 435778 150152 435830 150204
rect 441712 150152 441764 150204
rect 442862 150152 442914 150204
rect 443000 150152 443052 150204
rect 444150 150152 444202 150204
rect 444380 150152 444432 150204
rect 445438 150152 445490 150204
rect 456800 150152 456852 150204
rect 457674 150152 457726 150204
rect 458364 150152 458416 150204
rect 459514 150152 459566 150204
rect 477684 150152 477736 150204
rect 478834 150152 478886 150204
rect 478972 150152 479024 150204
rect 480122 150152 480174 150204
rect 480260 150152 480312 150204
rect 481410 150152 481462 150204
rect 481640 150152 481692 150204
rect 482698 150152 482750 150204
rect 97724 149880 97776 149932
rect 117228 149880 117280 149932
rect 89168 149812 89220 149864
rect 117136 149812 117188 149864
rect 78588 149744 78640 149796
rect 112812 149744 112864 149796
rect 71688 149676 71740 149728
rect 109684 149676 109736 149728
rect 75184 149608 75236 149660
rect 114284 149608 114336 149660
rect 68376 149540 68428 149592
rect 112720 149540 112772 149592
rect 64696 149472 64748 149524
rect 111340 149472 111392 149524
rect 61384 149404 61436 149456
rect 112628 149404 112680 149456
rect 57888 149336 57940 149388
rect 112536 149336 112588 149388
rect 44088 149268 44140 149320
rect 47584 149268 47636 149320
rect 50988 149268 51040 149320
rect 54576 149268 54628 149320
rect 111248 149268 111300 149320
rect 112444 149200 112496 149252
rect 111156 149132 111208 149184
rect 111064 149064 111116 149116
rect 109592 148996 109644 149048
rect 116124 148996 116176 149048
rect 111800 147568 111852 147620
rect 116124 147568 116176 147620
rect 109960 147092 110012 147144
rect 116032 147092 116084 147144
rect 110328 147024 110380 147076
rect 116400 147024 116452 147076
rect 110052 146956 110104 147008
rect 116768 146956 116820 147008
rect 110144 146888 110196 146940
rect 116860 146888 116912 146940
rect 110236 145528 110288 145580
rect 117044 145528 117096 145580
rect 113732 143556 113784 143608
rect 115204 143556 115256 143608
rect 114468 143488 114520 143540
rect 116124 143488 116176 143540
rect 114376 141720 114428 141772
rect 116492 141720 116544 141772
rect 114100 140700 114152 140752
rect 116492 140700 116544 140752
rect 112812 132404 112864 132456
rect 116124 132404 116176 132456
rect 114284 131044 114336 131096
rect 115940 131044 115992 131096
rect 109684 128256 109736 128308
rect 116124 128256 116176 128308
rect 112720 126896 112772 126948
rect 116124 126896 116176 126948
rect 111340 124108 111392 124160
rect 116124 124108 116176 124160
rect 112628 122748 112680 122800
rect 115940 122748 115992 122800
rect 112536 121388 112588 121440
rect 116124 121388 116176 121440
rect 114284 118736 114336 118788
rect 115296 118736 115348 118788
rect 111248 118600 111300 118652
rect 116124 118600 116176 118652
rect 112444 117240 112496 117292
rect 116124 117240 116176 117292
rect 111156 114452 111208 114504
rect 116124 114452 116176 114504
rect 111064 113092 111116 113144
rect 116124 113092 116176 113144
rect 113548 109624 113600 109676
rect 115388 109624 115440 109676
rect 114192 104796 114244 104848
rect 115940 104796 115992 104848
rect 114008 99288 114060 99340
rect 116492 99288 116544 99340
rect 114468 96840 114520 96892
rect 116768 96840 116820 96892
rect 113824 93576 113876 93628
rect 116492 93576 116544 93628
rect 113916 92420 113968 92472
rect 116124 92420 116176 92472
rect 115204 91604 115256 91656
rect 116860 91604 116912 91656
rect 114468 87184 114520 87236
rect 116676 87184 116728 87236
rect 114100 86912 114152 86964
rect 116216 86912 116268 86964
rect 113916 71748 113968 71800
rect 116492 71748 116544 71800
rect 114100 69028 114152 69080
rect 116308 69028 116360 69080
rect 114192 67600 114244 67652
rect 116216 67600 116268 67652
rect 113548 64744 113600 64796
rect 116584 64744 116636 64796
rect 112444 62092 112496 62144
rect 116124 62092 116176 62144
rect 113824 52436 113876 52488
rect 116400 52436 116452 52488
rect 113916 48288 113968 48340
rect 115940 48288 115992 48340
rect 111064 46928 111116 46980
rect 116032 46928 116084 46980
rect 113640 44140 113692 44192
rect 117136 44140 117188 44192
rect 114008 41420 114060 41472
rect 115940 41420 115992 41472
rect 114100 38632 114152 38684
rect 115940 38632 115992 38684
rect 114284 37272 114336 37324
rect 116400 37272 116452 37324
rect 114376 34484 114428 34536
rect 115940 34484 115992 34536
rect 113732 33124 113784 33176
rect 116400 33124 116452 33176
rect 114468 31764 114520 31816
rect 115940 31764 115992 31816
rect 111156 28976 111208 29028
rect 116124 28976 116176 29028
rect 111248 27616 111300 27668
rect 116124 27616 116176 27668
rect 112536 24828 112588 24880
rect 116124 24828 116176 24880
rect 114192 22108 114244 22160
rect 115940 22108 115992 22160
rect 111340 19320 111392 19372
rect 116124 19320 116176 19372
rect 113548 13812 113600 13864
rect 116216 13812 116268 13864
rect 113640 8236 113692 8288
rect 115204 8236 115256 8288
rect 109684 4904 109736 4956
rect 116492 4904 116544 4956
rect 109868 4836 109920 4888
rect 116400 4836 116452 4888
rect 109776 4768 109828 4820
rect 117136 4768 117188 4820
rect 109592 4496 109644 4548
rect 112444 4496 112496 4548
rect 109960 4156 110012 4208
rect 116124 4156 116176 4208
rect 110052 2932 110104 2984
rect 32496 2592 32548 2644
rect 98276 2592 98328 2644
rect 110420 2864 110472 2916
rect 106188 2320 106240 2372
rect 116584 2320 116636 2372
rect 102968 2252 103020 2304
rect 116676 2252 116728 2304
rect 99656 2184 99708 2236
rect 116768 2184 116820 2236
rect 96344 2116 96396 2168
rect 116860 2116 116912 2168
rect 89628 2048 89680 2100
rect 116952 2048 117004 2100
rect 82728 1980 82780 2032
rect 111064 1980 111116 2032
rect 76012 1912 76064 1964
rect 109776 1912 109828 1964
rect 62672 1844 62724 1896
rect 114376 1844 114428 1896
rect 491300 1844 491352 1896
rect 493922 1844 493974 1896
rect 59360 1776 59412 1828
rect 113732 1776 113784 1828
rect 49332 1708 49384 1760
rect 111156 1708 111208 1760
rect 46020 1640 46072 1692
rect 111248 1640 111300 1692
rect 35992 1572 36044 1624
rect 114192 1572 114244 1624
rect 39304 1504 39356 1556
rect 117228 1504 117280 1556
rect 15936 1436 15988 1488
rect 98644 1436 98696 1488
rect 110052 1436 110104 1488
rect 143632 1436 143684 1488
rect 12624 1368 12676 1420
rect 100760 1368 100812 1420
rect 110420 1368 110472 1420
rect 193588 1368 193640 1420
rect 92664 1300 92716 1352
rect 113824 1300 113876 1352
rect 22652 1232 22704 1284
rect 113640 1232 113692 1284
rect 42616 1164 42668 1216
rect 112536 1164 112588 1216
rect 52644 1096 52696 1148
rect 114468 1096 114520 1148
rect 65984 1028 66036 1080
rect 114284 1028 114336 1080
rect 69296 960 69348 1012
rect 114100 960 114152 1012
rect 72700 892 72752 944
rect 114008 892 114060 944
rect 79324 824 79376 876
rect 117044 824 117096 876
rect 86040 756 86092 808
rect 113916 756 113968 808
rect 2688 688 2740 740
rect 116124 688 116176 740
<< metal2 >>
rect 386 163200 442 164400
rect 1214 163200 1270 164400
rect 2042 163200 2098 164400
rect 2870 163200 2926 164400
rect 3698 163200 3754 164400
rect 3804 163254 4108 163282
rect 400 158778 428 163200
rect 388 158772 440 158778
rect 388 158714 440 158720
rect 1228 155242 1256 163200
rect 2056 161474 2084 163200
rect 2056 161446 2176 161474
rect 2044 158772 2096 158778
rect 2044 158714 2096 158720
rect 1216 155236 1268 155242
rect 1216 155178 1268 155184
rect 2056 151065 2084 158714
rect 2148 158030 2176 161446
rect 2136 158024 2188 158030
rect 2136 157966 2188 157972
rect 2884 155378 2912 163200
rect 3712 163146 3740 163200
rect 3804 163146 3832 163254
rect 3712 163118 3832 163146
rect 2872 155372 2924 155378
rect 2872 155314 2924 155320
rect 4080 153882 4108 163254
rect 4526 163200 4582 164400
rect 5354 163200 5410 164400
rect 6274 163200 6330 164400
rect 7102 163200 7158 164400
rect 7930 163200 7986 164400
rect 8758 163200 8814 164400
rect 9586 163200 9642 164400
rect 10414 163200 10470 164400
rect 11242 163200 11298 164400
rect 12162 163200 12218 164400
rect 12990 163200 13046 164400
rect 13818 163200 13874 164400
rect 14646 163200 14702 164400
rect 15474 163200 15530 164400
rect 16302 163200 16358 164400
rect 17130 163200 17186 164400
rect 18050 163200 18106 164400
rect 18878 163200 18934 164400
rect 19706 163200 19762 164400
rect 20534 163200 20590 164400
rect 21362 163200 21418 164400
rect 22190 163200 22246 164400
rect 23018 163200 23074 164400
rect 23124 163254 23428 163282
rect 4540 157214 4568 163200
rect 4528 157208 4580 157214
rect 4528 157150 4580 157156
rect 5368 155310 5396 163200
rect 5356 155304 5408 155310
rect 5356 155246 5408 155252
rect 4068 153876 4120 153882
rect 4068 153818 4120 153824
rect 6288 152522 6316 163200
rect 7116 153785 7144 163200
rect 7944 156641 7972 163200
rect 7930 156632 7986 156641
rect 7930 156567 7986 156576
rect 8772 155446 8800 163200
rect 8760 155440 8812 155446
rect 8760 155382 8812 155388
rect 7102 153776 7158 153785
rect 7102 153711 7158 153720
rect 6276 152516 6328 152522
rect 6276 152458 6328 152464
rect 9600 152425 9628 163200
rect 10428 153921 10456 163200
rect 11256 156738 11284 163200
rect 12176 158001 12204 163200
rect 13004 159390 13032 163200
rect 12992 159384 13044 159390
rect 12992 159326 13044 159332
rect 12162 157992 12218 158001
rect 12162 157927 12218 157936
rect 11244 156732 11296 156738
rect 11244 156674 11296 156680
rect 13832 154086 13860 163200
rect 14660 156670 14688 163200
rect 14648 156664 14700 156670
rect 14648 156606 14700 156612
rect 15488 155514 15516 163200
rect 15476 155508 15528 155514
rect 15476 155450 15528 155456
rect 13820 154080 13872 154086
rect 13820 154022 13872 154028
rect 10414 153912 10470 153921
rect 10414 153847 10470 153856
rect 16316 152561 16344 163200
rect 17144 153950 17172 163200
rect 18064 156806 18092 163200
rect 18892 158098 18920 163200
rect 19720 159361 19748 163200
rect 19706 159352 19762 159361
rect 19706 159287 19762 159296
rect 18880 158092 18932 158098
rect 18880 158034 18932 158040
rect 18052 156800 18104 156806
rect 18052 156742 18104 156748
rect 20548 154018 20576 163200
rect 21376 156874 21404 163200
rect 21364 156868 21416 156874
rect 21364 156810 21416 156816
rect 22204 155582 22232 163200
rect 23032 163146 23060 163200
rect 23124 163146 23152 163254
rect 23032 163118 23152 163146
rect 22192 155576 22244 155582
rect 22192 155518 22244 155524
rect 20536 154012 20588 154018
rect 20536 153954 20588 153960
rect 17132 153944 17184 153950
rect 17132 153886 17184 153892
rect 23400 152590 23428 163254
rect 23938 163200 23994 164400
rect 24766 163200 24822 164400
rect 25594 163200 25650 164400
rect 26422 163200 26478 164400
rect 27250 163200 27306 164400
rect 28078 163200 28134 164400
rect 28906 163200 28962 164400
rect 29826 163200 29882 164400
rect 30654 163200 30710 164400
rect 31482 163200 31538 164400
rect 32310 163200 32366 164400
rect 33138 163200 33194 164400
rect 33966 163200 34022 164400
rect 34072 163254 34468 163282
rect 23952 155650 23980 163200
rect 24780 156942 24808 163200
rect 24768 156936 24820 156942
rect 24768 156878 24820 156884
rect 23940 155644 23992 155650
rect 23940 155586 23992 155592
rect 25608 154154 25636 163200
rect 26436 159458 26464 163200
rect 26424 159452 26476 159458
rect 26424 159394 26476 159400
rect 27264 155281 27292 163200
rect 28092 156777 28120 163200
rect 28078 156768 28134 156777
rect 28078 156703 28134 156712
rect 27250 155272 27306 155281
rect 27250 155207 27306 155216
rect 25596 154148 25648 154154
rect 25596 154090 25648 154096
rect 23388 152584 23440 152590
rect 16302 152552 16358 152561
rect 23388 152526 23440 152532
rect 16302 152487 16358 152496
rect 9586 152416 9642 152425
rect 9586 152351 9642 152360
rect 23294 152280 23350 152289
rect 23294 152215 23350 152224
rect 12990 152144 13046 152153
rect 12990 152079 13046 152088
rect 9494 152008 9550 152017
rect 9494 151943 9550 151952
rect 2686 151872 2742 151881
rect 2686 151807 2742 151816
rect 2042 151056 2098 151065
rect 2042 150991 2098 151000
rect 2700 149940 2728 151807
rect 9508 149940 9536 151943
rect 13004 149940 13032 152079
rect 19798 150512 19854 150521
rect 19798 150447 19854 150456
rect 19812 149940 19840 150447
rect 23308 149940 23336 152215
rect 26700 152176 26752 152182
rect 26700 152118 26752 152124
rect 26712 149940 26740 152118
rect 28920 151201 28948 163200
rect 29840 152697 29868 163200
rect 30668 155417 30696 163200
rect 31496 158234 31524 163200
rect 31484 158228 31536 158234
rect 31484 158170 31536 158176
rect 32324 158137 32352 163200
rect 33152 159497 33180 163200
rect 33980 163146 34008 163200
rect 34072 163146 34100 163254
rect 33980 163118 34100 163146
rect 33138 159488 33194 159497
rect 33138 159423 33194 159432
rect 32310 158128 32366 158137
rect 32310 158063 32366 158072
rect 30654 155408 30710 155417
rect 30654 155343 30710 155352
rect 29826 152688 29882 152697
rect 34440 152658 34468 163254
rect 34794 163200 34850 164400
rect 35714 163200 35770 164400
rect 36542 163200 36598 164400
rect 37370 163200 37426 164400
rect 38198 163200 38254 164400
rect 38304 163254 38516 163282
rect 34808 154222 34836 163200
rect 35728 158166 35756 163200
rect 36556 160750 36584 163200
rect 36544 160744 36596 160750
rect 36544 160686 36596 160692
rect 37384 159118 37412 163200
rect 38212 163146 38240 163200
rect 38304 163146 38332 163254
rect 38212 163118 38332 163146
rect 37372 159112 37424 159118
rect 37372 159054 37424 159060
rect 35716 158160 35768 158166
rect 35716 158102 35768 158108
rect 34796 154216 34848 154222
rect 34796 154158 34848 154164
rect 38488 154057 38516 163254
rect 39026 163200 39082 164400
rect 39854 163200 39910 164400
rect 40682 163200 40738 164400
rect 41602 163200 41658 164400
rect 42430 163200 42486 164400
rect 43258 163200 43314 164400
rect 44086 163200 44142 164400
rect 44914 163200 44970 164400
rect 45742 163200 45798 164400
rect 46570 163200 46626 164400
rect 47490 163200 47546 164400
rect 48318 163200 48374 164400
rect 49146 163200 49202 164400
rect 49974 163200 50030 164400
rect 50802 163200 50858 164400
rect 51630 163200 51686 164400
rect 52458 163200 52514 164400
rect 53378 163200 53434 164400
rect 54206 163200 54262 164400
rect 55034 163200 55090 164400
rect 55862 163200 55918 164400
rect 56690 163200 56746 164400
rect 57518 163200 57574 164400
rect 57624 163254 57928 163282
rect 38568 159112 38620 159118
rect 38568 159054 38620 159060
rect 38474 154048 38530 154057
rect 38474 153983 38530 153992
rect 29826 152623 29882 152632
rect 34428 152652 34480 152658
rect 34428 152594 34480 152600
rect 33600 151904 33652 151910
rect 33600 151846 33652 151852
rect 28906 151192 28962 151201
rect 28906 151127 28962 151136
rect 33612 149940 33640 151846
rect 38580 151094 38608 159054
rect 39040 157010 39068 163200
rect 39868 162586 39896 163200
rect 39856 162580 39908 162586
rect 39856 162522 39908 162528
rect 40696 160818 40724 163200
rect 40684 160812 40736 160818
rect 40684 160754 40736 160760
rect 39028 157004 39080 157010
rect 39028 156946 39080 156952
rect 41616 155718 41644 163200
rect 42444 158273 42472 163200
rect 43272 162654 43300 163200
rect 43260 162648 43312 162654
rect 43260 162590 43312 162596
rect 42430 158264 42486 158273
rect 42430 158199 42486 158208
rect 41604 155712 41656 155718
rect 41604 155654 41656 155660
rect 40500 152040 40552 152046
rect 40500 151982 40552 151988
rect 38568 151088 38620 151094
rect 38568 151030 38620 151036
rect 37002 150648 37058 150657
rect 37002 150583 37058 150592
rect 37016 149940 37044 150583
rect 40512 149940 40540 151982
rect 44100 151337 44128 163200
rect 44928 154290 44956 163200
rect 45756 158302 45784 163200
rect 46584 159730 46612 163200
rect 47504 160886 47532 163200
rect 47492 160880 47544 160886
rect 47492 160822 47544 160828
rect 46572 159724 46624 159730
rect 46572 159666 46624 159672
rect 45744 158296 45796 158302
rect 45744 158238 45796 158244
rect 48332 155786 48360 163200
rect 49160 157078 49188 163200
rect 49988 160070 50016 163200
rect 50816 161474 50844 163200
rect 50816 161446 51028 161474
rect 49976 160064 50028 160070
rect 49976 160006 50028 160012
rect 49148 157072 49200 157078
rect 49148 157014 49200 157020
rect 48320 155780 48372 155786
rect 48320 155722 48372 155728
rect 44916 154284 44968 154290
rect 44916 154226 44968 154232
rect 44086 151328 44142 151337
rect 44086 151263 44142 151272
rect 51000 151162 51028 161446
rect 51644 154358 51672 163200
rect 52472 158370 52500 163200
rect 53392 159662 53420 163200
rect 54220 160954 54248 163200
rect 54208 160948 54260 160954
rect 54208 160890 54260 160896
rect 53380 159656 53432 159662
rect 53380 159598 53432 159604
rect 52460 158364 52512 158370
rect 52460 158306 52512 158312
rect 55048 155854 55076 163200
rect 55876 157146 55904 163200
rect 56704 161634 56732 163200
rect 57532 163146 57560 163200
rect 57624 163146 57652 163254
rect 57532 163118 57652 163146
rect 56692 161628 56744 161634
rect 56692 161570 56744 161576
rect 55864 157140 55916 157146
rect 55864 157082 55916 157088
rect 55036 155848 55088 155854
rect 55036 155790 55088 155796
rect 51632 154352 51684 154358
rect 51632 154294 51684 154300
rect 57900 151230 57928 163254
rect 58346 163200 58402 164400
rect 59266 163200 59322 164400
rect 60094 163200 60150 164400
rect 60922 163200 60978 164400
rect 61750 163200 61806 164400
rect 62578 163200 62634 164400
rect 63406 163200 63462 164400
rect 64234 163200 64290 164400
rect 65154 163200 65210 164400
rect 65982 163200 66038 164400
rect 66810 163200 66866 164400
rect 67638 163200 67694 164400
rect 68466 163200 68522 164400
rect 69294 163200 69350 164400
rect 70122 163200 70178 164400
rect 71042 163200 71098 164400
rect 71870 163200 71926 164400
rect 72698 163200 72754 164400
rect 73526 163200 73582 164400
rect 74354 163200 74410 164400
rect 75182 163200 75238 164400
rect 76010 163200 76066 164400
rect 76930 163200 76986 164400
rect 77758 163200 77814 164400
rect 78586 163200 78642 164400
rect 79414 163200 79470 164400
rect 80242 163200 80298 164400
rect 81070 163200 81126 164400
rect 81898 163200 81954 164400
rect 82818 163200 82874 164400
rect 83646 163200 83702 164400
rect 83752 163254 84148 163282
rect 58360 154426 58388 163200
rect 59280 158438 59308 163200
rect 60108 159798 60136 163200
rect 60936 161022 60964 163200
rect 61764 161702 61792 163200
rect 61752 161696 61804 161702
rect 61752 161638 61804 161644
rect 60924 161016 60976 161022
rect 60924 160958 60976 160964
rect 60096 159792 60148 159798
rect 60096 159734 60148 159740
rect 62592 158574 62620 163200
rect 62580 158568 62632 158574
rect 62580 158510 62632 158516
rect 59268 158432 59320 158438
rect 59268 158374 59320 158380
rect 58348 154420 58400 154426
rect 58348 154362 58400 154368
rect 63420 153746 63448 163200
rect 64248 158778 64276 163200
rect 65168 161838 65196 163200
rect 65156 161832 65208 161838
rect 65156 161774 65208 161780
rect 64236 158772 64288 158778
rect 64236 158714 64288 158720
rect 64788 158772 64840 158778
rect 64788 158714 64840 158720
rect 63408 153740 63460 153746
rect 63408 153682 63460 153688
rect 64800 151298 64828 158714
rect 65996 158506 66024 163200
rect 66824 160002 66852 163200
rect 67652 161090 67680 163200
rect 68480 161770 68508 163200
rect 68468 161764 68520 161770
rect 68468 161706 68520 161712
rect 67640 161084 67692 161090
rect 67640 161026 67692 161032
rect 66812 159996 66864 160002
rect 66812 159938 66864 159944
rect 65984 158500 66036 158506
rect 65984 158442 66036 158448
rect 69308 157282 69336 163200
rect 70136 159633 70164 163200
rect 70122 159624 70178 159633
rect 70122 159559 70178 159568
rect 71056 158778 71084 163200
rect 71884 162042 71912 163200
rect 71872 162036 71924 162042
rect 71872 161978 71924 161984
rect 71044 158772 71096 158778
rect 71044 158714 71096 158720
rect 71688 158772 71740 158778
rect 71688 158714 71740 158720
rect 69296 157276 69348 157282
rect 69296 157218 69348 157224
rect 71700 151473 71728 158714
rect 72712 155922 72740 163200
rect 72700 155916 72752 155922
rect 72700 155858 72752 155864
rect 73540 152726 73568 163200
rect 74368 160721 74396 163200
rect 75196 161906 75224 163200
rect 75184 161900 75236 161906
rect 75184 161842 75236 161848
rect 74354 160712 74410 160721
rect 74354 160647 74410 160656
rect 76024 157350 76052 163200
rect 76944 159934 76972 163200
rect 76932 159928 76984 159934
rect 76932 159870 76984 159876
rect 77772 158778 77800 163200
rect 78600 161974 78628 163200
rect 78588 161968 78640 161974
rect 78588 161910 78640 161916
rect 77760 158772 77812 158778
rect 77760 158714 77812 158720
rect 78588 158772 78640 158778
rect 78588 158714 78640 158720
rect 76012 157344 76064 157350
rect 76012 157286 76064 157292
rect 73528 152720 73580 152726
rect 73528 152662 73580 152668
rect 71686 151464 71742 151473
rect 71686 151399 71742 151408
rect 78600 151366 78628 158714
rect 79428 157826 79456 163200
rect 80256 159594 80284 163200
rect 81084 161158 81112 163200
rect 81912 162110 81940 163200
rect 81900 162104 81952 162110
rect 81900 162046 81952 162052
rect 81072 161152 81124 161158
rect 81072 161094 81124 161100
rect 80244 159588 80296 159594
rect 80244 159530 80296 159536
rect 79416 157820 79468 157826
rect 79416 157762 79468 157768
rect 82832 156913 82860 163200
rect 83660 163146 83688 163200
rect 83752 163146 83780 163254
rect 83660 163118 83780 163146
rect 82818 156904 82874 156913
rect 82818 156839 82874 156848
rect 84120 152794 84148 163254
rect 84474 163200 84530 164400
rect 85302 163200 85358 164400
rect 86130 163200 86186 164400
rect 86958 163200 87014 164400
rect 87786 163200 87842 164400
rect 88706 163200 88762 164400
rect 89534 163200 89590 164400
rect 90362 163200 90418 164400
rect 91190 163200 91246 164400
rect 92018 163200 92074 164400
rect 92846 163200 92902 164400
rect 93674 163200 93730 164400
rect 94594 163200 94650 164400
rect 95422 163200 95478 164400
rect 96250 163200 96306 164400
rect 97078 163200 97134 164400
rect 97906 163200 97962 164400
rect 98734 163200 98790 164400
rect 99562 163200 99618 164400
rect 100482 163200 100538 164400
rect 101310 163200 101366 164400
rect 102138 163200 102194 164400
rect 102966 163200 103022 164400
rect 103072 163254 103468 163282
rect 84488 158778 84516 163200
rect 84476 158772 84528 158778
rect 84476 158714 84528 158720
rect 85316 155553 85344 163200
rect 85488 158772 85540 158778
rect 85488 158714 85540 158720
rect 85302 155544 85358 155553
rect 85302 155479 85358 155488
rect 84108 152788 84160 152794
rect 84108 152730 84160 152736
rect 81716 151836 81768 151842
rect 81716 151778 81768 151784
rect 78588 151360 78640 151366
rect 78588 151302 78640 151308
rect 64788 151292 64840 151298
rect 64788 151234 64840 151240
rect 57888 151224 57940 151230
rect 57888 151166 57940 151172
rect 50988 151156 51040 151162
rect 50988 151098 51040 151104
rect 81728 149940 81756 151778
rect 85500 151609 85528 158714
rect 86144 158642 86172 163200
rect 86972 159866 87000 163200
rect 87800 160857 87828 163200
rect 88720 162178 88748 163200
rect 88708 162172 88760 162178
rect 88708 162114 88760 162120
rect 87786 160848 87842 160857
rect 87786 160783 87842 160792
rect 86960 159860 87012 159866
rect 86960 159802 87012 159808
rect 86132 158636 86184 158642
rect 86132 158578 86184 158584
rect 89548 155174 89576 163200
rect 89536 155168 89588 155174
rect 89536 155110 89588 155116
rect 90376 152862 90404 163200
rect 91204 159118 91232 163200
rect 92032 162246 92060 163200
rect 92020 162240 92072 162246
rect 92020 162182 92072 162188
rect 91192 159112 91244 159118
rect 91192 159054 91244 159060
rect 92388 159112 92440 159118
rect 92388 159054 92440 159060
rect 90364 152856 90416 152862
rect 90364 152798 90416 152804
rect 89168 152040 89220 152046
rect 89168 151982 89220 151988
rect 88616 151972 88668 151978
rect 88616 151914 88668 151920
rect 85486 151600 85542 151609
rect 85486 151535 85542 151544
rect 85212 150476 85264 150482
rect 85212 150418 85264 150424
rect 85224 149940 85252 150418
rect 88628 149940 88656 151914
rect 89180 149870 89208 151982
rect 92400 151434 92428 159054
rect 92860 154494 92888 163200
rect 93688 159322 93716 163200
rect 94608 161226 94636 163200
rect 95436 162382 95464 163200
rect 95424 162376 95476 162382
rect 95424 162318 95476 162324
rect 94596 161220 94648 161226
rect 94596 161162 94648 161168
rect 93676 159316 93728 159322
rect 93676 159258 93728 159264
rect 96264 156602 96292 163200
rect 96252 156596 96304 156602
rect 96252 156538 96304 156544
rect 92848 154488 92900 154494
rect 92848 154430 92900 154436
rect 97092 152930 97120 163200
rect 97080 152924 97132 152930
rect 97080 152866 97132 152872
rect 95516 152040 95568 152046
rect 95516 151982 95568 151988
rect 92388 151428 92440 151434
rect 92388 151370 92440 151376
rect 92020 150544 92072 150550
rect 92020 150486 92072 150492
rect 92032 149940 92060 150486
rect 95528 149940 95556 151982
rect 97724 151836 97776 151842
rect 97724 151778 97776 151784
rect 97736 149938 97764 151778
rect 97920 151502 97948 163200
rect 98748 162314 98776 163200
rect 98736 162308 98788 162314
rect 98736 162250 98788 162256
rect 99576 158710 99604 163200
rect 100496 159526 100524 163200
rect 101324 161294 101352 163200
rect 102152 162518 102180 163200
rect 102980 163146 103008 163200
rect 103072 163146 103100 163254
rect 102980 163118 103100 163146
rect 102140 162512 102192 162518
rect 102140 162454 102192 162460
rect 101312 161288 101364 161294
rect 101312 161230 101364 161236
rect 100484 159520 100536 159526
rect 100484 159462 100536 159468
rect 99564 158704 99616 158710
rect 99564 158646 99616 158652
rect 103440 154562 103468 163254
rect 103794 163200 103850 164400
rect 104622 163200 104678 164400
rect 105450 163200 105506 164400
rect 106370 163200 106426 164400
rect 107198 163200 107254 164400
rect 107304 163254 107516 163282
rect 103808 158778 103836 163200
rect 104636 161474 104664 163200
rect 104636 161446 104848 161474
rect 103796 158772 103848 158778
rect 103796 158714 103848 158720
rect 103428 154556 103480 154562
rect 103428 154498 103480 154504
rect 102324 152108 102376 152114
rect 102324 152050 102376 152056
rect 97908 151496 97960 151502
rect 97908 151438 97960 151444
rect 98920 150612 98972 150618
rect 98920 150554 98972 150560
rect 98932 149940 98960 150554
rect 102336 149940 102364 152050
rect 104820 151570 104848 161446
rect 105464 153814 105492 163200
rect 106384 157962 106412 163200
rect 107212 163146 107240 163200
rect 107304 163146 107332 163254
rect 107212 163118 107332 163146
rect 106372 157956 106424 157962
rect 106372 157898 106424 157904
rect 105452 153808 105504 153814
rect 105452 153750 105504 153756
rect 107488 152998 107516 163254
rect 108026 163200 108082 164400
rect 108854 163200 108910 164400
rect 109682 163200 109738 164400
rect 110510 163200 110566 164400
rect 111338 163200 111394 164400
rect 111444 163254 111748 163282
rect 108040 161362 108068 163200
rect 108868 162450 108896 163200
rect 108856 162444 108908 162450
rect 108856 162386 108908 162392
rect 108028 161356 108080 161362
rect 108028 161298 108080 161304
rect 109224 160064 109276 160070
rect 109224 160006 109276 160012
rect 109040 158772 109092 158778
rect 109040 158714 109092 158720
rect 109052 153202 109080 158714
rect 109132 157208 109184 157214
rect 109132 157150 109184 157156
rect 109040 153196 109092 153202
rect 109040 153138 109092 153144
rect 107476 152992 107528 152998
rect 107476 152934 107528 152940
rect 109144 152454 109172 157150
rect 109236 152833 109264 160006
rect 109696 159254 109724 163200
rect 109684 159248 109736 159254
rect 109684 159190 109736 159196
rect 110524 159186 110552 163200
rect 111352 163146 111380 163200
rect 111444 163146 111472 163254
rect 111352 163118 111472 163146
rect 110512 159180 110564 159186
rect 110512 159122 110564 159128
rect 109222 152824 109278 152833
rect 109222 152759 109278 152768
rect 109132 152448 109184 152454
rect 109132 152390 109184 152396
rect 110050 152280 110106 152289
rect 110050 152215 110106 152224
rect 109960 152108 110012 152114
rect 109960 152050 110012 152056
rect 105820 151836 105872 151842
rect 105740 151786 105820 151814
rect 104808 151564 104860 151570
rect 104808 151506 104860 151512
rect 105740 149954 105768 151786
rect 105820 151778 105872 151784
rect 106924 151836 106976 151842
rect 106924 151778 106976 151784
rect 97724 149932 97776 149938
rect 105740 149926 105846 149954
rect 97724 149874 97776 149880
rect 89168 149864 89220 149870
rect 78338 149802 78628 149818
rect 89168 149806 89220 149812
rect 78338 149796 78640 149802
rect 78338 149790 78588 149796
rect 78588 149738 78640 149744
rect 71688 149728 71740 149734
rect 71438 149676 71688 149682
rect 106936 149705 106964 151778
rect 109684 149728 109736 149734
rect 106922 149696 106978 149705
rect 71438 149670 71740 149676
rect 71438 149654 71728 149670
rect 74842 149666 75224 149682
rect 74842 149660 75236 149666
rect 74842 149654 75184 149660
rect 109684 149670 109736 149676
rect 106922 149631 106978 149640
rect 75184 149602 75236 149608
rect 68376 149592 68428 149598
rect 64538 149530 64736 149546
rect 68034 149540 68376 149546
rect 68034 149534 68428 149540
rect 64538 149524 64748 149530
rect 64538 149518 64696 149524
rect 68034 149518 68416 149534
rect 64696 149466 64748 149472
rect 61384 149456 61436 149462
rect 6366 149424 6422 149433
rect 6118 149382 6366 149410
rect 16486 149424 16542 149433
rect 16422 149382 16486 149410
rect 6366 149359 6422 149368
rect 30286 149424 30342 149433
rect 30222 149382 30286 149410
rect 16486 149359 16542 149368
rect 43930 149382 44128 149410
rect 47334 149382 47624 149410
rect 50830 149382 51028 149410
rect 54234 149382 54616 149410
rect 57730 149394 57928 149410
rect 61134 149404 61384 149410
rect 61134 149398 61436 149404
rect 57730 149388 57940 149394
rect 57730 149382 57888 149388
rect 30286 149359 30342 149368
rect 44100 149326 44128 149382
rect 47596 149326 47624 149382
rect 51000 149326 51028 149382
rect 54588 149326 54616 149382
rect 61134 149382 61424 149398
rect 109250 149382 109632 149410
rect 57888 149330 57940 149336
rect 44088 149320 44140 149326
rect 44088 149262 44140 149268
rect 47584 149320 47636 149326
rect 47584 149262 47636 149268
rect 50988 149320 51040 149326
rect 50988 149262 51040 149268
rect 54576 149320 54628 149326
rect 54576 149262 54628 149268
rect 109604 149054 109632 149382
rect 109592 149048 109644 149054
rect 109592 148990 109644 148996
rect 109696 128314 109724 149670
rect 109972 147150 110000 152050
rect 109960 147144 110012 147150
rect 109960 147086 110012 147092
rect 110064 147014 110092 152215
rect 110144 152176 110196 152182
rect 110144 152118 110196 152124
rect 110052 147008 110104 147014
rect 110052 146950 110104 146956
rect 110156 146946 110184 152118
rect 110328 151972 110380 151978
rect 110328 151914 110380 151920
rect 110236 151904 110288 151910
rect 110236 151846 110288 151852
rect 110144 146940 110196 146946
rect 110144 146882 110196 146888
rect 110248 145586 110276 151846
rect 110340 147082 110368 151914
rect 111720 151638 111748 163254
rect 112258 163200 112314 164400
rect 113086 163200 113142 164400
rect 113914 163200 113970 164400
rect 114742 163200 114798 164400
rect 115570 163200 115626 164400
rect 116398 163200 116454 164400
rect 117226 163200 117282 164400
rect 118146 163200 118202 164400
rect 118974 163200 119030 164400
rect 119802 163200 119858 164400
rect 120630 163200 120686 164400
rect 121458 163200 121514 164400
rect 122286 163200 122342 164400
rect 122392 163254 122696 163282
rect 112272 161498 112300 163200
rect 112260 161492 112312 161498
rect 112260 161434 112312 161440
rect 113100 157214 113128 163200
rect 113088 157208 113140 157214
rect 113088 157150 113140 157156
rect 113928 153066 113956 163200
rect 114756 161430 114784 163200
rect 115584 161566 115612 163200
rect 115572 161560 115624 161566
rect 115572 161502 115624 161508
rect 114744 161424 114796 161430
rect 114744 161366 114796 161372
rect 116412 156534 116440 163200
rect 116400 156528 116452 156534
rect 116400 156470 116452 156476
rect 117240 153134 117268 163200
rect 118160 154834 118188 163200
rect 118700 159248 118752 159254
rect 118700 159190 118752 159196
rect 118712 155106 118740 159190
rect 118988 158982 119016 163200
rect 118976 158976 119028 158982
rect 118976 158918 119028 158924
rect 118792 155236 118844 155242
rect 118792 155178 118844 155184
rect 118700 155100 118752 155106
rect 118700 155042 118752 155048
rect 118148 154828 118200 154834
rect 118148 154770 118200 154776
rect 118700 153740 118752 153746
rect 118700 153682 118752 153688
rect 117228 153128 117280 153134
rect 117228 153070 117280 153076
rect 113916 153060 113968 153066
rect 113916 153002 113968 153008
rect 118712 152386 118740 153682
rect 118700 152380 118752 152386
rect 118700 152322 118752 152328
rect 116214 152144 116270 152153
rect 116214 152079 116270 152088
rect 114376 152040 114428 152046
rect 113822 152008 113878 152017
rect 114376 151982 114428 151988
rect 113822 151943 113878 151952
rect 111708 151632 111760 151638
rect 111708 151574 111760 151580
rect 112812 149796 112864 149802
rect 112812 149738 112864 149744
rect 111798 149696 111854 149705
rect 111798 149631 111854 149640
rect 111340 149524 111392 149530
rect 111340 149466 111392 149472
rect 111248 149320 111300 149326
rect 111248 149262 111300 149268
rect 111156 149184 111208 149190
rect 111156 149126 111208 149132
rect 111064 149116 111116 149122
rect 111064 149058 111116 149064
rect 110328 147076 110380 147082
rect 110328 147018 110380 147024
rect 110236 145580 110288 145586
rect 110236 145522 110288 145528
rect 109684 128308 109736 128314
rect 109684 128250 109736 128256
rect 111076 113150 111104 149058
rect 111168 114510 111196 149126
rect 111260 118658 111288 149262
rect 111352 124166 111380 149466
rect 111812 147626 111840 149631
rect 112720 149592 112772 149598
rect 112720 149534 112772 149540
rect 112628 149456 112680 149462
rect 112628 149398 112680 149404
rect 112536 149388 112588 149394
rect 112536 149330 112588 149336
rect 112444 149252 112496 149258
rect 112444 149194 112496 149200
rect 111800 147620 111852 147626
rect 111800 147562 111852 147568
rect 111340 124160 111392 124166
rect 111340 124102 111392 124108
rect 111248 118652 111300 118658
rect 111248 118594 111300 118600
rect 112456 117298 112484 149194
rect 112548 121446 112576 149330
rect 112640 122806 112668 149398
rect 112732 126954 112760 149534
rect 112824 132462 112852 149738
rect 113730 144256 113786 144265
rect 113730 144191 113786 144200
rect 113744 143614 113772 144191
rect 113732 143608 113784 143614
rect 113732 143550 113784 143556
rect 112812 132456 112864 132462
rect 112812 132398 112864 132404
rect 112720 126948 112772 126954
rect 112720 126890 112772 126896
rect 112628 122800 112680 122806
rect 112628 122742 112680 122748
rect 112536 121440 112588 121446
rect 112536 121382 112588 121388
rect 112444 117292 112496 117298
rect 112444 117234 112496 117240
rect 111156 114504 111208 114510
rect 111156 114446 111208 114452
rect 111064 113144 111116 113150
rect 111064 113086 111116 113092
rect 113546 110120 113602 110129
rect 113546 110055 113602 110064
rect 113560 109682 113588 110055
rect 113548 109676 113600 109682
rect 113548 109618 113600 109624
rect 113836 93634 113864 151943
rect 114100 150544 114152 150550
rect 114006 150512 114062 150521
rect 114100 150486 114152 150492
rect 114006 150447 114062 150456
rect 113914 149152 113970 149161
rect 113914 149087 113970 149096
rect 113824 93628 113876 93634
rect 113824 93570 113876 93576
rect 113928 92478 113956 149087
rect 114020 99346 114048 150447
rect 114112 140758 114140 150486
rect 114284 149660 114336 149666
rect 114284 149602 114336 149608
rect 114190 149424 114246 149433
rect 114190 149359 114246 149368
rect 114100 140752 114152 140758
rect 114100 140694 114152 140700
rect 114098 132832 114154 132841
rect 114098 132767 114154 132776
rect 114008 99340 114060 99346
rect 114008 99282 114060 99288
rect 113916 92472 113968 92478
rect 113916 92414 113968 92420
rect 114112 86970 114140 132767
rect 114204 104854 114232 149359
rect 114296 131102 114324 149602
rect 114388 141778 114416 151982
rect 116228 151814 116256 152079
rect 118804 151814 118832 155178
rect 119816 153746 119844 163200
rect 120644 160070 120672 163200
rect 120632 160064 120684 160070
rect 120632 160006 120684 160012
rect 120172 159724 120224 159730
rect 120172 159666 120224 159672
rect 120080 158024 120132 158030
rect 120080 157966 120132 157972
rect 119804 153740 119856 153746
rect 119804 153682 119856 153688
rect 120092 151814 120120 157966
rect 120184 154970 120212 159666
rect 121472 158778 121500 163200
rect 122300 163146 122328 163200
rect 122392 163146 122420 163254
rect 122300 163118 122420 163146
rect 121460 158772 121512 158778
rect 121460 158714 121512 158720
rect 121092 155372 121144 155378
rect 121092 155314 121144 155320
rect 120172 154964 120224 154970
rect 120172 154906 120224 154912
rect 116228 151786 116716 151814
rect 118804 151786 119844 151814
rect 120092 151786 120488 151814
rect 114468 150612 114520 150618
rect 114468 150554 114520 150560
rect 114480 143546 114508 150554
rect 116308 150476 116360 150482
rect 116308 150418 116360 150424
rect 116124 149048 116176 149054
rect 116122 149016 116124 149025
rect 116176 149016 116178 149025
rect 116122 148951 116178 148960
rect 116124 147620 116176 147626
rect 116124 147562 116176 147568
rect 116032 147144 116084 147150
rect 116136 147121 116164 147562
rect 116032 147086 116084 147092
rect 116122 147112 116178 147121
rect 116044 145217 116072 147086
rect 116122 147047 116178 147056
rect 116030 145208 116086 145217
rect 116030 145143 116086 145152
rect 115204 143608 115256 143614
rect 115204 143550 115256 143556
rect 114468 143540 114520 143546
rect 114468 143482 114520 143488
rect 114376 141772 114428 141778
rect 114376 141714 114428 141720
rect 114284 131096 114336 131102
rect 114284 131038 114336 131044
rect 114282 121408 114338 121417
rect 114282 121343 114338 121352
rect 114296 118794 114324 121343
rect 114284 118788 114336 118794
rect 114284 118730 114336 118736
rect 114192 104848 114244 104854
rect 114192 104790 114244 104796
rect 114466 98696 114522 98705
rect 114466 98631 114522 98640
rect 114480 96898 114508 98631
rect 114468 96892 114520 96898
rect 114468 96834 114520 96840
rect 115216 91662 115244 143550
rect 116124 143540 116176 143546
rect 116124 143482 116176 143488
rect 116136 143313 116164 143482
rect 116122 143304 116178 143313
rect 116122 143239 116178 143248
rect 116320 135561 116348 150418
rect 116582 149288 116638 149297
rect 116582 149223 116638 149232
rect 116400 147076 116452 147082
rect 116400 147018 116452 147024
rect 116412 137601 116440 147018
rect 116492 141772 116544 141778
rect 116492 141714 116544 141720
rect 116504 141409 116532 141714
rect 116490 141400 116546 141409
rect 116490 141335 116546 141344
rect 116492 140752 116544 140758
rect 116492 140694 116544 140700
rect 116504 139505 116532 140694
rect 116490 139496 116546 139505
rect 116490 139431 116546 139440
rect 116398 137592 116454 137601
rect 116398 137527 116454 137536
rect 116306 135552 116362 135561
rect 116306 135487 116362 135496
rect 116124 132456 116176 132462
rect 116124 132398 116176 132404
rect 116136 131753 116164 132398
rect 116122 131744 116178 131753
rect 116122 131679 116178 131688
rect 115940 131096 115992 131102
rect 115940 131038 115992 131044
rect 115952 129849 115980 131038
rect 115938 129840 115994 129849
rect 115938 129775 115994 129784
rect 116124 128308 116176 128314
rect 116124 128250 116176 128256
rect 116136 127945 116164 128250
rect 116122 127936 116178 127945
rect 116122 127871 116178 127880
rect 116124 126948 116176 126954
rect 116124 126890 116176 126896
rect 116136 126041 116164 126890
rect 116122 126032 116178 126041
rect 116122 125967 116178 125976
rect 116124 124160 116176 124166
rect 116122 124128 116124 124137
rect 116176 124128 116178 124137
rect 116122 124063 116178 124072
rect 115940 122800 115992 122806
rect 115940 122742 115992 122748
rect 115952 122233 115980 122742
rect 115938 122224 115994 122233
rect 115938 122159 115994 122168
rect 116124 121440 116176 121446
rect 116124 121382 116176 121388
rect 116136 120193 116164 121382
rect 116122 120184 116178 120193
rect 116122 120119 116178 120128
rect 115296 118788 115348 118794
rect 115296 118730 115348 118736
rect 115204 91656 115256 91662
rect 115204 91598 115256 91604
rect 114466 87272 114522 87281
rect 114466 87207 114468 87216
rect 114520 87207 114522 87216
rect 114468 87178 114520 87184
rect 114100 86964 114152 86970
rect 114100 86906 114152 86912
rect 115308 83745 115336 118730
rect 116124 118652 116176 118658
rect 116124 118594 116176 118600
rect 116136 118289 116164 118594
rect 116122 118280 116178 118289
rect 116122 118215 116178 118224
rect 116124 117292 116176 117298
rect 116124 117234 116176 117240
rect 116136 116385 116164 117234
rect 116122 116376 116178 116385
rect 116122 116311 116178 116320
rect 116124 114504 116176 114510
rect 116122 114472 116124 114481
rect 116176 114472 116178 114481
rect 116122 114407 116178 114416
rect 116124 113144 116176 113150
rect 116124 113086 116176 113092
rect 116136 112577 116164 113086
rect 116122 112568 116178 112577
rect 116122 112503 116178 112512
rect 115388 109676 115440 109682
rect 115388 109618 115440 109624
rect 115294 83736 115350 83745
rect 115294 83671 115350 83680
rect 115400 81841 115428 109618
rect 115940 104848 115992 104854
rect 115938 104816 115940 104825
rect 115992 104816 115994 104825
rect 115938 104751 115994 104760
rect 116492 99340 116544 99346
rect 116492 99282 116544 99288
rect 116504 99113 116532 99282
rect 116490 99104 116546 99113
rect 116490 99039 116546 99048
rect 116596 97209 116624 149223
rect 116582 97200 116638 97209
rect 116582 97135 116638 97144
rect 116688 95305 116716 151786
rect 118974 151056 119030 151065
rect 118974 150991 119030 151000
rect 116950 150648 117006 150657
rect 116950 150583 117006 150592
rect 116768 147008 116820 147014
rect 116768 146950 116820 146956
rect 116780 101017 116808 146950
rect 116860 146940 116912 146946
rect 116860 146882 116912 146888
rect 116872 102921 116900 146882
rect 116964 108769 116992 150583
rect 118988 149954 119016 150991
rect 119816 150226 119844 151786
rect 120460 150226 120488 151786
rect 121104 150226 121132 155314
rect 122668 153882 122696 163254
rect 123114 163200 123170 164400
rect 124034 163200 124090 164400
rect 124862 163200 124918 164400
rect 125690 163200 125746 164400
rect 126518 163200 126574 164400
rect 127346 163200 127402 164400
rect 128174 163200 128230 164400
rect 129002 163200 129058 164400
rect 129922 163200 129978 164400
rect 130750 163200 130806 164400
rect 131578 163200 131634 164400
rect 132406 163200 132462 164400
rect 133234 163200 133290 164400
rect 134062 163200 134118 164400
rect 134890 163200 134946 164400
rect 135810 163200 135866 164400
rect 136638 163200 136694 164400
rect 137466 163200 137522 164400
rect 138294 163200 138350 164400
rect 139122 163200 139178 164400
rect 139950 163200 140006 164400
rect 140778 163200 140834 164400
rect 141698 163200 141754 164400
rect 142526 163200 142582 164400
rect 143354 163200 143410 164400
rect 144182 163200 144238 164400
rect 145010 163200 145066 164400
rect 145838 163200 145894 164400
rect 146666 163200 146722 164400
rect 147586 163200 147642 164400
rect 148414 163200 148470 164400
rect 149242 163200 149298 164400
rect 150070 163200 150126 164400
rect 150898 163200 150954 164400
rect 151726 163200 151782 164400
rect 152554 163200 152610 164400
rect 153474 163200 153530 164400
rect 154302 163200 154358 164400
rect 155130 163200 155186 164400
rect 155958 163200 156014 164400
rect 156786 163200 156842 164400
rect 157614 163200 157670 164400
rect 158442 163200 158498 164400
rect 159362 163200 159418 164400
rect 160190 163200 160246 164400
rect 161018 163200 161074 164400
rect 161124 163254 161428 163282
rect 122748 158772 122800 158778
rect 122748 158714 122800 158720
rect 121736 153876 121788 153882
rect 121736 153818 121788 153824
rect 122656 153876 122708 153882
rect 122656 153818 122708 153824
rect 121748 150226 121776 153818
rect 122380 152448 122432 152454
rect 122380 152390 122432 152396
rect 122392 150226 122420 152390
rect 122760 151706 122788 158714
rect 123128 157894 123156 163200
rect 124048 159730 124076 163200
rect 124876 160682 124904 163200
rect 125704 161474 125732 163200
rect 125704 161446 125824 161474
rect 124864 160676 124916 160682
rect 124864 160618 124916 160624
rect 124036 159724 124088 159730
rect 124036 159666 124088 159672
rect 123944 159384 123996 159390
rect 123944 159326 123996 159332
rect 123116 157888 123168 157894
rect 123116 157830 123168 157836
rect 123024 155304 123076 155310
rect 123024 155246 123076 155252
rect 122748 151700 122800 151706
rect 122748 151642 122800 151648
rect 119816 150198 119890 150226
rect 120460 150198 120534 150226
rect 121104 150198 121178 150226
rect 121748 150198 121822 150226
rect 122392 150198 122466 150226
rect 117228 149932 117280 149938
rect 118988 149926 119324 149954
rect 119862 149940 119890 150198
rect 120506 149940 120534 150198
rect 121150 149940 121178 150198
rect 121794 149940 121822 150198
rect 122438 149940 122466 150198
rect 123036 150192 123064 155246
rect 123668 152516 123720 152522
rect 123668 152458 123720 152464
rect 123680 150192 123708 152458
rect 123956 152454 123984 159326
rect 125508 158976 125560 158982
rect 125508 158918 125560 158924
rect 124770 156632 124826 156641
rect 124770 156567 124826 156576
rect 124310 153776 124366 153785
rect 124310 153711 124366 153720
rect 123944 152448 123996 152454
rect 123944 152390 123996 152396
rect 124324 150192 124352 153711
rect 124784 151814 124812 156567
rect 125520 153785 125548 158918
rect 125692 156732 125744 156738
rect 125692 156674 125744 156680
rect 125600 155440 125652 155446
rect 125600 155382 125652 155388
rect 125506 153776 125562 153785
rect 125506 153711 125562 153720
rect 124784 151786 124996 151814
rect 124968 150226 124996 151786
rect 124968 150198 125042 150226
rect 123036 150164 123110 150192
rect 123680 150164 123754 150192
rect 124324 150164 124398 150192
rect 123082 149940 123110 150164
rect 123726 149940 123754 150164
rect 124370 149940 124398 150164
rect 125014 149940 125042 150198
rect 125612 150192 125640 155382
rect 125704 152522 125732 156674
rect 125796 155242 125824 161446
rect 126532 156738 126560 163200
rect 127360 159118 127388 163200
rect 127622 159352 127678 159361
rect 127622 159287 127678 159296
rect 127348 159112 127400 159118
rect 127348 159054 127400 159060
rect 127070 157992 127126 158001
rect 127070 157927 127126 157936
rect 126520 156732 126572 156738
rect 126520 156674 126572 156680
rect 125784 155236 125836 155242
rect 125784 155178 125836 155184
rect 126886 153912 126942 153921
rect 126886 153847 126942 153856
rect 125692 152516 125744 152522
rect 125692 152458 125744 152464
rect 126334 152416 126390 152425
rect 126334 152351 126390 152360
rect 126348 150226 126376 152351
rect 126302 150198 126376 150226
rect 125612 150164 125686 150192
rect 125658 149940 125686 150164
rect 126302 149940 126330 150198
rect 126900 150192 126928 153847
rect 127084 150210 127112 157927
rect 127532 152516 127584 152522
rect 127532 152458 127584 152464
rect 127072 150204 127124 150210
rect 126900 150164 126974 150192
rect 126946 149940 126974 150164
rect 127544 150192 127572 152458
rect 127636 151910 127664 159287
rect 128188 155038 128216 163200
rect 128360 159656 128412 159662
rect 128360 159598 128412 159604
rect 128176 155032 128228 155038
rect 128176 154974 128228 154980
rect 128372 153678 128400 159598
rect 129016 158778 129044 163200
rect 129832 159452 129884 159458
rect 129832 159394 129884 159400
rect 129004 158772 129056 158778
rect 129004 158714 129056 158720
rect 129740 156664 129792 156670
rect 129740 156606 129792 156612
rect 129464 154080 129516 154086
rect 129464 154022 129516 154028
rect 128360 153672 128412 153678
rect 128360 153614 128412 153620
rect 128820 152448 128872 152454
rect 128820 152390 128872 152396
rect 127624 151904 127676 151910
rect 127624 151846 127676 151852
rect 128222 150204 128274 150210
rect 127544 150164 127618 150192
rect 127072 150146 127124 150152
rect 127590 149940 127618 150164
rect 128832 150192 128860 152390
rect 129476 150192 129504 154022
rect 129752 151814 129780 156606
rect 129844 152454 129872 159394
rect 129936 156670 129964 163200
rect 130764 159662 130792 163200
rect 130752 159656 130804 159662
rect 130752 159598 130804 159604
rect 131592 158778 131620 163200
rect 132420 159390 132448 163200
rect 132408 159384 132460 159390
rect 132408 159326 132460 159332
rect 131120 158772 131172 158778
rect 131120 158714 131172 158720
rect 131580 158772 131632 158778
rect 131580 158714 131632 158720
rect 132408 158772 132460 158778
rect 132408 158714 132460 158720
rect 129924 156664 129976 156670
rect 129924 156606 129976 156612
rect 130292 155508 130344 155514
rect 130292 155450 130344 155456
rect 129832 152448 129884 152454
rect 129832 152390 129884 152396
rect 130304 151814 130332 155450
rect 131132 154086 131160 158714
rect 131120 154080 131172 154086
rect 131120 154022 131172 154028
rect 132040 153944 132092 153950
rect 132040 153886 132092 153892
rect 131394 152552 131450 152561
rect 131394 152487 131450 152496
rect 129752 151786 130148 151814
rect 130304 151786 130792 151814
rect 130120 150226 130148 151786
rect 130764 150226 130792 151786
rect 130120 150198 130194 150226
rect 130764 150198 130838 150226
rect 128832 150164 128906 150192
rect 129476 150164 129550 150192
rect 128222 150146 128274 150152
rect 128234 149940 128262 150146
rect 128878 149940 128906 150164
rect 129522 149940 129550 150164
rect 130166 149940 130194 150198
rect 130810 149940 130838 150198
rect 131408 150192 131436 152487
rect 132052 150192 132080 153886
rect 132420 151774 132448 158714
rect 132500 158092 132552 158098
rect 132500 158034 132552 158040
rect 132408 151768 132460 151774
rect 132408 151710 132460 151716
rect 132512 150210 132540 158034
rect 133248 158030 133276 163200
rect 133512 159792 133564 159798
rect 133512 159734 133564 159740
rect 133236 158024 133288 158030
rect 133236 157966 133288 157972
rect 132684 156800 132736 156806
rect 132684 156742 132736 156748
rect 132696 150226 132724 156742
rect 133524 156398 133552 159734
rect 133512 156392 133564 156398
rect 133512 156334 133564 156340
rect 134076 152522 134104 163200
rect 134904 154902 134932 163200
rect 135824 161474 135852 163200
rect 135824 161446 135944 161474
rect 135628 159996 135680 160002
rect 135628 159938 135680 159944
rect 135260 156868 135312 156874
rect 135260 156810 135312 156816
rect 134892 154896 134944 154902
rect 134892 154838 134944 154844
rect 134616 154012 134668 154018
rect 134616 153954 134668 153960
rect 134064 152516 134116 152522
rect 134064 152458 134116 152464
rect 133972 151904 134024 151910
rect 133972 151846 134024 151852
rect 133984 150226 134012 151846
rect 134628 150226 134656 153954
rect 135272 150226 135300 156810
rect 135640 156466 135668 159938
rect 135628 156460 135680 156466
rect 135628 156402 135680 156408
rect 135812 155576 135864 155582
rect 135812 155518 135864 155524
rect 135824 151814 135852 155518
rect 135916 153950 135944 161446
rect 136362 159488 136418 159497
rect 136362 159423 136418 159432
rect 136088 159384 136140 159390
rect 136088 159326 136140 159332
rect 136100 155310 136128 159326
rect 136088 155304 136140 155310
rect 136088 155246 136140 155252
rect 135904 153944 135956 153950
rect 135904 153886 135956 153892
rect 136376 151978 136404 159423
rect 136652 156806 136680 163200
rect 137480 159497 137508 163200
rect 137466 159488 137522 159497
rect 137466 159423 137522 159432
rect 137836 156936 137888 156942
rect 137836 156878 137888 156884
rect 136640 156800 136692 156806
rect 136640 156742 136692 156748
rect 136732 155644 136784 155650
rect 136732 155586 136784 155592
rect 136548 152584 136600 152590
rect 136548 152526 136600 152532
rect 136364 151972 136416 151978
rect 136364 151914 136416 151920
rect 135824 151786 135944 151814
rect 135916 150226 135944 151786
rect 136560 150226 136588 152526
rect 136744 151814 136772 155586
rect 136744 151786 137232 151814
rect 137204 150226 137232 151786
rect 137848 150226 137876 156878
rect 138308 155446 138336 163200
rect 139136 159458 139164 163200
rect 139124 159452 139176 159458
rect 139124 159394 139176 159400
rect 139492 158228 139544 158234
rect 139492 158170 139544 158176
rect 139398 156768 139454 156777
rect 139398 156703 139454 156712
rect 138296 155440 138348 155446
rect 138296 155382 138348 155388
rect 138480 154148 138532 154154
rect 138480 154090 138532 154096
rect 138492 150226 138520 154090
rect 139124 152448 139176 152454
rect 139124 152390 139176 152396
rect 139136 150226 139164 152390
rect 132500 150204 132552 150210
rect 131408 150164 131482 150192
rect 132052 150164 132126 150192
rect 131454 149940 131482 150164
rect 132098 149940 132126 150164
rect 132696 150198 132770 150226
rect 132500 150146 132552 150152
rect 132742 149940 132770 150198
rect 133374 150204 133426 150210
rect 133984 150198 134058 150226
rect 134628 150198 134702 150226
rect 135272 150198 135346 150226
rect 135916 150198 135990 150226
rect 136560 150198 136634 150226
rect 137204 150198 137278 150226
rect 137848 150198 137922 150226
rect 138492 150198 138566 150226
rect 139136 150198 139210 150226
rect 139412 150210 139440 156703
rect 139504 151910 139532 158170
rect 139964 158098 139992 163200
rect 140792 159390 140820 163200
rect 141712 160614 141740 163200
rect 141700 160608 141752 160614
rect 141700 160550 141752 160556
rect 140780 159384 140832 159390
rect 140780 159326 140832 159332
rect 139952 158092 140004 158098
rect 139952 158034 140004 158040
rect 142342 155408 142398 155417
rect 142342 155343 142398 155352
rect 139766 155272 139822 155281
rect 139766 155207 139822 155216
rect 139492 151904 139544 151910
rect 139492 151846 139544 151852
rect 139780 150226 139808 155207
rect 141698 152688 141754 152697
rect 141698 152623 141754 152632
rect 141054 151192 141110 151201
rect 141054 151127 141110 151136
rect 133374 150146 133426 150152
rect 133386 149940 133414 150146
rect 134030 149940 134058 150198
rect 134674 149940 134702 150198
rect 135318 149940 135346 150198
rect 135962 149940 135990 150198
rect 136606 149940 136634 150198
rect 137250 149940 137278 150198
rect 137894 149940 137922 150198
rect 138538 149940 138566 150198
rect 139182 149940 139210 150198
rect 139400 150204 139452 150210
rect 139780 150198 139854 150226
rect 139400 150146 139452 150152
rect 139826 149940 139854 150198
rect 140458 150204 140510 150210
rect 140458 150146 140510 150152
rect 140470 149940 140498 150146
rect 141068 150090 141096 151127
rect 141712 150226 141740 152623
rect 142356 150226 142384 155343
rect 142540 155281 142568 163200
rect 142526 155272 142582 155281
rect 142526 155207 142582 155216
rect 143368 154018 143396 163200
rect 144196 159254 144224 163200
rect 144184 159248 144236 159254
rect 144184 159190 144236 159196
rect 145024 158778 145052 163200
rect 145852 158846 145880 163200
rect 145930 159624 145986 159633
rect 145930 159559 145986 159568
rect 145840 158840 145892 158846
rect 145840 158782 145892 158788
rect 145012 158772 145064 158778
rect 145012 158714 145064 158720
rect 145104 158160 145156 158166
rect 143630 158128 143686 158137
rect 145104 158102 145156 158108
rect 143630 158063 143686 158072
rect 143356 154012 143408 154018
rect 143356 153954 143408 153960
rect 142988 151904 143040 151910
rect 142988 151846 143040 151852
rect 143000 150226 143028 151846
rect 143644 150226 143672 158063
rect 144828 154828 144880 154834
rect 144828 154770 144880 154776
rect 144840 152454 144868 154770
rect 144920 152652 144972 152658
rect 144920 152594 144972 152600
rect 144828 152448 144880 152454
rect 144828 152390 144880 152396
rect 144276 151972 144328 151978
rect 144276 151914 144328 151920
rect 144288 150226 144316 151914
rect 144932 150226 144960 152594
rect 141712 150198 141786 150226
rect 142356 150198 142430 150226
rect 143000 150198 143074 150226
rect 143644 150198 143718 150226
rect 144288 150198 144362 150226
rect 144932 150198 145006 150226
rect 145116 150210 145144 158102
rect 145564 154216 145616 154222
rect 145564 154158 145616 154164
rect 145576 150226 145604 154158
rect 145944 153921 145972 159559
rect 146024 159316 146076 159322
rect 146024 159258 146076 159264
rect 146036 157758 146064 159258
rect 146116 159180 146168 159186
rect 146116 159122 146168 159128
rect 146128 158001 146156 159122
rect 146208 158772 146260 158778
rect 146208 158714 146260 158720
rect 146114 157992 146170 158001
rect 146114 157927 146170 157936
rect 146116 157820 146168 157826
rect 146116 157762 146168 157768
rect 146024 157752 146076 157758
rect 146024 157694 146076 157700
rect 145930 153912 145986 153921
rect 145930 153847 145986 153856
rect 146128 152250 146156 157762
rect 146116 152244 146168 152250
rect 146116 152186 146168 152192
rect 146220 151026 146248 158714
rect 146680 155378 146708 163200
rect 146852 160744 146904 160750
rect 146852 160686 146904 160692
rect 146668 155372 146720 155378
rect 146668 155314 146720 155320
rect 146208 151020 146260 151026
rect 146208 150962 146260 150968
rect 146864 150226 146892 160686
rect 147600 152590 147628 163200
rect 148428 160750 148456 163200
rect 149152 160812 149204 160818
rect 149152 160754 149204 160760
rect 148416 160744 148468 160750
rect 148416 160686 148468 160692
rect 147772 159928 147824 159934
rect 147772 159870 147824 159876
rect 147680 159112 147732 159118
rect 147680 159054 147732 159060
rect 147692 157826 147720 159054
rect 147680 157820 147732 157826
rect 147680 157762 147732 157768
rect 147680 157004 147732 157010
rect 147680 156946 147732 156952
rect 147588 152584 147640 152590
rect 147588 152526 147640 152532
rect 147496 151088 147548 151094
rect 147496 151030 147548 151036
rect 141068 150062 141142 150090
rect 141114 149940 141142 150062
rect 141758 149940 141786 150198
rect 142402 149940 142430 150198
rect 143046 149940 143074 150198
rect 143690 149940 143718 150198
rect 144334 149940 144362 150198
rect 144978 149940 145006 150198
rect 145104 150204 145156 150210
rect 145576 150198 145650 150226
rect 145104 150146 145156 150152
rect 145622 149940 145650 150198
rect 146254 150204 146306 150210
rect 146864 150198 146938 150226
rect 146254 150146 146306 150152
rect 146266 149940 146294 150146
rect 146910 149940 146938 150198
rect 147508 150090 147536 151030
rect 147692 150210 147720 156946
rect 147784 154222 147812 159870
rect 147772 154216 147824 154222
rect 147772 154158 147824 154164
rect 148138 154048 148194 154057
rect 148138 153983 148194 153992
rect 148152 150226 148180 153983
rect 147680 150204 147732 150210
rect 148152 150198 148226 150226
rect 149164 150210 149192 160754
rect 149256 160546 149284 163200
rect 149428 162580 149480 162586
rect 149428 162522 149480 162528
rect 149244 160540 149296 160546
rect 149244 160482 149296 160488
rect 149440 150226 149468 162522
rect 150084 156874 150112 163200
rect 150912 159934 150940 163200
rect 150900 159928 150952 159934
rect 150900 159870 150952 159876
rect 150440 158840 150492 158846
rect 150440 158782 150492 158788
rect 150072 156868 150124 156874
rect 150072 156810 150124 156816
rect 150452 155582 150480 158782
rect 150530 158264 150586 158273
rect 150530 158199 150586 158208
rect 150440 155576 150492 155582
rect 150440 155518 150492 155524
rect 147680 150146 147732 150152
rect 147508 150062 147582 150090
rect 147554 149940 147582 150062
rect 148198 149940 148226 150198
rect 148830 150204 148882 150210
rect 148830 150146 148882 150152
rect 149152 150204 149204 150210
rect 149440 150198 149514 150226
rect 150544 150210 150572 158199
rect 150624 155712 150676 155718
rect 150624 155654 150676 155660
rect 150636 150226 150664 155654
rect 151740 151094 151768 163200
rect 151912 162648 151964 162654
rect 151912 162590 151964 162596
rect 151728 151088 151780 151094
rect 151728 151030 151780 151036
rect 149152 150146 149204 150152
rect 148842 149940 148870 150146
rect 149486 149940 149514 150198
rect 150026 150204 150078 150210
rect 150026 150146 150078 150152
rect 150532 150204 150584 150210
rect 150636 150198 150710 150226
rect 150532 150146 150584 150152
rect 150038 149940 150066 150146
rect 150682 149940 150710 150198
rect 151314 150204 151366 150210
rect 151924 150192 151952 162590
rect 152568 158778 152596 163200
rect 152556 158772 152608 158778
rect 152556 158714 152608 158720
rect 153108 158772 153160 158778
rect 153108 158714 153160 158720
rect 152554 151328 152610 151337
rect 152554 151263 152610 151272
rect 151924 150164 151998 150192
rect 151314 150146 151366 150152
rect 151326 149940 151354 150146
rect 151970 149940 151998 150164
rect 152568 150090 152596 151263
rect 153120 150958 153148 158714
rect 153384 158296 153436 158302
rect 153384 158238 153436 158244
rect 153200 154284 153252 154290
rect 153200 154226 153252 154232
rect 153108 150952 153160 150958
rect 153108 150894 153160 150900
rect 153212 150192 153240 154226
rect 153396 151814 153424 158238
rect 153488 158166 153516 163200
rect 153476 158160 153528 158166
rect 153476 158102 153528 158108
rect 154212 154964 154264 154970
rect 154212 154906 154264 154912
rect 154224 151814 154252 154906
rect 154316 154290 154344 163200
rect 155040 160880 155092 160886
rect 155040 160822 155092 160828
rect 154672 155780 154724 155786
rect 154672 155722 154724 155728
rect 154304 154284 154356 154290
rect 154304 154226 154356 154232
rect 153396 151786 153884 151814
rect 154224 151786 154528 151814
rect 153856 150226 153884 151786
rect 154500 150226 154528 151786
rect 153856 150198 153930 150226
rect 154500 150198 154574 150226
rect 154684 150210 154712 155722
rect 155052 151814 155080 160822
rect 155144 160818 155172 163200
rect 155132 160812 155184 160818
rect 155132 160754 155184 160760
rect 155972 159186 156000 163200
rect 155960 159180 156012 159186
rect 155960 159122 156012 159128
rect 156420 157072 156472 157078
rect 156420 157014 156472 157020
rect 155052 151786 155172 151814
rect 155144 150226 155172 151786
rect 153212 150164 153286 150192
rect 152568 150062 152642 150090
rect 152614 149940 152642 150062
rect 153258 149940 153286 150164
rect 153902 149940 153930 150198
rect 154546 149940 154574 150198
rect 154672 150204 154724 150210
rect 155144 150198 155218 150226
rect 154672 150146 154724 150152
rect 155190 149940 155218 150198
rect 155822 150204 155874 150210
rect 156432 150192 156460 157014
rect 156800 155514 156828 163200
rect 157628 159798 157656 163200
rect 158456 161474 158484 163200
rect 158456 161446 158668 161474
rect 157616 159792 157668 159798
rect 157616 159734 157668 159740
rect 158444 159588 158496 159594
rect 158444 159530 158496 159536
rect 157340 159452 157392 159458
rect 157340 159394 157392 159400
rect 156788 155508 156840 155514
rect 156788 155450 156840 155456
rect 157352 154970 157380 159394
rect 157340 154964 157392 154970
rect 157340 154906 157392 154912
rect 156604 154420 156656 154426
rect 156604 154362 156656 154368
rect 156616 154154 156644 154362
rect 158456 154358 158484 159530
rect 158352 154352 158404 154358
rect 158352 154294 158404 154300
rect 158444 154352 158496 154358
rect 158444 154294 158496 154300
rect 156604 154148 156656 154154
rect 156604 154090 156656 154096
rect 157062 152824 157118 152833
rect 157062 152759 157118 152768
rect 157076 150192 157104 152759
rect 157708 151156 157760 151162
rect 157708 151098 157760 151104
rect 156432 150164 156506 150192
rect 157076 150164 157150 150192
rect 155822 150146 155874 150152
rect 155834 149940 155862 150146
rect 156478 149940 156506 150164
rect 157122 149940 157150 150164
rect 157720 150090 157748 151098
rect 158364 150192 158392 154294
rect 158640 151162 158668 161446
rect 159376 159361 159404 163200
rect 159362 159352 159418 159361
rect 159362 159287 159418 159296
rect 158996 158364 159048 158370
rect 158996 158306 159048 158312
rect 158628 151156 158680 151162
rect 158628 151098 158680 151104
rect 159008 150192 159036 158306
rect 160204 156942 160232 163200
rect 161032 163146 161060 163200
rect 161124 163146 161152 163254
rect 161032 163118 161152 163146
rect 160376 160948 160428 160954
rect 160376 160890 160428 160896
rect 160284 159860 160336 159866
rect 160284 159802 160336 159808
rect 160192 156936 160244 156942
rect 160192 156878 160244 156884
rect 160100 155848 160152 155854
rect 160100 155790 160152 155796
rect 159640 153672 159692 153678
rect 159640 153614 159692 153620
rect 159652 150192 159680 153614
rect 160112 150210 160140 155790
rect 160296 155650 160324 159802
rect 160284 155644 160336 155650
rect 160284 155586 160336 155592
rect 160388 150226 160416 160890
rect 161400 152425 161428 163254
rect 161846 163200 161902 164400
rect 162674 163200 162730 164400
rect 163502 163200 163558 164400
rect 164330 163200 164386 164400
rect 165250 163200 165306 164400
rect 166078 163200 166134 164400
rect 166906 163200 166962 164400
rect 167734 163200 167790 164400
rect 168562 163200 168618 164400
rect 169390 163200 169446 164400
rect 170218 163200 170274 164400
rect 171138 163200 171194 164400
rect 171966 163200 172022 164400
rect 172072 163254 172468 163282
rect 161480 161628 161532 161634
rect 161480 161570 161532 161576
rect 161386 152416 161442 152425
rect 161386 152351 161442 152360
rect 160100 150204 160152 150210
rect 158364 150164 158438 150192
rect 159008 150164 159082 150192
rect 159652 150164 159726 150192
rect 157720 150062 157794 150090
rect 157766 149940 157794 150062
rect 158410 149940 158438 150164
rect 159054 149940 159082 150164
rect 159698 149940 159726 150164
rect 160100 150146 160152 150152
rect 160342 150198 160416 150226
rect 161492 150210 161520 161570
rect 161860 160886 161888 163200
rect 161848 160880 161900 160886
rect 161848 160822 161900 160828
rect 161572 157140 161624 157146
rect 161572 157082 161624 157088
rect 161584 150226 161612 157082
rect 162688 156641 162716 163200
rect 163044 158432 163096 158438
rect 163044 158374 163096 158380
rect 162674 156632 162730 156641
rect 162674 156567 162730 156576
rect 162860 151224 162912 151230
rect 162860 151166 162912 151172
rect 160974 150204 161026 150210
rect 160342 149940 160370 150198
rect 160974 150146 161026 150152
rect 161480 150204 161532 150210
rect 161584 150198 161658 150226
rect 161480 150146 161532 150152
rect 160986 149940 161014 150146
rect 161630 149940 161658 150198
rect 162262 150204 162314 150210
rect 162262 150146 162314 150152
rect 162274 149940 162302 150146
rect 162872 150090 162900 151166
rect 163056 150210 163084 158374
rect 163516 158234 163544 163200
rect 164344 160002 164372 163200
rect 164332 159996 164384 160002
rect 164332 159938 164384 159944
rect 165264 158778 165292 163200
rect 165620 161696 165672 161702
rect 165620 161638 165672 161644
rect 165436 161016 165488 161022
rect 165436 160958 165488 160964
rect 165252 158772 165304 158778
rect 165252 158714 165304 158720
rect 163504 158228 163556 158234
rect 163504 158170 163556 158176
rect 164424 156392 164476 156398
rect 164424 156334 164476 156340
rect 163504 154148 163556 154154
rect 163504 154090 163556 154096
rect 163516 150226 163544 154090
rect 164436 151814 164464 156334
rect 164436 151786 164832 151814
rect 164804 150226 164832 151786
rect 165448 150226 165476 160958
rect 165632 151814 165660 161638
rect 166092 160954 166120 163200
rect 166080 160948 166132 160954
rect 166080 160890 166132 160896
rect 166724 158568 166776 158574
rect 166724 158510 166776 158516
rect 165632 151786 166120 151814
rect 166092 150226 166120 151786
rect 166736 150226 166764 158510
rect 166920 150890 166948 163200
rect 167644 158772 167696 158778
rect 167644 158714 167696 158720
rect 167368 152380 167420 152386
rect 167368 152322 167420 152328
rect 166908 150884 166960 150890
rect 166908 150826 166960 150832
rect 167380 150226 167408 152322
rect 167656 151298 167684 158714
rect 167748 152658 167776 163200
rect 168472 161832 168524 161838
rect 168472 161774 168524 161780
rect 168380 158500 168432 158506
rect 168380 158442 168432 158448
rect 167736 152652 167788 152658
rect 167736 152594 167788 152600
rect 167644 151292 167696 151298
rect 167644 151234 167696 151240
rect 168012 151224 168064 151230
rect 168012 151166 168064 151172
rect 168104 151224 168156 151230
rect 168104 151166 168156 151172
rect 163044 150204 163096 150210
rect 163516 150198 163590 150226
rect 163044 150146 163096 150152
rect 162872 150062 162946 150090
rect 162918 149940 162946 150062
rect 163562 149940 163590 150198
rect 164194 150204 164246 150210
rect 164804 150198 164878 150226
rect 165448 150198 165522 150226
rect 166092 150198 166166 150226
rect 166736 150198 166810 150226
rect 167380 150198 167454 150226
rect 164194 150146 164246 150152
rect 164206 149940 164234 150146
rect 164850 149940 164878 150198
rect 165494 149940 165522 150198
rect 166138 149940 166166 150198
rect 166782 149940 166810 150198
rect 167426 149940 167454 150198
rect 168024 150090 168052 151166
rect 168116 150890 168144 151166
rect 168104 150884 168156 150890
rect 168104 150826 168156 150832
rect 168392 150210 168420 158442
rect 168484 151814 168512 161774
rect 168576 153678 168604 163200
rect 169404 157010 169432 163200
rect 169760 161084 169812 161090
rect 169760 161026 169812 161032
rect 169392 157004 169444 157010
rect 169392 156946 169444 156952
rect 168564 153672 168616 153678
rect 168564 153614 168616 153620
rect 168484 151786 168696 151814
rect 168668 150226 168696 151786
rect 168380 150204 168432 150210
rect 168668 150198 168742 150226
rect 169772 150210 169800 161026
rect 170232 159594 170260 163200
rect 171152 159866 171180 163200
rect 171980 163146 172008 163200
rect 172072 163146 172100 163254
rect 171980 163118 172100 163146
rect 171324 161764 171376 161770
rect 171324 161706 171376 161712
rect 171140 159860 171192 159866
rect 171140 159802 171192 159808
rect 170220 159588 170272 159594
rect 170220 159530 170272 159536
rect 171140 157276 171192 157282
rect 171140 157218 171192 157224
rect 169944 156460 169996 156466
rect 169944 156402 169996 156408
rect 169956 150226 169984 156402
rect 168380 150146 168432 150152
rect 168024 150062 168098 150090
rect 168070 149940 168098 150062
rect 168714 149940 168742 150198
rect 169346 150204 169398 150210
rect 169346 150146 169398 150152
rect 169760 150204 169812 150210
rect 169956 150198 170030 150226
rect 171152 150210 171180 157218
rect 171336 150226 171364 161706
rect 172440 154154 172468 163254
rect 172794 163200 172850 164400
rect 173622 163200 173678 164400
rect 174450 163200 174506 164400
rect 175278 163200 175334 164400
rect 176106 163200 176162 164400
rect 177026 163200 177082 164400
rect 177854 163200 177910 164400
rect 178682 163200 178738 164400
rect 179510 163200 179566 164400
rect 180338 163200 180394 164400
rect 180444 163254 180748 163282
rect 172704 162036 172756 162042
rect 172704 161978 172756 161984
rect 172428 154148 172480 154154
rect 172428 154090 172480 154096
rect 172518 153912 172574 153921
rect 172518 153847 172574 153856
rect 169760 150146 169812 150152
rect 169358 149940 169386 150146
rect 170002 149940 170030 150198
rect 170634 150204 170686 150210
rect 170634 150146 170686 150152
rect 171140 150204 171192 150210
rect 171140 150146 171192 150152
rect 171290 150198 171364 150226
rect 172532 150226 172560 153847
rect 171922 150204 171974 150210
rect 170646 149940 170674 150146
rect 171290 149940 171318 150198
rect 172532 150198 172606 150226
rect 172716 150210 172744 161978
rect 172808 157146 172836 163200
rect 173636 158302 173664 163200
rect 173992 159384 174044 159390
rect 173992 159326 174044 159332
rect 173624 158296 173676 158302
rect 173624 158238 173676 158244
rect 172796 157140 172848 157146
rect 172796 157082 172848 157088
rect 174004 152318 174032 159326
rect 174464 159118 174492 163200
rect 175292 161022 175320 163200
rect 175556 161900 175608 161906
rect 175556 161842 175608 161848
rect 175280 161016 175332 161022
rect 175280 160958 175332 160964
rect 175462 160712 175518 160721
rect 175462 160647 175518 160656
rect 174452 159112 174504 159118
rect 174452 159054 174504 159060
rect 174452 155916 174504 155922
rect 174452 155858 174504 155864
rect 173992 152312 174044 152318
rect 173992 152254 174044 152260
rect 173162 151464 173218 151473
rect 173162 151399 173218 151408
rect 171922 150146 171974 150152
rect 171934 149940 171962 150146
rect 172578 149940 172606 150198
rect 172704 150204 172756 150210
rect 172704 150146 172756 150152
rect 173176 150090 173204 151399
rect 174464 150226 174492 155858
rect 175096 152720 175148 152726
rect 175096 152662 175148 152668
rect 175108 150226 175136 152662
rect 173854 150204 173906 150210
rect 174464 150198 174538 150226
rect 175108 150198 175182 150226
rect 173854 150146 173906 150152
rect 173176 150062 173250 150090
rect 173222 149940 173250 150062
rect 173866 149940 173894 150146
rect 174510 149940 174538 150198
rect 175154 149940 175182 150198
rect 175476 150192 175504 160647
rect 175568 151814 175596 161842
rect 176120 157078 176148 163200
rect 176660 159588 176712 159594
rect 176660 159530 176712 159536
rect 176108 157072 176160 157078
rect 176108 157014 176160 157020
rect 176672 156466 176700 159530
rect 177040 158370 177068 163200
rect 177868 159458 177896 163200
rect 178224 161968 178276 161974
rect 178224 161910 178276 161916
rect 177856 159452 177908 159458
rect 177856 159394 177908 159400
rect 177028 158364 177080 158370
rect 177028 158306 177080 158312
rect 177028 157344 177080 157350
rect 177028 157286 177080 157292
rect 176660 156460 176712 156466
rect 176660 156402 176712 156408
rect 175568 151786 176424 151814
rect 176396 150226 176424 151786
rect 177040 150226 177068 157286
rect 177672 154216 177724 154222
rect 177672 154158 177724 154164
rect 177684 150226 177712 154158
rect 178236 151814 178264 161910
rect 178696 153921 178724 163200
rect 179420 159520 179472 159526
rect 179420 159462 179472 159468
rect 178682 153912 178738 153921
rect 178682 153847 178738 153856
rect 179432 152726 179460 159462
rect 179524 157282 179552 163200
rect 180352 163146 180380 163200
rect 180444 163146 180472 163254
rect 180352 163118 180472 163146
rect 179512 157276 179564 157282
rect 179512 157218 179564 157224
rect 180248 154352 180300 154358
rect 180248 154294 180300 154300
rect 179420 152720 179472 152726
rect 179420 152662 179472 152668
rect 179604 152244 179656 152250
rect 179604 152186 179656 152192
rect 178236 151786 179000 151814
rect 178316 151360 178368 151366
rect 178316 151302 178368 151308
rect 176396 150198 176470 150226
rect 177040 150198 177114 150226
rect 177684 150198 177758 150226
rect 175476 150164 175826 150192
rect 175798 149940 175826 150164
rect 176442 149940 176470 150198
rect 177086 149940 177114 150198
rect 177730 149940 177758 150198
rect 178328 150090 178356 151302
rect 178972 150226 179000 151786
rect 179616 150226 179644 152186
rect 180260 150226 180288 154294
rect 180720 151366 180748 163254
rect 181166 163200 181222 164400
rect 181994 163200 182050 164400
rect 182914 163200 182970 164400
rect 183742 163200 183798 164400
rect 184570 163200 184626 164400
rect 185398 163200 185454 164400
rect 186226 163200 186282 164400
rect 187054 163200 187110 164400
rect 187882 163200 187938 164400
rect 188802 163200 188858 164400
rect 189630 163200 189686 164400
rect 190458 163200 190514 164400
rect 191286 163200 191342 164400
rect 192114 163200 192170 164400
rect 192942 163200 192998 164400
rect 193770 163200 193826 164400
rect 194690 163200 194746 164400
rect 195518 163200 195574 164400
rect 195624 163254 195928 163282
rect 181076 162104 181128 162110
rect 181076 162046 181128 162052
rect 180892 161152 180944 161158
rect 180892 161094 180944 161100
rect 180708 151360 180760 151366
rect 180708 151302 180760 151308
rect 180904 150226 180932 161094
rect 180982 156904 181038 156913
rect 180982 156839 181038 156848
rect 178972 150198 179046 150226
rect 179616 150198 179690 150226
rect 180260 150198 180334 150226
rect 178328 150062 178402 150090
rect 178374 149940 178402 150062
rect 179018 149940 179046 150198
rect 179662 149940 179690 150198
rect 180306 149940 180334 150198
rect 180858 150198 180932 150226
rect 180996 150210 181024 156839
rect 181088 151814 181116 162046
rect 181180 159322 181208 163200
rect 181168 159316 181220 159322
rect 181168 159258 181220 159264
rect 182008 154222 182036 163200
rect 182928 156777 182956 163200
rect 183756 161090 183784 163200
rect 183744 161084 183796 161090
rect 183744 161026 183796 161032
rect 183284 160064 183336 160070
rect 183284 160006 183336 160012
rect 182914 156768 182970 156777
rect 182914 156703 182970 156712
rect 183296 154834 183324 160006
rect 184584 159526 184612 163200
rect 184572 159520 184624 159526
rect 184572 159462 184624 159468
rect 183560 158636 183612 158642
rect 183560 158578 183612 158584
rect 183284 154828 183336 154834
rect 183284 154770 183336 154776
rect 183284 154284 183336 154290
rect 183284 154226 183336 154232
rect 181996 154216 182048 154222
rect 181996 154158 182048 154164
rect 182732 152788 182784 152794
rect 182732 152730 182784 152736
rect 181088 151786 181484 151814
rect 181456 150226 181484 151786
rect 180984 150204 181036 150210
rect 180858 149940 180886 150198
rect 181456 150198 181530 150226
rect 180984 150146 181036 150152
rect 181502 149940 181530 150198
rect 182134 150204 182186 150210
rect 182744 150192 182772 152730
rect 183296 152386 183324 154226
rect 183284 152380 183336 152386
rect 183284 152322 183336 152328
rect 183374 151600 183430 151609
rect 183374 151535 183430 151544
rect 182744 150164 182818 150192
rect 182134 150146 182186 150152
rect 182146 149940 182174 150146
rect 182790 149940 182818 150164
rect 183388 150090 183416 151535
rect 183572 150210 183600 158578
rect 185032 155644 185084 155650
rect 185032 155586 185084 155592
rect 184018 155544 184074 155553
rect 184018 155479 184074 155488
rect 183560 150204 183612 150210
rect 184032 150192 184060 155479
rect 185044 151814 185072 155586
rect 185412 154358 185440 163200
rect 185950 160848 186006 160857
rect 185950 160783 186006 160792
rect 185400 154352 185452 154358
rect 185400 154294 185452 154300
rect 185044 151786 185348 151814
rect 185320 150226 185348 151786
rect 184710 150204 184762 150210
rect 184032 150164 184106 150192
rect 183560 150146 183612 150152
rect 183388 150062 183462 150090
rect 183434 149940 183462 150062
rect 184078 149940 184106 150164
rect 185320 150198 185394 150226
rect 184710 150146 184762 150152
rect 184722 149940 184750 150146
rect 185366 149940 185394 150198
rect 185964 150192 185992 160783
rect 186240 155650 186268 163200
rect 186320 162172 186372 162178
rect 186320 162114 186372 162120
rect 186228 155644 186280 155650
rect 186228 155586 186280 155592
rect 186332 151814 186360 162114
rect 187068 158438 187096 163200
rect 187896 160070 187924 163200
rect 187884 160064 187936 160070
rect 187884 160006 187936 160012
rect 187700 159724 187752 159730
rect 187700 159666 187752 159672
rect 187056 158432 187108 158438
rect 187056 158374 187108 158380
rect 187240 155168 187292 155174
rect 187240 155110 187292 155116
rect 186332 151786 186636 151814
rect 186608 150226 186636 151786
rect 186608 150198 186682 150226
rect 185964 150164 186038 150192
rect 186010 149940 186038 150164
rect 186654 149940 186682 150198
rect 187252 150192 187280 155110
rect 187712 152794 187740 159666
rect 188816 154290 188844 163200
rect 189172 162240 189224 162246
rect 189172 162182 189224 162188
rect 188804 154284 188856 154290
rect 188804 154226 188856 154232
rect 187884 152856 187936 152862
rect 187884 152798 187936 152804
rect 187700 152788 187752 152794
rect 187700 152730 187752 152736
rect 187896 150192 187924 152798
rect 188528 151428 188580 151434
rect 188528 151370 188580 151376
rect 187252 150164 187326 150192
rect 187896 150164 187970 150192
rect 187298 149940 187326 150164
rect 187942 149940 187970 150164
rect 188540 150090 188568 151370
rect 189184 150192 189212 162182
rect 189644 155417 189672 163200
rect 190472 158506 190500 163200
rect 190736 162376 190788 162382
rect 190736 162318 190788 162324
rect 190460 158500 190512 158506
rect 190460 158442 190512 158448
rect 190460 157752 190512 157758
rect 190460 157694 190512 157700
rect 189630 155408 189686 155417
rect 189630 155343 189686 155352
rect 189816 154488 189868 154494
rect 189816 154430 189868 154436
rect 189828 150192 189856 154430
rect 190472 150226 190500 157694
rect 190472 150198 190546 150226
rect 190748 150210 190776 162318
rect 191104 161220 191156 161226
rect 191104 161162 191156 161168
rect 191116 150226 191144 161162
rect 191300 159390 191328 163200
rect 191288 159384 191340 159390
rect 191288 159326 191340 159332
rect 192128 154426 192156 163200
rect 192576 159248 192628 159254
rect 192576 159190 192628 159196
rect 192392 156596 192444 156602
rect 192392 156538 192444 156544
rect 192116 154420 192168 154426
rect 192116 154362 192168 154368
rect 192404 150226 192432 156538
rect 192588 152862 192616 159190
rect 192956 155718 192984 163200
rect 193404 162308 193456 162314
rect 193404 162250 193456 162256
rect 192944 155712 192996 155718
rect 192944 155654 192996 155660
rect 193036 152924 193088 152930
rect 193036 152866 193088 152872
rect 192576 152856 192628 152862
rect 192576 152798 192628 152804
rect 193048 150226 193076 152866
rect 193416 151814 193444 162250
rect 193784 157350 193812 163200
rect 194704 159730 194732 163200
rect 195532 163146 195560 163200
rect 195624 163146 195652 163254
rect 195532 163118 195652 163146
rect 194692 159724 194744 159730
rect 194692 159666 194744 159672
rect 195244 159656 195296 159662
rect 195244 159598 195296 159604
rect 194968 158704 195020 158710
rect 194968 158646 195020 158652
rect 193772 157344 193824 157350
rect 193772 157286 193824 157292
rect 193416 151786 194364 151814
rect 193680 151496 193732 151502
rect 193680 151438 193732 151444
rect 189184 150164 189258 150192
rect 189828 150164 189902 150192
rect 188540 150062 188614 150090
rect 188586 149940 188614 150062
rect 189230 149940 189258 150164
rect 189874 149940 189902 150164
rect 190518 149940 190546 150198
rect 190736 150204 190788 150210
rect 191116 150198 191190 150226
rect 190736 150146 190788 150152
rect 191162 149940 191190 150198
rect 191794 150204 191846 150210
rect 192404 150198 192478 150226
rect 193048 150198 193122 150226
rect 191794 150146 191846 150152
rect 191806 149940 191834 150146
rect 192450 149940 192478 150198
rect 193094 149940 193122 150198
rect 193692 150090 193720 151438
rect 194336 150226 194364 151786
rect 194980 150226 195008 158646
rect 195256 152561 195284 159598
rect 195612 152720 195664 152726
rect 195612 152662 195664 152668
rect 195242 152552 195298 152561
rect 195242 152487 195298 152496
rect 195624 150226 195652 152662
rect 195900 151434 195928 163254
rect 196346 163200 196402 164400
rect 197174 163200 197230 164400
rect 198002 163200 198058 164400
rect 198830 163200 198886 164400
rect 199658 163200 199714 164400
rect 200578 163200 200634 164400
rect 201406 163200 201462 164400
rect 202234 163200 202290 164400
rect 203062 163200 203118 164400
rect 203890 163200 203946 164400
rect 204718 163200 204774 164400
rect 205546 163200 205602 164400
rect 206466 163200 206522 164400
rect 207294 163200 207350 164400
rect 208122 163200 208178 164400
rect 208950 163200 209006 164400
rect 209778 163200 209834 164400
rect 210606 163200 210662 164400
rect 211434 163200 211490 164400
rect 212354 163200 212410 164400
rect 213182 163200 213238 164400
rect 214010 163200 214066 164400
rect 214838 163200 214894 164400
rect 215666 163200 215722 164400
rect 216494 163200 216550 164400
rect 217322 163200 217378 164400
rect 218242 163200 218298 164400
rect 219070 163200 219126 164400
rect 219898 163200 219954 164400
rect 220726 163200 220782 164400
rect 221554 163200 221610 164400
rect 222382 163200 222438 164400
rect 223210 163200 223266 164400
rect 224130 163200 224186 164400
rect 224958 163200 225014 164400
rect 225786 163200 225842 164400
rect 226614 163200 226670 164400
rect 227442 163200 227498 164400
rect 228270 163200 228326 164400
rect 229098 163200 229154 164400
rect 230018 163200 230074 164400
rect 230846 163200 230902 164400
rect 231674 163200 231730 164400
rect 232502 163200 232558 164400
rect 233330 163200 233386 164400
rect 234158 163200 234214 164400
rect 234986 163200 235042 164400
rect 235906 163200 235962 164400
rect 236734 163200 236790 164400
rect 237562 163200 237618 164400
rect 238390 163200 238446 164400
rect 239218 163200 239274 164400
rect 240046 163200 240102 164400
rect 240874 163200 240930 164400
rect 241794 163200 241850 164400
rect 242622 163200 242678 164400
rect 243450 163200 243506 164400
rect 244278 163200 244334 164400
rect 245106 163200 245162 164400
rect 245934 163200 245990 164400
rect 246762 163200 246818 164400
rect 247682 163200 247738 164400
rect 248510 163200 248566 164400
rect 249338 163200 249394 164400
rect 250166 163200 250222 164400
rect 250994 163200 251050 164400
rect 251822 163200 251878 164400
rect 252650 163200 252706 164400
rect 253570 163200 253626 164400
rect 254398 163200 254454 164400
rect 255226 163200 255282 164400
rect 256054 163200 256110 164400
rect 256882 163200 256938 164400
rect 257710 163200 257766 164400
rect 258538 163200 258594 164400
rect 259458 163200 259514 164400
rect 260286 163200 260342 164400
rect 261114 163200 261170 164400
rect 261942 163200 261998 164400
rect 262770 163200 262826 164400
rect 263598 163200 263654 164400
rect 264426 163200 264482 164400
rect 265346 163200 265402 164400
rect 266174 163200 266230 164400
rect 267002 163200 267058 164400
rect 267830 163200 267886 164400
rect 268658 163200 268714 164400
rect 269486 163200 269542 164400
rect 270314 163200 270370 164400
rect 271234 163200 271290 164400
rect 272062 163200 272118 164400
rect 272890 163200 272946 164400
rect 273718 163200 273774 164400
rect 274546 163200 274602 164400
rect 275374 163200 275430 164400
rect 276202 163200 276258 164400
rect 277122 163200 277178 164400
rect 277950 163200 278006 164400
rect 278778 163200 278834 164400
rect 279606 163200 279662 164400
rect 280434 163200 280490 164400
rect 281262 163200 281318 164400
rect 282090 163200 282146 164400
rect 283010 163200 283066 164400
rect 283838 163200 283894 164400
rect 284666 163200 284722 164400
rect 285494 163200 285550 164400
rect 286322 163200 286378 164400
rect 287150 163200 287206 164400
rect 287978 163200 288034 164400
rect 288898 163200 288954 164400
rect 289726 163200 289782 164400
rect 290554 163200 290610 164400
rect 291382 163200 291438 164400
rect 292210 163200 292266 164400
rect 293038 163200 293094 164400
rect 293866 163200 293922 164400
rect 294786 163200 294842 164400
rect 295614 163200 295670 164400
rect 295720 163254 295932 163282
rect 196256 161288 196308 161294
rect 196256 161230 196308 161236
rect 195888 151428 195940 151434
rect 195888 151370 195940 151376
rect 196268 150226 196296 161230
rect 196360 158846 196388 163200
rect 196900 162512 196952 162518
rect 196900 162454 196952 162460
rect 196348 158840 196400 158846
rect 196348 158782 196400 158788
rect 196912 150226 196940 162454
rect 197188 158574 197216 163200
rect 198016 159594 198044 163200
rect 198844 161158 198872 163200
rect 198832 161152 198884 161158
rect 198832 161094 198884 161100
rect 198004 159588 198056 159594
rect 198004 159530 198056 159536
rect 197636 159180 197688 159186
rect 197636 159122 197688 159128
rect 197176 158568 197228 158574
rect 197176 158510 197228 158516
rect 197452 155032 197504 155038
rect 197452 154974 197504 154980
rect 197360 154896 197412 154902
rect 197360 154838 197412 154844
rect 197372 152250 197400 154838
rect 197360 152244 197412 152250
rect 197360 152186 197412 152192
rect 197464 152182 197492 154974
rect 197544 154556 197596 154562
rect 197544 154498 197596 154504
rect 197452 152176 197504 152182
rect 197452 152118 197504 152124
rect 197556 150226 197584 154498
rect 197648 153610 197676 159122
rect 198740 158840 198792 158846
rect 198740 158782 198792 158788
rect 198752 154494 198780 158782
rect 199672 155786 199700 163200
rect 200304 161356 200356 161362
rect 200304 161298 200356 161304
rect 200120 157956 200172 157962
rect 200120 157898 200172 157904
rect 199660 155780 199712 155786
rect 199660 155722 199712 155728
rect 198740 154488 198792 154494
rect 198740 154430 198792 154436
rect 199476 153808 199528 153814
rect 199476 153750 199528 153756
rect 197636 153604 197688 153610
rect 197636 153546 197688 153552
rect 198188 153196 198240 153202
rect 198188 153138 198240 153144
rect 198200 150226 198228 153138
rect 198832 151564 198884 151570
rect 198832 151506 198884 151512
rect 194336 150198 194410 150226
rect 194980 150198 195054 150226
rect 195624 150198 195698 150226
rect 196268 150198 196342 150226
rect 196912 150198 196986 150226
rect 197556 150198 197630 150226
rect 198200 150198 198274 150226
rect 193692 150062 193766 150090
rect 193738 149940 193766 150062
rect 194382 149940 194410 150198
rect 195026 149940 195054 150198
rect 195670 149940 195698 150198
rect 196314 149940 196342 150198
rect 196958 149940 196986 150198
rect 197602 149940 197630 150198
rect 198246 149940 198274 150198
rect 198844 150090 198872 151506
rect 199488 150226 199516 153750
rect 200132 150226 200160 157898
rect 199488 150198 199562 150226
rect 200132 150198 200206 150226
rect 200316 150210 200344 161298
rect 200592 158642 200620 163200
rect 201314 159488 201370 159497
rect 201314 159423 201370 159432
rect 200580 158636 200632 158642
rect 200580 158578 200632 158584
rect 201328 157758 201356 159423
rect 201420 159186 201448 163200
rect 202052 162444 202104 162450
rect 202052 162386 202104 162392
rect 201408 159180 201460 159186
rect 201408 159122 201460 159128
rect 201316 157752 201368 157758
rect 201316 157694 201368 157700
rect 201592 155100 201644 155106
rect 201592 155042 201644 155048
rect 200764 152992 200816 152998
rect 200764 152934 200816 152940
rect 200776 150226 200804 152934
rect 198844 150062 198918 150090
rect 198890 149940 198918 150062
rect 199534 149940 199562 150198
rect 200178 149940 200206 150198
rect 200304 150204 200356 150210
rect 200776 150198 200850 150226
rect 201604 150210 201632 155042
rect 202064 150226 202092 162386
rect 202248 158778 202276 163200
rect 202972 159112 203024 159118
rect 202972 159054 203024 159060
rect 202236 158772 202288 158778
rect 202236 158714 202288 158720
rect 202788 158772 202840 158778
rect 202788 158714 202840 158720
rect 202800 151502 202828 158714
rect 202984 153202 203012 159054
rect 203076 158778 203104 163200
rect 203064 158772 203116 158778
rect 203064 158714 203116 158720
rect 203338 157992 203394 158001
rect 203338 157927 203394 157936
rect 202972 153196 203024 153202
rect 202972 153138 203024 153144
rect 202788 151496 202840 151502
rect 202788 151438 202840 151444
rect 203352 150226 203380 157927
rect 203904 155922 203932 163200
rect 204260 161492 204312 161498
rect 204260 161434 204312 161440
rect 203892 155916 203944 155922
rect 203892 155858 203944 155864
rect 204272 151814 204300 161434
rect 204732 159497 204760 163200
rect 205560 161226 205588 163200
rect 206192 161424 206244 161430
rect 206192 161366 206244 161372
rect 205548 161220 205600 161226
rect 205548 161162 205600 161168
rect 204718 159488 204774 159497
rect 204718 159423 204774 159432
rect 205640 157888 205692 157894
rect 205640 157830 205692 157836
rect 205272 157208 205324 157214
rect 205272 157150 205324 157156
rect 204272 151786 204668 151814
rect 203984 151632 204036 151638
rect 203984 151574 204036 151580
rect 200304 150146 200356 150152
rect 200822 149940 200850 150198
rect 201454 150204 201506 150210
rect 201454 150146 201506 150152
rect 201592 150204 201644 150210
rect 202064 150198 202138 150226
rect 201592 150146 201644 150152
rect 201466 149940 201494 150146
rect 202110 149940 202138 150198
rect 202742 150204 202794 150210
rect 203352 150198 203426 150226
rect 202742 150146 202794 150152
rect 202754 149940 202782 150146
rect 203398 149940 203426 150198
rect 203996 150090 204024 151574
rect 204640 150226 204668 151786
rect 205284 150226 205312 157150
rect 205652 152998 205680 157830
rect 205916 153060 205968 153066
rect 205916 153002 205968 153008
rect 205640 152992 205692 152998
rect 205640 152934 205692 152940
rect 205928 150226 205956 153002
rect 206204 151814 206232 161366
rect 206480 155854 206508 163200
rect 207204 161560 207256 161566
rect 207204 161502 207256 161508
rect 207020 159928 207072 159934
rect 207020 159870 207072 159876
rect 207032 157962 207060 159870
rect 207020 157956 207072 157962
rect 207020 157898 207072 157904
rect 207020 156528 207072 156534
rect 207020 156470 207072 156476
rect 206468 155848 206520 155854
rect 206468 155790 206520 155796
rect 206204 151786 206600 151814
rect 206572 150226 206600 151786
rect 204640 150198 204714 150226
rect 205284 150198 205358 150226
rect 205928 150198 206002 150226
rect 206572 150198 206646 150226
rect 207032 150210 207060 156470
rect 207216 150226 207244 161502
rect 207308 158001 207336 163200
rect 208136 159254 208164 163200
rect 208964 159934 208992 163200
rect 208952 159928 209004 159934
rect 208952 159870 209004 159876
rect 208124 159248 208176 159254
rect 208124 159190 208176 159196
rect 208492 158772 208544 158778
rect 208492 158714 208544 158720
rect 207294 157992 207350 158001
rect 207294 157927 207350 157936
rect 208504 153814 208532 158714
rect 209792 157214 209820 163200
rect 210148 160064 210200 160070
rect 210148 160006 210200 160012
rect 209780 157208 209832 157214
rect 209780 157150 209832 157156
rect 209964 154828 210016 154834
rect 209964 154770 210016 154776
rect 208492 153808 208544 153814
rect 208492 153750 208544 153756
rect 209778 153776 209834 153785
rect 208400 153740 208452 153746
rect 209778 153711 209834 153720
rect 208400 153682 208452 153688
rect 208412 151842 208440 153682
rect 208492 153128 208544 153134
rect 208492 153070 208544 153076
rect 208400 151836 208452 151842
rect 208400 151778 208452 151784
rect 208504 150226 208532 153070
rect 209136 152448 209188 152454
rect 209136 152390 209188 152396
rect 209148 150226 209176 152390
rect 209792 150226 209820 153711
rect 203996 150062 204070 150090
rect 204042 149940 204070 150062
rect 204686 149940 204714 150198
rect 205330 149940 205358 150198
rect 205974 149940 206002 150198
rect 206618 149940 206646 150198
rect 207020 150204 207072 150210
rect 207216 150198 207290 150226
rect 207020 150146 207072 150152
rect 207262 149940 207290 150198
rect 207894 150204 207946 150210
rect 208504 150198 208578 150226
rect 209148 150198 209222 150226
rect 209792 150198 209866 150226
rect 209976 150210 210004 154770
rect 210160 152930 210188 160006
rect 210620 159050 210648 163200
rect 211448 159662 211476 163200
rect 212368 161474 212396 163200
rect 212368 161446 212488 161474
rect 211436 159656 211488 159662
rect 211436 159598 211488 159604
rect 211896 159180 211948 159186
rect 211896 159122 211948 159128
rect 210608 159044 210660 159050
rect 210608 158986 210660 158992
rect 210148 152924 210200 152930
rect 210148 152866 210200 152872
rect 211908 152726 211936 159122
rect 212264 153876 212316 153882
rect 212264 153818 212316 153824
rect 211896 152720 211948 152726
rect 211896 152662 211948 152668
rect 210424 151836 210476 151842
rect 210424 151778 210476 151784
rect 210436 150226 210464 151778
rect 211620 151700 211672 151706
rect 211620 151642 211672 151648
rect 207894 150146 207946 150152
rect 207906 149940 207934 150146
rect 208550 149940 208578 150198
rect 209194 149940 209222 150198
rect 209838 149940 209866 150198
rect 209964 150204 210016 150210
rect 210436 150198 210510 150226
rect 209964 150146 210016 150152
rect 210482 149940 210510 150198
rect 211114 150204 211166 150210
rect 211114 150146 211166 150152
rect 211126 149940 211154 150146
rect 211632 150090 211660 151642
rect 212276 150226 212304 153818
rect 212460 151570 212488 161446
rect 213196 153882 213224 163200
rect 213920 160676 213972 160682
rect 213920 160618 213972 160624
rect 213644 159724 213696 159730
rect 213644 159666 213696 159672
rect 213184 153876 213236 153882
rect 213184 153818 213236 153824
rect 213656 152998 213684 159666
rect 212908 152992 212960 152998
rect 212908 152934 212960 152940
rect 213644 152992 213696 152998
rect 213644 152934 213696 152940
rect 212448 151564 212500 151570
rect 212448 151506 212500 151512
rect 212920 150226 212948 152934
rect 213552 152788 213604 152794
rect 213552 152730 213604 152736
rect 213564 150226 213592 152730
rect 213932 151814 213960 160618
rect 214024 159118 214052 163200
rect 214852 159730 214880 163200
rect 214840 159724 214892 159730
rect 214840 159666 214892 159672
rect 214012 159112 214064 159118
rect 214012 159054 214064 159060
rect 215024 159044 215076 159050
rect 215024 158986 215076 158992
rect 215036 156602 215064 158986
rect 215392 157820 215444 157826
rect 215392 157762 215444 157768
rect 215024 156596 215076 156602
rect 215024 156538 215076 156544
rect 214840 155236 214892 155242
rect 214840 155178 214892 155184
rect 213932 151786 214236 151814
rect 214208 150226 214236 151786
rect 214852 150226 214880 155178
rect 215300 153672 215352 153678
rect 215300 153614 215352 153620
rect 215312 153134 215340 153614
rect 215300 153128 215352 153134
rect 215300 153070 215352 153076
rect 212276 150198 212350 150226
rect 212920 150198 212994 150226
rect 213564 150198 213638 150226
rect 214208 150198 214282 150226
rect 214852 150198 214926 150226
rect 215404 150210 215432 157762
rect 215484 156732 215536 156738
rect 215484 156674 215536 156680
rect 215496 150226 215524 156674
rect 215680 154562 215708 163200
rect 216508 155242 216536 163200
rect 217336 160070 217364 163200
rect 217324 160064 217376 160070
rect 217324 160006 217376 160012
rect 218256 159798 218284 163200
rect 216772 159792 216824 159798
rect 216772 159734 216824 159740
rect 218244 159792 218296 159798
rect 218244 159734 218296 159740
rect 216680 159112 216732 159118
rect 216680 159054 216732 159060
rect 216692 156738 216720 159054
rect 216680 156732 216732 156738
rect 216680 156674 216732 156680
rect 216496 155236 216548 155242
rect 216496 155178 216548 155184
rect 215668 154556 215720 154562
rect 215668 154498 215720 154504
rect 216784 153066 216812 159734
rect 218060 156664 218112 156670
rect 218060 156606 218112 156612
rect 217416 154080 217468 154086
rect 217416 154022 217468 154028
rect 216772 153060 216824 153066
rect 216772 153002 216824 153008
rect 216772 152176 216824 152182
rect 216772 152118 216824 152124
rect 216784 150226 216812 152118
rect 217428 150226 217456 154022
rect 218072 150226 218100 156606
rect 219084 155174 219112 163200
rect 219532 155304 219584 155310
rect 219532 155246 219584 155252
rect 219072 155168 219124 155174
rect 219072 155110 219124 155116
rect 218702 152552 218758 152561
rect 218702 152487 218758 152496
rect 218716 150226 218744 152487
rect 219544 151814 219572 155246
rect 219912 154086 219940 163200
rect 220176 159928 220228 159934
rect 220176 159870 220228 159876
rect 220188 158710 220216 159870
rect 220740 158778 220768 163200
rect 220728 158772 220780 158778
rect 220728 158714 220780 158720
rect 220176 158704 220228 158710
rect 220176 158646 220228 158652
rect 220636 158024 220688 158030
rect 220636 157966 220688 157972
rect 219900 154080 219952 154086
rect 219900 154022 219952 154028
rect 219544 151786 220032 151814
rect 219348 151768 219400 151774
rect 219348 151710 219400 151716
rect 211632 150062 211706 150090
rect 211678 149940 211706 150062
rect 212322 149940 212350 150198
rect 212966 149940 212994 150198
rect 213610 149940 213638 150198
rect 214254 149940 214282 150198
rect 214898 149940 214926 150198
rect 215392 150204 215444 150210
rect 215496 150198 215570 150226
rect 215392 150146 215444 150152
rect 215542 149940 215570 150198
rect 216174 150204 216226 150210
rect 216784 150198 216858 150226
rect 217428 150198 217502 150226
rect 218072 150198 218146 150226
rect 218716 150198 218790 150226
rect 216174 150146 216226 150152
rect 216186 149940 216214 150146
rect 216830 149940 216858 150198
rect 217474 149940 217502 150198
rect 218118 149940 218146 150198
rect 218762 149940 218790 150198
rect 219360 150090 219388 151710
rect 220004 150226 220032 151786
rect 220004 150198 220078 150226
rect 219360 150062 219434 150090
rect 219406 149940 219434 150062
rect 220050 149940 220078 150198
rect 220648 150192 220676 157966
rect 221568 157894 221596 163200
rect 221924 159996 221976 160002
rect 221924 159938 221976 159944
rect 221556 157888 221608 157894
rect 221556 157830 221608 157836
rect 221280 152516 221332 152522
rect 221280 152458 221332 152464
rect 221292 150192 221320 152458
rect 221936 152454 221964 159938
rect 222396 159934 222424 163200
rect 222384 159928 222436 159934
rect 222384 159870 222436 159876
rect 222108 159248 222160 159254
rect 222108 159190 222160 159196
rect 222016 155440 222068 155446
rect 222016 155382 222068 155388
rect 222028 152794 222056 155382
rect 222016 152788 222068 152794
rect 222016 152730 222068 152736
rect 222120 152561 222148 159190
rect 222752 156800 222804 156806
rect 222752 156742 222804 156748
rect 222568 153944 222620 153950
rect 222568 153886 222620 153892
rect 222106 152552 222162 152561
rect 222106 152487 222162 152496
rect 221924 152448 221976 152454
rect 221924 152390 221976 152396
rect 221924 152244 221976 152250
rect 221924 152186 221976 152192
rect 221936 150192 221964 152186
rect 222580 150192 222608 153886
rect 222764 151814 222792 156742
rect 223224 155310 223252 163200
rect 223488 160064 223540 160070
rect 223488 160006 223540 160012
rect 223212 155304 223264 155310
rect 223212 155246 223264 155252
rect 223500 153785 223528 160006
rect 224144 158982 224172 163200
rect 224972 159730 225000 163200
rect 225696 159928 225748 159934
rect 225696 159870 225748 159876
rect 224592 159724 224644 159730
rect 224592 159666 224644 159672
rect 224960 159724 225012 159730
rect 224960 159666 225012 159672
rect 224132 158976 224184 158982
rect 224132 158918 224184 158924
rect 223856 157752 223908 157758
rect 223856 157694 223908 157700
rect 223486 153776 223542 153785
rect 223486 153711 223542 153720
rect 222764 151786 223252 151814
rect 223224 150226 223252 151786
rect 223224 150198 223298 150226
rect 220648 150164 220722 150192
rect 221292 150164 221366 150192
rect 221936 150164 222010 150192
rect 222580 150164 222654 150192
rect 220694 149940 220722 150164
rect 221338 149940 221366 150164
rect 221982 149940 222010 150164
rect 222626 149940 222654 150164
rect 223270 149940 223298 150198
rect 223868 150192 223896 157694
rect 224604 152794 224632 159666
rect 224960 158092 225012 158098
rect 224960 158034 225012 158040
rect 224500 152788 224552 152794
rect 224500 152730 224552 152736
rect 224592 152788 224644 152794
rect 224592 152730 224644 152736
rect 224512 150192 224540 152730
rect 224972 150210 225000 158034
rect 225708 158030 225736 159870
rect 225696 158024 225748 158030
rect 225696 157966 225748 157972
rect 225800 155446 225828 163200
rect 225788 155440 225840 155446
rect 225788 155382 225840 155388
rect 226628 155106 226656 163200
rect 227076 160608 227128 160614
rect 227076 160550 227128 160556
rect 226616 155100 226668 155106
rect 226616 155042 226668 155048
rect 225144 154964 225196 154970
rect 225144 154906 225196 154912
rect 224960 150204 225012 150210
rect 223868 150164 223942 150192
rect 224512 150164 224586 150192
rect 223914 149940 223942 150164
rect 224558 149940 224586 150164
rect 225156 150192 225184 154906
rect 226432 152312 226484 152318
rect 226432 152254 226484 152260
rect 225834 150204 225886 150210
rect 225156 150164 225230 150192
rect 224960 150146 225012 150152
rect 225202 149940 225230 150164
rect 226444 150192 226472 152254
rect 227088 150192 227116 160550
rect 227456 159254 227484 163200
rect 228284 160070 228312 163200
rect 228272 160064 228324 160070
rect 228272 160006 228324 160012
rect 227444 159248 227496 159254
rect 227444 159190 227496 159196
rect 227720 158976 227772 158982
rect 227720 158918 227772 158924
rect 227732 156534 227760 158918
rect 227904 158772 227956 158778
rect 227904 158714 227956 158720
rect 227720 156528 227772 156534
rect 227720 156470 227772 156476
rect 227916 155281 227944 158714
rect 229112 158098 229140 163200
rect 229100 158092 229152 158098
rect 229100 158034 229152 158040
rect 230032 155582 230060 163200
rect 230388 159860 230440 159866
rect 230388 159802 230440 159808
rect 229192 155576 229244 155582
rect 229192 155518 229244 155524
rect 230020 155576 230072 155582
rect 230020 155518 230072 155524
rect 227718 155272 227774 155281
rect 227718 155207 227774 155216
rect 227902 155272 227958 155281
rect 227902 155207 227958 155216
rect 227732 150192 227760 155207
rect 228364 154012 228416 154018
rect 228364 153954 228416 153960
rect 228376 150192 228404 153954
rect 229008 152856 229060 152862
rect 229008 152798 229060 152804
rect 229020 150226 229048 152798
rect 229020 150198 229094 150226
rect 229204 150210 229232 155518
rect 230400 152250 230428 159802
rect 230664 159316 230716 159322
rect 230664 159258 230716 159264
rect 230676 152318 230704 159258
rect 230860 158778 230888 163200
rect 231688 159866 231716 163200
rect 232228 160744 232280 160750
rect 232228 160686 232280 160692
rect 231952 160540 232004 160546
rect 231952 160482 232004 160488
rect 231676 159860 231728 159866
rect 231676 159802 231728 159808
rect 230848 158772 230900 158778
rect 230848 158714 230900 158720
rect 230940 155372 230992 155378
rect 230940 155314 230992 155320
rect 230664 152312 230716 152318
rect 230664 152254 230716 152260
rect 230388 152244 230440 152250
rect 230388 152186 230440 152192
rect 229652 151020 229704 151026
rect 229652 150962 229704 150968
rect 226444 150164 226518 150192
rect 227088 150164 227162 150192
rect 227732 150164 227806 150192
rect 228376 150164 228450 150192
rect 225834 150146 225886 150152
rect 225846 149940 225874 150146
rect 226490 149940 226518 150164
rect 227134 149940 227162 150164
rect 227778 149940 227806 150164
rect 228422 149940 228450 150164
rect 229066 149940 229094 150198
rect 229192 150204 229244 150210
rect 229192 150146 229244 150152
rect 229664 150090 229692 150962
rect 230952 150226 230980 155314
rect 231584 152584 231636 152590
rect 231584 152526 231636 152532
rect 231596 150226 231624 152526
rect 230342 150204 230394 150210
rect 230952 150198 231026 150226
rect 231596 150198 231670 150226
rect 231964 150210 231992 160482
rect 232240 150226 232268 160686
rect 232516 155378 232544 163200
rect 233240 157956 233292 157962
rect 233240 157898 233292 157904
rect 232504 155372 232556 155378
rect 232504 155314 232556 155320
rect 230342 150146 230394 150152
rect 229664 150062 229738 150090
rect 229710 149940 229738 150062
rect 230354 149940 230382 150146
rect 230998 149940 231026 150198
rect 231642 149940 231670 150198
rect 231952 150204 232004 150210
rect 232240 150198 232314 150226
rect 233252 150210 233280 157898
rect 233344 153950 233372 163200
rect 234172 160002 234200 163200
rect 234160 159996 234212 160002
rect 234160 159938 234212 159944
rect 233516 156868 233568 156874
rect 233516 156810 233568 156816
rect 233332 153944 233384 153950
rect 233332 153886 233384 153892
rect 233528 150226 233556 156810
rect 235000 152522 235028 163200
rect 235920 158137 235948 163200
rect 235998 159352 236054 159361
rect 235998 159287 236054 159296
rect 235906 158128 235962 158137
rect 235906 158063 235962 158072
rect 234988 152516 235040 152522
rect 234988 152458 235040 152464
rect 236012 151910 236040 159287
rect 236092 158160 236144 158166
rect 236092 158102 236144 158108
rect 236000 151904 236052 151910
rect 236000 151846 236052 151852
rect 234804 151088 234856 151094
rect 234804 151030 234856 151036
rect 231952 150146 232004 150152
rect 232286 149940 232314 150198
rect 232918 150204 232970 150210
rect 232918 150146 232970 150152
rect 233240 150204 233292 150210
rect 233528 150198 233602 150226
rect 233240 150146 233292 150152
rect 232930 149940 232958 150146
rect 233574 149940 233602 150198
rect 234206 150204 234258 150210
rect 234206 150146 234258 150152
rect 234218 149940 234246 150146
rect 234816 150090 234844 151030
rect 235448 150952 235500 150958
rect 235448 150894 235500 150900
rect 235460 150090 235488 150894
rect 236104 150226 236132 158102
rect 236748 156806 236776 163200
rect 237380 160812 237432 160818
rect 237380 160754 237432 160760
rect 236736 156800 236788 156806
rect 236736 156742 236788 156748
rect 236736 152380 236788 152386
rect 236736 152322 236788 152328
rect 236748 150226 236776 152322
rect 237392 150226 237420 160754
rect 237576 159322 237604 163200
rect 238404 159934 238432 163200
rect 238392 159928 238444 159934
rect 238392 159870 238444 159876
rect 237564 159316 237616 159322
rect 237564 159258 237616 159264
rect 238668 158772 238720 158778
rect 238668 158714 238720 158720
rect 238680 155514 238708 158714
rect 239232 157962 239260 163200
rect 239956 160064 240008 160070
rect 239956 160006 240008 160012
rect 239220 157956 239272 157962
rect 239220 157898 239272 157904
rect 238576 155508 238628 155514
rect 238576 155450 238628 155456
rect 238668 155508 238720 155514
rect 238668 155450 238720 155456
rect 238024 153604 238076 153610
rect 238024 153546 238076 153552
rect 238036 150226 238064 153546
rect 238588 151814 238616 155450
rect 239968 153066 239996 160006
rect 240060 156670 240088 163200
rect 240888 160070 240916 163200
rect 240876 160064 240928 160070
rect 240876 160006 240928 160012
rect 241704 159452 241756 159458
rect 241704 159394 241756 159400
rect 241244 156936 241296 156942
rect 241244 156878 241296 156884
rect 240048 156664 240100 156670
rect 240048 156606 240100 156612
rect 239312 153060 239364 153066
rect 239312 153002 239364 153008
rect 239956 153060 240008 153066
rect 239956 153002 240008 153008
rect 238588 151786 238708 151814
rect 238680 150226 238708 151786
rect 239324 150226 239352 153002
rect 240600 151904 240652 151910
rect 240600 151846 240652 151852
rect 239956 151156 240008 151162
rect 239956 151098 240008 151104
rect 236104 150198 236178 150226
rect 236748 150198 236822 150226
rect 237392 150198 237466 150226
rect 238036 150198 238110 150226
rect 238680 150198 238754 150226
rect 239324 150198 239398 150226
rect 234816 150062 234890 150090
rect 235460 150062 235534 150090
rect 234862 149940 234890 150062
rect 235506 149940 235534 150062
rect 236150 149940 236178 150198
rect 236794 149940 236822 150198
rect 237438 149940 237466 150198
rect 238082 149940 238110 150198
rect 238726 149940 238754 150198
rect 239370 149940 239398 150198
rect 239968 150090 239996 151098
rect 240612 150226 240640 151846
rect 241256 150226 241284 156878
rect 241716 152182 241744 159394
rect 241808 158778 241836 163200
rect 242072 160880 242124 160886
rect 242072 160822 242124 160828
rect 241796 158772 241848 158778
rect 241796 158714 241848 158720
rect 241886 152416 241942 152425
rect 241886 152351 241942 152360
rect 241704 152176 241756 152182
rect 241704 152118 241756 152124
rect 241900 150226 241928 152351
rect 242084 151814 242112 160822
rect 242636 158166 242664 163200
rect 242900 158228 242952 158234
rect 242900 158170 242952 158176
rect 242624 158160 242676 158166
rect 242624 158102 242676 158108
rect 242084 151786 242480 151814
rect 242452 150226 242480 151786
rect 240612 150198 240686 150226
rect 241256 150198 241330 150226
rect 241900 150198 241974 150226
rect 242452 150198 242526 150226
rect 242912 150210 242940 158170
rect 243082 156632 243138 156641
rect 243082 156567 243138 156576
rect 243096 150226 243124 156567
rect 243464 154018 243492 163200
rect 243452 154012 243504 154018
rect 243452 153954 243504 153960
rect 244292 153746 244320 163200
rect 245120 159458 245148 163200
rect 245752 160948 245804 160954
rect 245752 160890 245804 160896
rect 245108 159452 245160 159458
rect 245108 159394 245160 159400
rect 244648 158772 244700 158778
rect 244648 158714 244700 158720
rect 244280 153740 244332 153746
rect 244280 153682 244332 153688
rect 244660 152862 244688 158714
rect 245660 157888 245712 157894
rect 245660 157830 245712 157836
rect 244648 152856 244700 152862
rect 244648 152798 244700 152804
rect 245672 152454 245700 157830
rect 244372 152448 244424 152454
rect 244372 152390 244424 152396
rect 245660 152448 245712 152454
rect 245660 152390 245712 152396
rect 244384 150226 244412 152390
rect 245016 151292 245068 151298
rect 245016 151234 245068 151240
rect 239968 150062 240042 150090
rect 240014 149940 240042 150062
rect 240658 149940 240686 150198
rect 241302 149940 241330 150198
rect 241946 149940 241974 150198
rect 242498 149940 242526 150198
rect 242900 150204 242952 150210
rect 243096 150198 243170 150226
rect 242900 150146 242952 150152
rect 243142 149940 243170 150198
rect 243774 150204 243826 150210
rect 244384 150198 244458 150226
rect 243774 150146 243826 150152
rect 243786 149940 243814 150146
rect 244430 149940 244458 150198
rect 245028 150090 245056 151234
rect 245764 150226 245792 160890
rect 245948 158234 245976 163200
rect 245936 158228 245988 158234
rect 245936 158170 245988 158176
rect 246776 156874 246804 163200
rect 247224 159520 247276 159526
rect 247224 159462 247276 159468
rect 247040 159248 247092 159254
rect 247040 159190 247092 159196
rect 246764 156868 246816 156874
rect 246764 156810 246816 156816
rect 247052 156641 247080 159190
rect 247132 157004 247184 157010
rect 247132 156946 247184 156952
rect 247038 156632 247094 156641
rect 247038 156567 247094 156576
rect 246948 152652 247000 152658
rect 246948 152594 247000 152600
rect 246304 151224 246356 151230
rect 246304 151166 246356 151172
rect 245718 150198 245792 150226
rect 245028 150062 245102 150090
rect 245074 149940 245102 150062
rect 245718 149940 245746 150198
rect 246316 150090 246344 151166
rect 246960 150226 246988 152594
rect 246960 150198 247034 150226
rect 247144 150210 247172 156946
rect 247236 152386 247264 159462
rect 247696 159118 247724 163200
rect 247684 159112 247736 159118
rect 247684 159054 247736 159060
rect 247592 153128 247644 153134
rect 247592 153070 247644 153076
rect 247224 152380 247276 152386
rect 247224 152322 247276 152328
rect 247604 150226 247632 153070
rect 248524 152590 248552 163200
rect 249352 156942 249380 163200
rect 250180 161474 250208 163200
rect 250180 161446 250300 161474
rect 249340 156936 249392 156942
rect 249340 156878 249392 156884
rect 248880 156460 248932 156466
rect 248880 156402 248932 156408
rect 248512 152584 248564 152590
rect 248512 152526 248564 152532
rect 248892 150226 248920 156402
rect 250272 154154 250300 161446
rect 251008 159254 251036 163200
rect 251836 159526 251864 163200
rect 251824 159520 251876 159526
rect 251824 159462 251876 159468
rect 251732 159316 251784 159322
rect 251732 159258 251784 159264
rect 250996 159248 251048 159254
rect 250996 159190 251048 159196
rect 251456 158296 251508 158302
rect 251456 158238 251508 158244
rect 250812 157140 250864 157146
rect 250812 157082 250864 157088
rect 250168 154148 250220 154154
rect 250168 154090 250220 154096
rect 250260 154148 250312 154154
rect 250260 154090 250312 154096
rect 249524 152244 249576 152250
rect 249524 152186 249576 152192
rect 249536 150226 249564 152186
rect 250180 150226 250208 154090
rect 250824 150226 250852 157082
rect 251468 150226 251496 158238
rect 251744 156466 251772 159258
rect 252664 158302 252692 163200
rect 252744 161016 252796 161022
rect 252744 160958 252796 160964
rect 252652 158296 252704 158302
rect 252652 158238 252704 158244
rect 252008 157956 252060 157962
rect 252008 157898 252060 157904
rect 251732 156460 251784 156466
rect 251732 156402 251784 156408
rect 252020 153134 252048 157898
rect 252560 157072 252612 157078
rect 252560 157014 252612 157020
rect 252100 153196 252152 153202
rect 252100 153138 252152 153144
rect 252008 153128 252060 153134
rect 252008 153070 252060 153076
rect 252112 150226 252140 153138
rect 246316 150062 246390 150090
rect 246362 149940 246390 150062
rect 247006 149940 247034 150198
rect 247132 150204 247184 150210
rect 247604 150198 247678 150226
rect 247132 150146 247184 150152
rect 247650 149940 247678 150198
rect 248282 150204 248334 150210
rect 248892 150198 248966 150226
rect 249536 150198 249610 150226
rect 250180 150198 250254 150226
rect 250824 150198 250898 150226
rect 251468 150198 251542 150226
rect 252112 150198 252186 150226
rect 252572 150210 252600 157014
rect 252756 150226 252784 160958
rect 253584 157010 253612 163200
rect 254032 158364 254084 158370
rect 254032 158306 254084 158312
rect 253572 157004 253624 157010
rect 253572 156946 253624 156952
rect 254044 150226 254072 158306
rect 254412 157078 254440 163200
rect 254400 157072 254452 157078
rect 254400 157014 254452 157020
rect 255240 152658 255268 163200
rect 255504 159996 255556 160002
rect 255504 159938 255556 159944
rect 255516 153921 255544 159938
rect 256068 158370 256096 163200
rect 256896 158778 256924 163200
rect 257344 159384 257396 159390
rect 257344 159326 257396 159332
rect 256884 158772 256936 158778
rect 256884 158714 256936 158720
rect 256056 158364 256108 158370
rect 256056 158306 256108 158312
rect 255872 157276 255924 157282
rect 255872 157218 255924 157224
rect 255318 153912 255374 153921
rect 255318 153847 255374 153856
rect 255502 153912 255558 153921
rect 255502 153847 255558 153856
rect 255228 152652 255280 152658
rect 255228 152594 255280 152600
rect 254676 152176 254728 152182
rect 254676 152118 254728 152124
rect 254688 150226 254716 152118
rect 255332 150226 255360 153847
rect 255884 151814 255912 157218
rect 257356 152318 257384 159326
rect 257724 159186 257752 163200
rect 258080 161084 258132 161090
rect 258080 161026 258132 161032
rect 257712 159180 257764 159186
rect 257712 159122 257764 159128
rect 257988 158772 258040 158778
rect 257988 158714 258040 158720
rect 258000 154222 258028 158714
rect 257896 154216 257948 154222
rect 257896 154158 257948 154164
rect 257988 154216 258040 154222
rect 257988 154158 258040 154164
rect 257252 152312 257304 152318
rect 257252 152254 257304 152260
rect 257344 152312 257396 152318
rect 257344 152254 257396 152260
rect 255884 151786 256004 151814
rect 255976 150226 256004 151786
rect 256608 151360 256660 151366
rect 256608 151302 256660 151308
rect 248282 150146 248334 150152
rect 248294 149940 248322 150146
rect 248938 149940 248966 150198
rect 249582 149940 249610 150198
rect 250226 149940 250254 150198
rect 250870 149940 250898 150198
rect 251514 149940 251542 150198
rect 252158 149940 252186 150198
rect 252560 150204 252612 150210
rect 252756 150198 252830 150226
rect 252560 150146 252612 150152
rect 252802 149940 252830 150198
rect 253434 150204 253486 150210
rect 254044 150198 254118 150226
rect 254688 150198 254762 150226
rect 255332 150198 255406 150226
rect 255976 150198 256050 150226
rect 253434 150146 253486 150152
rect 253446 149940 253474 150146
rect 254090 149940 254118 150198
rect 254734 149940 254762 150198
rect 255378 149940 255406 150198
rect 256022 149940 256050 150198
rect 256620 150090 256648 151302
rect 257264 150226 257292 152254
rect 257908 150226 257936 154158
rect 257264 150198 257338 150226
rect 257908 150198 257982 150226
rect 258092 150210 258120 161026
rect 258552 160002 258580 163200
rect 258540 159996 258592 160002
rect 258540 159938 258592 159944
rect 259472 157962 259500 163200
rect 259644 159588 259696 159594
rect 259644 159530 259696 159536
rect 259460 157956 259512 157962
rect 259460 157898 259512 157904
rect 258538 156768 258594 156777
rect 258538 156703 258594 156712
rect 258552 150226 258580 156703
rect 259656 153202 259684 159530
rect 260300 157146 260328 163200
rect 261128 158778 261156 163200
rect 261956 158846 261984 163200
rect 262128 159112 262180 159118
rect 262128 159054 262180 159060
rect 261944 158840 261996 158846
rect 261944 158782 261996 158788
rect 261116 158772 261168 158778
rect 261116 158714 261168 158720
rect 260840 158432 260892 158438
rect 260840 158374 260892 158380
rect 260288 157140 260340 157146
rect 260288 157082 260340 157088
rect 260472 154352 260524 154358
rect 260472 154294 260524 154300
rect 259644 153196 259696 153202
rect 259644 153138 259696 153144
rect 259828 152380 259880 152386
rect 259828 152322 259880 152328
rect 259840 150226 259868 152322
rect 260484 150226 260512 154294
rect 256620 150062 256694 150090
rect 256666 149940 256694 150062
rect 257310 149940 257338 150198
rect 257954 149940 257982 150198
rect 258080 150204 258132 150210
rect 258552 150198 258626 150226
rect 258080 150146 258132 150152
rect 258598 149940 258626 150198
rect 259230 150204 259282 150210
rect 259840 150198 259914 150226
rect 260484 150198 260558 150226
rect 260852 150210 260880 158374
rect 261116 155644 261168 155650
rect 261116 155586 261168 155592
rect 261128 150226 261156 155586
rect 262140 154970 262168 159054
rect 262784 158438 262812 163200
rect 263416 158840 263468 158846
rect 263416 158782 263468 158788
rect 262772 158432 262824 158438
rect 262772 158374 262824 158380
rect 262128 154964 262180 154970
rect 262128 154906 262180 154912
rect 263048 154284 263100 154290
rect 263048 154226 263100 154232
rect 262404 152924 262456 152930
rect 262404 152866 262456 152872
rect 262416 150226 262444 152866
rect 263060 150226 263088 154226
rect 263428 152930 263456 158782
rect 263612 154290 263640 163200
rect 263876 160064 263928 160070
rect 263876 160006 263928 160012
rect 263784 158500 263836 158506
rect 263784 158442 263836 158448
rect 263690 155408 263746 155417
rect 263690 155343 263746 155352
rect 263600 154284 263652 154290
rect 263600 154226 263652 154232
rect 263600 153672 263652 153678
rect 263600 153614 263652 153620
rect 263416 152924 263468 152930
rect 263416 152866 263468 152872
rect 259230 150146 259282 150152
rect 259242 149940 259270 150146
rect 259886 149940 259914 150198
rect 260530 149940 260558 150198
rect 260840 150204 260892 150210
rect 261128 150198 261202 150226
rect 260840 150146 260892 150152
rect 261174 149940 261202 150198
rect 261806 150204 261858 150210
rect 262416 150198 262490 150226
rect 263060 150198 263134 150226
rect 263612 150210 263640 153614
rect 263704 150226 263732 155343
rect 263796 153678 263824 158442
rect 263888 155417 263916 160006
rect 264440 159118 264468 163200
rect 265360 160070 265388 163200
rect 265348 160064 265400 160070
rect 265348 160006 265400 160012
rect 265070 159488 265126 159497
rect 265070 159423 265126 159432
rect 264428 159112 264480 159118
rect 264428 159054 264480 159060
rect 263874 155408 263930 155417
rect 263874 155343 263930 155352
rect 263784 153672 263836 153678
rect 263784 153614 263836 153620
rect 265084 152318 265112 159423
rect 266188 158506 266216 163200
rect 266176 158500 266228 158506
rect 266176 158442 266228 158448
rect 266912 157344 266964 157350
rect 266912 157286 266964 157292
rect 265164 155712 265216 155718
rect 265164 155654 265216 155660
rect 264980 152312 265032 152318
rect 264980 152254 265032 152260
rect 265072 152312 265124 152318
rect 265072 152254 265124 152260
rect 264992 150226 265020 152254
rect 261806 150146 261858 150152
rect 261818 149940 261846 150146
rect 262462 149940 262490 150198
rect 263106 149940 263134 150198
rect 263600 150204 263652 150210
rect 263704 150198 263778 150226
rect 263600 150146 263652 150152
rect 263750 149940 263778 150198
rect 264382 150204 264434 150210
rect 264992 150198 265066 150226
rect 265176 150210 265204 155654
rect 265716 154420 265768 154426
rect 265716 154362 265768 154368
rect 265728 150226 265756 154362
rect 264382 150146 264434 150152
rect 264394 149940 264422 150146
rect 265038 149940 265066 150198
rect 265164 150204 265216 150210
rect 265164 150146 265216 150152
rect 265682 150198 265756 150226
rect 266924 150226 266952 157286
rect 267016 154426 267044 163200
rect 267844 159050 267872 163200
rect 267832 159044 267884 159050
rect 267832 158986 267884 158992
rect 268672 158846 268700 163200
rect 268936 159656 268988 159662
rect 268936 159598 268988 159604
rect 268660 158840 268712 158846
rect 268660 158782 268712 158788
rect 268844 154488 268896 154494
rect 268844 154430 268896 154436
rect 267004 154420 267056 154426
rect 267004 154362 267056 154368
rect 267556 152992 267608 152998
rect 267556 152934 267608 152940
rect 267568 150226 267596 152934
rect 268200 151428 268252 151434
rect 268200 151370 268252 151376
rect 266314 150204 266366 150210
rect 265682 149940 265710 150198
rect 266924 150198 266998 150226
rect 267568 150198 267642 150226
rect 266314 150146 266366 150152
rect 266326 149940 266354 150146
rect 266970 149940 266998 150198
rect 267614 149940 267642 150198
rect 268212 150090 268240 151370
rect 268856 150226 268884 154430
rect 268948 152386 268976 159598
rect 269028 158772 269080 158778
rect 269028 158714 269080 158720
rect 269040 155038 269068 158714
rect 269396 158568 269448 158574
rect 269396 158510 269448 158516
rect 269028 155032 269080 155038
rect 269028 154974 269080 154980
rect 268936 152380 268988 152386
rect 268936 152322 268988 152328
rect 269408 151814 269436 158510
rect 269500 157894 269528 163200
rect 269488 157888 269540 157894
rect 269488 157830 269540 157836
rect 270328 154358 270356 163200
rect 270500 161152 270552 161158
rect 270500 161094 270552 161100
rect 270316 154352 270368 154358
rect 270316 154294 270368 154300
rect 270132 153196 270184 153202
rect 270132 153138 270184 153144
rect 269408 151786 269528 151814
rect 269500 150226 269528 151786
rect 270144 150226 270172 153138
rect 270512 151814 270540 161094
rect 271248 159322 271276 163200
rect 272076 159594 272104 163200
rect 272524 159792 272576 159798
rect 272524 159734 272576 159740
rect 272064 159588 272116 159594
rect 272064 159530 272116 159536
rect 271236 159316 271288 159322
rect 271236 159258 271288 159264
rect 271696 158840 271748 158846
rect 271696 158782 271748 158788
rect 271052 155780 271104 155786
rect 271052 155722 271104 155728
rect 271064 151814 271092 155722
rect 271708 152998 271736 158782
rect 272064 158636 272116 158642
rect 272064 158578 272116 158584
rect 271696 152992 271748 152998
rect 271696 152934 271748 152940
rect 270512 151786 270816 151814
rect 271064 151786 271460 151814
rect 270788 150226 270816 151786
rect 271432 150226 271460 151786
rect 272076 150226 272104 158578
rect 272536 153202 272564 159734
rect 272904 158574 272932 163200
rect 272892 158568 272944 158574
rect 272892 158510 272944 158516
rect 273444 155916 273496 155922
rect 273444 155858 273496 155864
rect 272524 153196 272576 153202
rect 272524 153138 272576 153144
rect 272708 152720 272760 152726
rect 272708 152662 272760 152668
rect 272720 150226 272748 152662
rect 273260 151496 273312 151502
rect 273260 151438 273312 151444
rect 268856 150198 268930 150226
rect 269500 150198 269574 150226
rect 270144 150198 270218 150226
rect 270788 150198 270862 150226
rect 271432 150198 271506 150226
rect 272076 150198 272150 150226
rect 272720 150198 272794 150226
rect 268212 150062 268286 150090
rect 268258 149940 268286 150062
rect 268902 149940 268930 150198
rect 269546 149940 269574 150198
rect 270190 149940 270218 150198
rect 270834 149940 270862 150198
rect 271478 149940 271506 150198
rect 272122 149940 272150 150198
rect 272766 149940 272794 150198
rect 273272 150090 273300 151438
rect 273456 150210 273484 155858
rect 273732 155650 273760 163200
rect 274560 158642 274588 163200
rect 275192 161220 275244 161226
rect 275192 161162 275244 161168
rect 274640 159248 274692 159254
rect 274640 159190 274692 159196
rect 274548 158636 274600 158642
rect 274548 158578 274600 158584
rect 273720 155644 273772 155650
rect 273720 155586 273772 155592
rect 274652 154494 274680 159190
rect 274640 154488 274692 154494
rect 274640 154430 274692 154436
rect 273904 153808 273956 153814
rect 273904 153750 273956 153756
rect 273916 150226 273944 153750
rect 275100 152312 275152 152318
rect 275100 152254 275152 152260
rect 275112 150498 275140 152254
rect 275204 151814 275232 161162
rect 275388 158914 275416 163200
rect 275376 158908 275428 158914
rect 275376 158850 275428 158856
rect 276018 157992 276074 158001
rect 276018 157927 276074 157936
rect 275204 151786 275876 151814
rect 275112 150470 275232 150498
rect 275204 150226 275232 150470
rect 275848 150226 275876 151786
rect 273444 150204 273496 150210
rect 273916 150198 273990 150226
rect 273444 150146 273496 150152
rect 273272 150062 273346 150090
rect 273318 149940 273346 150062
rect 273962 149940 273990 150198
rect 274594 150204 274646 150210
rect 275204 150198 275278 150226
rect 275848 150198 275922 150226
rect 276032 150210 276060 157927
rect 276216 157282 276244 163200
rect 276204 157276 276256 157282
rect 276204 157218 276256 157224
rect 276480 155848 276532 155854
rect 276480 155790 276532 155796
rect 276492 150226 276520 155790
rect 277136 155718 277164 163200
rect 277964 159798 277992 163200
rect 277952 159792 278004 159798
rect 277952 159734 278004 159740
rect 278792 158982 278820 163200
rect 279516 159044 279568 159050
rect 279516 158986 279568 158992
rect 278780 158976 278832 158982
rect 278780 158918 278832 158924
rect 278320 158908 278372 158914
rect 278320 158850 278372 158856
rect 277952 158704 278004 158710
rect 277952 158646 278004 158652
rect 277124 155712 277176 155718
rect 277124 155654 277176 155660
rect 277766 152552 277822 152561
rect 277766 152487 277822 152496
rect 277780 150226 277808 152487
rect 277964 151814 277992 158646
rect 278332 152726 278360 158850
rect 279056 157208 279108 157214
rect 279056 157150 279108 157156
rect 278780 156596 278832 156602
rect 278780 156538 278832 156544
rect 278320 152720 278372 152726
rect 278320 152662 278372 152668
rect 277964 151786 278452 151814
rect 278424 150226 278452 151786
rect 274594 150146 274646 150152
rect 274606 149940 274634 150146
rect 275250 149940 275278 150198
rect 275894 149940 275922 150198
rect 276020 150204 276072 150210
rect 276492 150198 276566 150226
rect 276020 150146 276072 150152
rect 276538 149940 276566 150198
rect 277170 150204 277222 150210
rect 277780 150198 277854 150226
rect 278424 150198 278498 150226
rect 278792 150210 278820 156538
rect 279068 150226 279096 157150
rect 279528 156398 279556 158986
rect 279620 158710 279648 163200
rect 280068 159180 280120 159186
rect 280068 159122 280120 159128
rect 279608 158704 279660 158710
rect 279608 158646 279660 158652
rect 279516 156392 279568 156398
rect 279516 156334 279568 156340
rect 280080 153814 280108 159122
rect 280448 155786 280476 163200
rect 281276 158778 281304 163200
rect 282104 159730 282132 163200
rect 281448 159724 281500 159730
rect 281448 159666 281500 159672
rect 282092 159724 282144 159730
rect 282092 159666 282144 159672
rect 281264 158772 281316 158778
rect 281264 158714 281316 158720
rect 280436 155780 280488 155786
rect 280436 155722 280488 155728
rect 280068 153808 280120 153814
rect 280068 153750 280120 153756
rect 280344 152380 280396 152386
rect 280344 152322 280396 152328
rect 280356 150226 280384 152322
rect 281460 152318 281488 159666
rect 282552 158772 282604 158778
rect 282552 158714 282604 158720
rect 282092 156732 282144 156738
rect 282092 156674 282144 156680
rect 281632 153876 281684 153882
rect 281632 153818 281684 153824
rect 281448 152312 281500 152318
rect 281448 152254 281500 152260
rect 280988 151564 281040 151570
rect 280988 151506 281040 151512
rect 277170 150146 277222 150152
rect 277182 149940 277210 150146
rect 277826 149940 277854 150198
rect 278470 149940 278498 150198
rect 278780 150204 278832 150210
rect 279068 150198 279142 150226
rect 278780 150146 278832 150152
rect 279114 149940 279142 150198
rect 279746 150204 279798 150210
rect 280356 150198 280430 150226
rect 279746 150146 279798 150152
rect 279758 149940 279786 150146
rect 280402 149940 280430 150198
rect 281000 150090 281028 151506
rect 281644 150226 281672 153818
rect 282104 151814 282132 156674
rect 282564 153882 282592 158714
rect 283024 156738 283052 163200
rect 283012 156732 283064 156738
rect 283012 156674 283064 156680
rect 283852 155242 283880 163200
rect 284392 159860 284444 159866
rect 284392 159802 284444 159808
rect 284300 159112 284352 159118
rect 284300 159054 284352 159060
rect 283104 155236 283156 155242
rect 283104 155178 283156 155184
rect 283840 155236 283892 155242
rect 283840 155178 283892 155184
rect 282552 153876 282604 153882
rect 282552 153818 282604 153824
rect 282920 152788 282972 152794
rect 282920 152730 282972 152736
rect 282104 151786 282316 151814
rect 282288 150226 282316 151786
rect 282932 150226 282960 152730
rect 281644 150198 281718 150226
rect 282288 150198 282362 150226
rect 282932 150198 283006 150226
rect 283116 150210 283144 155178
rect 284312 154562 284340 159054
rect 283564 154556 283616 154562
rect 283564 154498 283616 154504
rect 284300 154556 284352 154562
rect 284300 154498 284352 154504
rect 283576 150226 283604 154498
rect 284404 152794 284432 159802
rect 284680 159254 284708 163200
rect 285508 159662 285536 163200
rect 285496 159656 285548 159662
rect 285496 159598 285548 159604
rect 284668 159248 284720 159254
rect 284668 159190 284720 159196
rect 286336 158778 286364 163200
rect 287060 159792 287112 159798
rect 287060 159734 287112 159740
rect 287072 159390 287100 159734
rect 287060 159384 287112 159390
rect 287060 159326 287112 159332
rect 286324 158772 286376 158778
rect 286324 158714 286376 158720
rect 286876 158772 286928 158778
rect 286876 158714 286928 158720
rect 286140 155168 286192 155174
rect 286140 155110 286192 155116
rect 284850 153776 284906 153785
rect 284850 153711 284906 153720
rect 284392 152788 284444 152794
rect 284392 152730 284444 152736
rect 284864 150226 284892 153711
rect 285496 153196 285548 153202
rect 285496 153138 285548 153144
rect 285508 150226 285536 153138
rect 286152 150226 286180 155110
rect 286888 154086 286916 158714
rect 287164 155854 287192 163200
rect 287992 159798 288020 163200
rect 288348 159928 288400 159934
rect 288348 159870 288400 159876
rect 287980 159792 288032 159798
rect 287980 159734 288032 159740
rect 287152 155848 287204 155854
rect 287152 155790 287204 155796
rect 287426 155272 287482 155281
rect 287426 155207 287482 155216
rect 286784 154080 286836 154086
rect 286784 154022 286836 154028
rect 286876 154080 286928 154086
rect 286876 154022 286928 154028
rect 286796 150226 286824 154022
rect 287440 150226 287468 155207
rect 288072 152448 288124 152454
rect 288072 152390 288124 152396
rect 288084 150226 288112 152390
rect 288360 152386 288388 159870
rect 288624 159792 288676 159798
rect 288624 159734 288676 159740
rect 288440 158024 288492 158030
rect 288440 157966 288492 157972
rect 288348 152380 288400 152386
rect 288348 152322 288400 152328
rect 288452 151814 288480 157966
rect 288636 157214 288664 159734
rect 288912 159050 288940 163200
rect 288900 159044 288952 159050
rect 288900 158986 288952 158992
rect 289740 158030 289768 163200
rect 289912 159724 289964 159730
rect 289912 159666 289964 159672
rect 289728 158024 289780 158030
rect 289728 157966 289780 157972
rect 288624 157208 288676 157214
rect 288624 157150 288676 157156
rect 289360 155304 289412 155310
rect 289360 155246 289412 155252
rect 288452 151786 288756 151814
rect 288728 150226 288756 151786
rect 289372 150226 289400 155246
rect 289924 152454 289952 159666
rect 290004 156528 290056 156534
rect 290004 156470 290056 156476
rect 289912 152448 289964 152454
rect 289912 152390 289964 152396
rect 290016 150226 290044 156470
rect 290568 155310 290596 163200
rect 291396 159934 291424 163200
rect 291384 159928 291436 159934
rect 291384 159870 291436 159876
rect 292224 159730 292252 163200
rect 292212 159724 292264 159730
rect 292212 159666 292264 159672
rect 291476 159384 291528 159390
rect 291476 159326 291528 159332
rect 291292 155440 291344 155446
rect 291292 155382 291344 155388
rect 290556 155304 290608 155310
rect 290556 155246 290608 155252
rect 291200 155100 291252 155106
rect 291200 155042 291252 155048
rect 290648 152312 290700 152318
rect 290648 152254 290700 152260
rect 290660 150226 290688 152254
rect 281000 150062 281074 150090
rect 281046 149940 281074 150062
rect 281690 149940 281718 150198
rect 282334 149940 282362 150198
rect 282978 149940 283006 150198
rect 283104 150204 283156 150210
rect 283576 150198 283650 150226
rect 283104 150146 283156 150152
rect 283622 149940 283650 150198
rect 284254 150204 284306 150210
rect 284864 150198 284938 150226
rect 285508 150198 285582 150226
rect 286152 150198 286226 150226
rect 286796 150198 286870 150226
rect 287440 150198 287514 150226
rect 288084 150198 288158 150226
rect 288728 150198 288802 150226
rect 289372 150198 289446 150226
rect 290016 150198 290090 150226
rect 290660 150198 290734 150226
rect 291212 150210 291240 155042
rect 291304 150226 291332 155382
rect 291488 155174 291516 159326
rect 292304 159044 292356 159050
rect 292304 158986 292356 158992
rect 291476 155168 291528 155174
rect 291476 155110 291528 155116
rect 292316 153202 292344 158986
rect 293052 158098 293080 163200
rect 292764 158092 292816 158098
rect 292764 158034 292816 158040
rect 293040 158092 293092 158098
rect 293040 158034 293092 158040
rect 292578 156632 292634 156641
rect 292578 156567 292634 156576
rect 292304 153196 292356 153202
rect 292304 153138 292356 153144
rect 292592 150226 292620 156567
rect 284254 150146 284306 150152
rect 284266 149940 284294 150146
rect 284910 149940 284938 150198
rect 285554 149940 285582 150198
rect 286198 149940 286226 150198
rect 286842 149940 286870 150198
rect 287486 149940 287514 150198
rect 288130 149940 288158 150198
rect 288774 149940 288802 150198
rect 289418 149940 289446 150198
rect 290062 149940 290090 150198
rect 290706 149940 290734 150198
rect 291200 150204 291252 150210
rect 291304 150198 291378 150226
rect 291200 150146 291252 150152
rect 291350 149940 291378 150198
rect 291982 150204 292034 150210
rect 292592 150198 292666 150226
rect 292776 150210 292804 158034
rect 293880 155446 293908 163200
rect 294512 155576 294564 155582
rect 294512 155518 294564 155524
rect 294052 155508 294104 155514
rect 294052 155450 294104 155456
rect 293868 155440 293920 155446
rect 293868 155382 293920 155388
rect 293224 153060 293276 153066
rect 293224 153002 293276 153008
rect 293236 150226 293264 153002
rect 291982 150146 292034 150152
rect 291994 149940 292022 150146
rect 292638 149940 292666 150198
rect 292764 150204 292816 150210
rect 293236 150198 293310 150226
rect 294064 150210 294092 155450
rect 294524 150226 294552 155518
rect 294800 155514 294828 163200
rect 295628 163146 295656 163200
rect 295720 163146 295748 163254
rect 295628 163118 295748 163146
rect 294788 155508 294840 155514
rect 294788 155450 294840 155456
rect 295904 152794 295932 163254
rect 296442 163200 296498 164400
rect 297270 163200 297326 164400
rect 298098 163200 298154 164400
rect 298926 163200 298982 164400
rect 299754 163200 299810 164400
rect 300674 163200 300730 164400
rect 301502 163200 301558 164400
rect 302330 163200 302386 164400
rect 303158 163200 303214 164400
rect 303986 163200 304042 164400
rect 304814 163200 304870 164400
rect 305642 163200 305698 164400
rect 306562 163200 306618 164400
rect 307390 163200 307446 164400
rect 308218 163200 308274 164400
rect 309046 163200 309102 164400
rect 309874 163200 309930 164400
rect 310702 163200 310758 164400
rect 311530 163200 311586 164400
rect 312450 163200 312506 164400
rect 313278 163200 313334 164400
rect 314106 163200 314162 164400
rect 314934 163200 314990 164400
rect 315762 163200 315818 164400
rect 316590 163200 316646 164400
rect 317418 163200 317474 164400
rect 318338 163200 318394 164400
rect 319166 163200 319222 164400
rect 319994 163200 320050 164400
rect 320822 163200 320878 164400
rect 321650 163200 321706 164400
rect 322478 163200 322534 164400
rect 322584 163254 322796 163282
rect 296456 157350 296484 163200
rect 296812 159316 296864 159322
rect 296812 159258 296864 159264
rect 296444 157344 296496 157350
rect 296444 157286 296496 157292
rect 296444 155372 296496 155378
rect 296444 155314 296496 155320
rect 295800 152788 295852 152794
rect 295800 152730 295852 152736
rect 295892 152788 295944 152794
rect 295892 152730 295944 152736
rect 295812 150226 295840 152730
rect 296456 150226 296484 155314
rect 296824 153678 296852 159258
rect 297284 155582 297312 163200
rect 298112 159322 298140 163200
rect 298940 159798 298968 163200
rect 298928 159792 298980 159798
rect 298928 159734 298980 159740
rect 298744 159452 298796 159458
rect 298744 159394 298796 159400
rect 298100 159316 298152 159322
rect 298100 159258 298152 159264
rect 298650 158128 298706 158137
rect 298650 158063 298706 158072
rect 297272 155576 297324 155582
rect 297272 155518 297324 155524
rect 297088 153944 297140 153950
rect 297088 153886 297140 153892
rect 297730 153912 297786 153921
rect 296812 153672 296864 153678
rect 296812 153614 296864 153620
rect 297100 150226 297128 153886
rect 297730 153847 297786 153856
rect 297744 150226 297772 153847
rect 298376 152516 298428 152522
rect 298376 152458 298428 152464
rect 298388 150226 298416 152458
rect 298664 151814 298692 158063
rect 298756 153066 298784 159394
rect 299768 156806 299796 163200
rect 299480 156800 299532 156806
rect 299480 156742 299532 156748
rect 299756 156800 299808 156806
rect 299756 156742 299808 156748
rect 298744 153060 298796 153066
rect 298744 153002 298796 153008
rect 299492 151814 299520 156742
rect 300308 156460 300360 156466
rect 300308 156402 300360 156408
rect 298664 151786 299060 151814
rect 299492 151786 299704 151814
rect 299032 150226 299060 151786
rect 299676 150226 299704 151786
rect 300320 150226 300348 156402
rect 300688 155378 300716 163200
rect 301516 158778 301544 163200
rect 301688 159520 301740 159526
rect 301688 159462 301740 159468
rect 301504 158772 301556 158778
rect 301504 158714 301556 158720
rect 300676 155372 300728 155378
rect 300676 155314 300728 155320
rect 301700 153134 301728 159462
rect 302240 156664 302292 156670
rect 302240 156606 302292 156612
rect 301596 153128 301648 153134
rect 301596 153070 301648 153076
rect 301688 153128 301740 153134
rect 301688 153070 301740 153076
rect 300952 152380 301004 152386
rect 300952 152322 301004 152328
rect 300964 150226 300992 152322
rect 301608 150226 301636 153070
rect 292764 150146 292816 150152
rect 293282 149940 293310 150198
rect 293914 150204 293966 150210
rect 293914 150146 293966 150152
rect 294052 150204 294104 150210
rect 294524 150198 294598 150226
rect 294052 150146 294104 150152
rect 293926 149940 293954 150146
rect 294570 149940 294598 150198
rect 295202 150204 295254 150210
rect 295812 150198 295886 150226
rect 296456 150198 296530 150226
rect 297100 150198 297174 150226
rect 297744 150198 297818 150226
rect 298388 150198 298462 150226
rect 299032 150198 299106 150226
rect 299676 150198 299750 150226
rect 300320 150198 300394 150226
rect 300964 150198 301038 150226
rect 301608 150198 301682 150226
rect 295202 150146 295254 150152
rect 295214 149940 295242 150146
rect 295858 149940 295886 150198
rect 296502 149940 296530 150198
rect 297146 149940 297174 150198
rect 297790 149940 297818 150198
rect 298434 149940 298462 150198
rect 299078 149940 299106 150198
rect 299722 149940 299750 150198
rect 300366 149940 300394 150198
rect 301010 149940 301038 150198
rect 301654 149940 301682 150198
rect 302252 150090 302280 156606
rect 302344 152522 302372 163200
rect 303172 156602 303200 163200
rect 304000 156670 304028 163200
rect 304828 159186 304856 163200
rect 305000 159996 305052 160002
rect 305000 159938 305052 159944
rect 304816 159180 304868 159186
rect 304816 159122 304868 159128
rect 304816 158772 304868 158778
rect 304816 158714 304868 158720
rect 304080 158160 304132 158166
rect 304080 158102 304132 158108
rect 303988 156664 304040 156670
rect 303988 156606 304040 156612
rect 303160 156596 303212 156602
rect 303160 156538 303212 156544
rect 302882 155408 302938 155417
rect 302882 155343 302938 155352
rect 302332 152516 302384 152522
rect 302332 152458 302384 152464
rect 302896 150090 302924 155343
rect 303528 152856 303580 152862
rect 303528 152798 303580 152804
rect 303540 150090 303568 152798
rect 304092 150226 304120 158102
rect 304828 154018 304856 158714
rect 304724 154012 304776 154018
rect 304724 153954 304776 153960
rect 304816 154012 304868 154018
rect 304816 153954 304868 153960
rect 304092 150198 304166 150226
rect 302252 150062 302326 150090
rect 302896 150062 302970 150090
rect 303540 150062 303614 150090
rect 302298 149940 302326 150062
rect 302942 149940 302970 150062
rect 303586 149940 303614 150062
rect 304138 149940 304166 150198
rect 304736 150090 304764 153954
rect 305012 152862 305040 159938
rect 305656 159866 305684 163200
rect 306576 161474 306604 163200
rect 306576 161446 306696 161474
rect 305644 159860 305696 159866
rect 305644 159802 305696 159808
rect 305460 159248 305512 159254
rect 305460 159190 305512 159196
rect 305472 153746 305500 159190
rect 306380 158228 306432 158234
rect 306380 158170 306432 158176
rect 306392 157334 306420 158170
rect 306392 157306 306604 157334
rect 306380 156936 306432 156942
rect 306380 156878 306432 156884
rect 306392 156466 306420 156878
rect 306380 156460 306432 156466
rect 306380 156402 306432 156408
rect 305368 153740 305420 153746
rect 305368 153682 305420 153688
rect 305460 153740 305512 153746
rect 305460 153682 305512 153688
rect 305000 152856 305052 152862
rect 305000 152798 305052 152804
rect 305380 150090 305408 153682
rect 306012 153060 306064 153066
rect 306012 153002 306064 153008
rect 306024 150090 306052 153002
rect 306576 150226 306604 157306
rect 306668 156874 306696 161446
rect 307404 158166 307432 163200
rect 308232 159526 308260 163200
rect 308220 159520 308272 159526
rect 308220 159462 308272 159468
rect 307392 158160 307444 158166
rect 307392 158102 307444 158108
rect 307024 157004 307076 157010
rect 307024 156946 307076 156952
rect 306656 156868 306708 156874
rect 306656 156810 306708 156816
rect 307036 156534 307064 156946
rect 307300 156936 307352 156942
rect 307300 156878 307352 156884
rect 307024 156528 307076 156534
rect 307024 156470 307076 156476
rect 306576 150198 306742 150226
rect 304736 150062 304810 150090
rect 305380 150062 305454 150090
rect 306024 150062 306098 150090
rect 304782 149940 304810 150062
rect 305426 149940 305454 150062
rect 306070 149940 306098 150062
rect 306714 149940 306742 150198
rect 307312 150090 307340 156878
rect 307944 154964 307996 154970
rect 307944 154906 307996 154912
rect 307956 150090 307984 154906
rect 309060 152590 309088 163200
rect 309888 161474 309916 163200
rect 309888 161446 310008 161474
rect 309232 156460 309284 156466
rect 309232 156402 309284 156408
rect 308588 152584 308640 152590
rect 308588 152526 308640 152532
rect 309048 152584 309100 152590
rect 309048 152526 309100 152532
rect 308600 150090 308628 152526
rect 309244 150090 309272 156402
rect 309876 154148 309928 154154
rect 309876 154090 309928 154096
rect 309888 150090 309916 154090
rect 309980 153950 310008 161446
rect 310612 158296 310664 158302
rect 310612 158238 310664 158244
rect 310520 154488 310572 154494
rect 310520 154430 310572 154436
rect 309968 153944 310020 153950
rect 309968 153886 310020 153892
rect 310532 150090 310560 154430
rect 310624 150210 310652 158238
rect 310716 156942 310744 163200
rect 311072 160064 311124 160070
rect 311072 160006 311124 160012
rect 310704 156936 310756 156942
rect 310704 156878 310756 156884
rect 311084 153066 311112 160006
rect 311544 160002 311572 163200
rect 311532 159996 311584 160002
rect 311532 159938 311584 159944
rect 311900 159928 311952 159934
rect 311900 159870 311952 159876
rect 311912 157826 311940 159870
rect 312464 159458 312492 163200
rect 312452 159452 312504 159458
rect 312452 159394 312504 159400
rect 311992 159316 312044 159322
rect 311992 159258 312044 159264
rect 311900 157820 311952 157826
rect 311900 157762 311952 157768
rect 311900 157072 311952 157078
rect 311900 157014 311952 157020
rect 311164 153128 311216 153134
rect 311164 153070 311216 153076
rect 311072 153060 311124 153066
rect 311072 153002 311124 153008
rect 310612 150204 310664 150210
rect 310612 150146 310664 150152
rect 311176 150090 311204 153070
rect 311912 151814 311940 157014
rect 312004 156466 312032 159258
rect 312452 156528 312504 156534
rect 312452 156470 312504 156476
rect 311992 156460 312044 156466
rect 311992 156402 312044 156408
rect 311912 151786 312032 151814
rect 312004 150210 312032 151786
rect 312464 150226 312492 156470
rect 313292 154154 313320 163200
rect 314120 158234 314148 163200
rect 314384 158364 314436 158370
rect 314384 158306 314436 158312
rect 314108 158228 314160 158234
rect 314108 158170 314160 158176
rect 313280 154148 313332 154154
rect 313280 154090 313332 154096
rect 313740 152652 313792 152658
rect 313740 152594 313792 152600
rect 313752 150226 313780 152594
rect 314396 150226 314424 158306
rect 314948 152658 314976 163200
rect 315776 158846 315804 163200
rect 315764 158840 315816 158846
rect 315764 158782 315816 158788
rect 316604 154222 316632 163200
rect 317432 158370 317460 163200
rect 318352 160070 318380 163200
rect 318340 160064 318392 160070
rect 318340 160006 318392 160012
rect 319180 159526 319208 163200
rect 317788 159520 317840 159526
rect 317788 159462 317840 159468
rect 319168 159520 319220 159526
rect 319168 159462 319220 159468
rect 317420 158364 317472 158370
rect 317420 158306 317472 158312
rect 316960 157956 317012 157962
rect 316960 157898 317012 157904
rect 315028 154216 315080 154222
rect 315028 154158 315080 154164
rect 316592 154216 316644 154222
rect 316592 154158 316644 154164
rect 314936 152652 314988 152658
rect 314936 152594 314988 152600
rect 315040 150226 315068 154158
rect 315672 153808 315724 153814
rect 315672 153750 315724 153756
rect 315684 150226 315712 153750
rect 316316 152856 316368 152862
rect 316316 152798 316368 152804
rect 316328 150226 316356 152798
rect 316972 150226 317000 157898
rect 317420 157140 317472 157146
rect 317420 157082 317472 157088
rect 317432 151814 317460 157082
rect 317800 156534 317828 159462
rect 318708 158840 318760 158846
rect 318708 158782 318760 158788
rect 317788 156528 317840 156534
rect 317788 156470 317840 156476
rect 317972 155032 318024 155038
rect 317972 154974 318024 154980
rect 317984 151814 318012 154974
rect 318720 153066 318748 158782
rect 319536 158432 319588 158438
rect 319536 158374 319588 158380
rect 318708 153060 318760 153066
rect 318708 153002 318760 153008
rect 318892 152924 318944 152930
rect 318892 152866 318944 152872
rect 317432 151786 317644 151814
rect 317984 151786 318288 151814
rect 317616 150226 317644 151786
rect 318260 150226 318288 151786
rect 318904 150226 318932 152866
rect 319548 150226 319576 158374
rect 320008 154494 320036 163200
rect 320732 159588 320784 159594
rect 320732 159530 320784 159536
rect 319996 154488 320048 154494
rect 319996 154430 320048 154436
rect 320180 154284 320232 154290
rect 320180 154226 320232 154232
rect 320192 150226 320220 154226
rect 320744 151910 320772 159530
rect 320836 158302 320864 163200
rect 320824 158296 320876 158302
rect 320824 158238 320876 158244
rect 321664 157962 321692 163200
rect 322492 163146 322520 163200
rect 322584 163146 322612 163254
rect 322492 163118 322612 163146
rect 322112 158500 322164 158506
rect 322112 158442 322164 158448
rect 321652 157956 321704 157962
rect 321652 157898 321704 157904
rect 320916 154556 320968 154562
rect 320916 154498 320968 154504
rect 320732 151904 320784 151910
rect 320732 151846 320784 151852
rect 320928 150226 320956 154498
rect 321468 153128 321520 153134
rect 321468 153070 321520 153076
rect 311854 150204 311906 150210
rect 311854 150146 311906 150152
rect 311992 150204 312044 150210
rect 312464 150198 312538 150226
rect 311992 150146 312044 150152
rect 307312 150062 307386 150090
rect 307956 150062 308030 150090
rect 308600 150062 308674 150090
rect 309244 150062 309318 150090
rect 309888 150062 309962 150090
rect 310532 150062 310606 150090
rect 311176 150062 311250 150090
rect 307358 149940 307386 150062
rect 308002 149940 308030 150062
rect 308646 149940 308674 150062
rect 309290 149940 309318 150062
rect 309934 149940 309962 150062
rect 310578 149940 310606 150062
rect 311222 149940 311250 150062
rect 311866 149940 311894 150146
rect 312510 149940 312538 150198
rect 313142 150204 313194 150210
rect 313752 150198 313826 150226
rect 314396 150198 314470 150226
rect 315040 150198 315114 150226
rect 315684 150198 315758 150226
rect 316328 150198 316402 150226
rect 316972 150198 317046 150226
rect 317616 150198 317690 150226
rect 318260 150198 318334 150226
rect 318904 150198 318978 150226
rect 319548 150198 319622 150226
rect 320192 150198 320266 150226
rect 313142 150146 313194 150152
rect 313154 149940 313182 150146
rect 313798 149940 313826 150198
rect 314442 149940 314470 150198
rect 315086 149940 315114 150198
rect 315730 149940 315758 150198
rect 316374 149940 316402 150198
rect 317018 149940 317046 150198
rect 317662 149940 317690 150198
rect 318306 149940 318334 150198
rect 318950 149940 318978 150198
rect 319594 149940 319622 150198
rect 320238 149940 320266 150198
rect 320882 150198 320956 150226
rect 321480 150226 321508 153070
rect 322124 150226 322152 158442
rect 322768 152862 322796 163254
rect 323306 163200 323362 164400
rect 324226 163200 324282 164400
rect 325054 163200 325110 164400
rect 325882 163200 325938 164400
rect 326710 163200 326766 164400
rect 326816 163254 327028 163282
rect 322848 154420 322900 154426
rect 322848 154362 322900 154368
rect 322756 152856 322808 152862
rect 322756 152798 322808 152804
rect 322860 150226 322888 154362
rect 323320 154290 323348 163200
rect 323400 156392 323452 156398
rect 323400 156334 323452 156340
rect 323308 154284 323360 154290
rect 323308 154226 323360 154232
rect 321480 150198 321554 150226
rect 322124 150198 322198 150226
rect 320882 149940 320910 150198
rect 321526 149940 321554 150198
rect 322170 149940 322198 150198
rect 322814 150198 322888 150226
rect 323412 150226 323440 156334
rect 324240 155922 324268 163200
rect 325068 159322 325096 163200
rect 325896 159934 325924 163200
rect 326724 163146 326752 163200
rect 326816 163146 326844 163254
rect 326724 163118 326844 163146
rect 325884 159928 325936 159934
rect 325884 159870 325936 159876
rect 325056 159316 325108 159322
rect 325056 159258 325108 159264
rect 324320 159180 324372 159186
rect 324320 159122 324372 159128
rect 324332 157894 324360 159122
rect 324320 157888 324372 157894
rect 324320 157830 324372 157836
rect 324688 157820 324740 157826
rect 324688 157762 324740 157768
rect 324228 155916 324280 155922
rect 324228 155858 324280 155864
rect 324044 152992 324096 152998
rect 324044 152934 324096 152940
rect 324056 150226 324084 152934
rect 324700 150226 324728 157762
rect 327000 154358 327028 163254
rect 327538 163200 327594 164400
rect 328366 163200 328422 164400
rect 329194 163200 329250 164400
rect 330114 163200 330170 164400
rect 330942 163200 330998 164400
rect 331770 163200 331826 164400
rect 332598 163200 332654 164400
rect 333426 163200 333482 164400
rect 334254 163200 334310 164400
rect 335082 163200 335138 164400
rect 336002 163200 336058 164400
rect 336830 163200 336886 164400
rect 337658 163200 337714 164400
rect 337764 163254 338068 163282
rect 327552 158982 327580 163200
rect 328380 161474 328408 163200
rect 328288 161446 328408 161474
rect 329208 161474 329236 163200
rect 329208 161446 329328 161474
rect 327540 158976 327592 158982
rect 327540 158918 327592 158924
rect 327080 158568 327132 158574
rect 327080 158510 327132 158516
rect 325332 154352 325384 154358
rect 325332 154294 325384 154300
rect 326988 154352 327040 154358
rect 326988 154294 327040 154300
rect 325344 150226 325372 154294
rect 325976 153672 326028 153678
rect 325976 153614 326028 153620
rect 325988 150226 326016 153614
rect 326620 151904 326672 151910
rect 326620 151846 326672 151852
rect 326632 150226 326660 151846
rect 327092 151814 327120 158510
rect 327908 155644 327960 155650
rect 327908 155586 327960 155592
rect 327092 151786 327304 151814
rect 327276 150226 327304 151786
rect 327920 150226 327948 155586
rect 328288 152930 328316 161446
rect 328368 158976 328420 158982
rect 328368 158918 328420 158924
rect 328380 155650 328408 158918
rect 328552 158636 328604 158642
rect 328552 158578 328604 158584
rect 328368 155644 328420 155650
rect 328368 155586 328420 155592
rect 328276 152924 328328 152930
rect 328276 152866 328328 152872
rect 328564 150226 328592 158578
rect 329300 152726 329328 161446
rect 330128 158438 330156 163200
rect 330208 159996 330260 160002
rect 330208 159938 330260 159944
rect 330116 158432 330168 158438
rect 330116 158374 330168 158380
rect 329840 157276 329892 157282
rect 329840 157218 329892 157224
rect 329196 152720 329248 152726
rect 329196 152662 329248 152668
rect 329288 152720 329340 152726
rect 329288 152662 329340 152668
rect 329208 150226 329236 152662
rect 329852 150226 329880 157218
rect 330024 155712 330076 155718
rect 330024 155654 330076 155660
rect 330036 151814 330064 155654
rect 330220 155106 330248 159938
rect 330956 157010 330984 163200
rect 331784 159390 331812 163200
rect 332612 160002 332640 163200
rect 332600 159996 332652 160002
rect 332600 159938 332652 159944
rect 332600 159656 332652 159662
rect 332600 159598 332652 159604
rect 331772 159384 331824 159390
rect 331772 159326 331824 159332
rect 331772 158908 331824 158914
rect 331772 158850 331824 158856
rect 331312 158704 331364 158710
rect 331312 158646 331364 158652
rect 330944 157004 330996 157010
rect 330944 156946 330996 156952
rect 331128 155168 331180 155174
rect 331128 155110 331180 155116
rect 330208 155100 330260 155106
rect 330208 155042 330260 155048
rect 330036 151786 330524 151814
rect 330496 150226 330524 151786
rect 331140 150226 331168 155110
rect 323412 150198 323486 150226
rect 324056 150198 324130 150226
rect 324700 150198 324774 150226
rect 325344 150198 325418 150226
rect 325988 150198 326062 150226
rect 326632 150198 326706 150226
rect 327276 150198 327350 150226
rect 327920 150198 327994 150226
rect 328564 150198 328638 150226
rect 329208 150198 329282 150226
rect 329852 150198 329926 150226
rect 330496 150198 330570 150226
rect 331140 150198 331214 150226
rect 331324 150210 331352 158646
rect 331784 150226 331812 158850
rect 332612 151910 332640 159598
rect 333060 155780 333112 155786
rect 333060 155722 333112 155728
rect 332600 151904 332652 151910
rect 332600 151846 332652 151852
rect 333072 150226 333100 155722
rect 333440 153814 333468 163200
rect 334268 155718 334296 163200
rect 334900 156732 334952 156738
rect 334900 156674 334952 156680
rect 334256 155712 334308 155718
rect 334256 155654 334308 155660
rect 333704 153876 333756 153882
rect 333704 153818 333756 153824
rect 333428 153808 333480 153814
rect 333428 153750 333480 153756
rect 333716 150226 333744 153818
rect 334348 152448 334400 152454
rect 334348 152390 334400 152396
rect 334360 150226 334388 152390
rect 334912 150226 334940 156674
rect 335096 154426 335124 163200
rect 336016 158846 336044 163200
rect 336648 160064 336700 160070
rect 336648 160006 336700 160012
rect 336004 158840 336056 158846
rect 336004 158782 336056 158788
rect 336660 155786 336688 160006
rect 336844 157078 336872 163200
rect 337672 163146 337700 163200
rect 337764 163146 337792 163254
rect 337672 163118 337792 163146
rect 337936 158840 337988 158846
rect 337936 158782 337988 158788
rect 336832 157072 336884 157078
rect 336832 157014 336884 157020
rect 336648 155780 336700 155786
rect 336648 155722 336700 155728
rect 335544 155236 335596 155242
rect 335544 155178 335596 155184
rect 335084 154420 335136 154426
rect 335084 154362 335136 154368
rect 335556 150226 335584 155178
rect 337476 154080 337528 154086
rect 337476 154022 337528 154028
rect 336188 153740 336240 153746
rect 336188 153682 336240 153688
rect 336200 150226 336228 153682
rect 336832 151904 336884 151910
rect 336832 151846 336884 151852
rect 336844 150226 336872 151846
rect 337488 150226 337516 154022
rect 337948 152998 337976 158782
rect 338040 154086 338068 163254
rect 338486 163200 338542 164400
rect 339314 163200 339370 164400
rect 340142 163200 340198 164400
rect 340970 163200 341026 164400
rect 341890 163200 341946 164400
rect 342718 163200 342774 164400
rect 343546 163200 343602 164400
rect 344374 163200 344430 164400
rect 345202 163200 345258 164400
rect 346030 163200 346086 164400
rect 346858 163200 346914 164400
rect 347778 163200 347834 164400
rect 348606 163200 348662 164400
rect 349434 163200 349490 164400
rect 350262 163200 350318 164400
rect 351090 163200 351146 164400
rect 351918 163200 351974 164400
rect 352746 163200 352802 164400
rect 353666 163200 353722 164400
rect 354494 163200 354550 164400
rect 355322 163200 355378 164400
rect 356150 163200 356206 164400
rect 356978 163200 357034 164400
rect 357084 163254 357388 163282
rect 338500 158506 338528 163200
rect 338764 159724 338816 159730
rect 338764 159666 338816 159672
rect 338488 158500 338540 158506
rect 338488 158442 338540 158448
rect 338672 157208 338724 157214
rect 338672 157150 338724 157156
rect 338120 155848 338172 155854
rect 338120 155790 338172 155796
rect 338028 154080 338080 154086
rect 338028 154022 338080 154028
rect 337936 152992 337988 152998
rect 337936 152934 337988 152940
rect 338132 150226 338160 155790
rect 338684 151814 338712 157150
rect 338776 154562 338804 159666
rect 339328 159594 339356 163200
rect 339316 159588 339368 159594
rect 339316 159530 339368 159536
rect 340156 158030 340184 163200
rect 340052 158024 340104 158030
rect 340052 157966 340104 157972
rect 340144 158024 340196 158030
rect 340144 157966 340196 157972
rect 339592 155304 339644 155310
rect 339592 155246 339644 155252
rect 338764 154556 338816 154562
rect 338764 154498 338816 154504
rect 338764 154420 338816 154426
rect 338764 154362 338816 154368
rect 338776 153134 338804 154362
rect 339408 153196 339460 153202
rect 339408 153138 339460 153144
rect 338764 153128 338816 153134
rect 338764 153070 338816 153076
rect 338684 151786 338804 151814
rect 338776 150226 338804 151786
rect 339420 150226 339448 153138
rect 322814 149940 322842 150198
rect 323458 149940 323486 150198
rect 324102 149940 324130 150198
rect 324746 149940 324774 150198
rect 325390 149940 325418 150198
rect 326034 149940 326062 150198
rect 326678 149940 326706 150198
rect 327322 149940 327350 150198
rect 327966 149940 327994 150198
rect 328610 149940 328638 150198
rect 329254 149940 329282 150198
rect 329898 149940 329926 150198
rect 330542 149940 330570 150198
rect 331186 149940 331214 150198
rect 331312 150204 331364 150210
rect 331784 150198 331858 150226
rect 331312 150146 331364 150152
rect 331830 149940 331858 150198
rect 332462 150204 332514 150210
rect 333072 150198 333146 150226
rect 333716 150198 333790 150226
rect 334360 150198 334434 150226
rect 334912 150198 334986 150226
rect 335556 150198 335630 150226
rect 336200 150198 336274 150226
rect 336844 150198 336918 150226
rect 337488 150198 337562 150226
rect 338132 150198 338206 150226
rect 338776 150198 338850 150226
rect 339420 150198 339494 150226
rect 339604 150210 339632 155246
rect 340064 150226 340092 157966
rect 340984 154426 341012 163200
rect 341340 157820 341392 157826
rect 341340 157762 341392 157768
rect 340972 154420 341024 154426
rect 340972 154362 341024 154368
rect 341352 150226 341380 157762
rect 341904 156738 341932 163200
rect 342732 160070 342760 163200
rect 342720 160064 342772 160070
rect 342720 160006 342772 160012
rect 342260 158092 342312 158098
rect 342260 158034 342312 158040
rect 341892 156732 341944 156738
rect 341892 156674 341944 156680
rect 341984 154556 342036 154562
rect 341984 154498 342036 154504
rect 341996 150226 342024 154498
rect 342272 151814 342300 158034
rect 343272 155440 343324 155446
rect 343272 155382 343324 155388
rect 342272 151786 342668 151814
rect 342640 150226 342668 151786
rect 343284 150226 343312 155382
rect 343560 155242 343588 163200
rect 343640 159792 343692 159798
rect 343640 159734 343692 159740
rect 343548 155236 343600 155242
rect 343548 155178 343600 155184
rect 343652 151910 343680 159734
rect 343916 155508 343968 155514
rect 343916 155450 343968 155456
rect 343640 151904 343692 151910
rect 343640 151846 343692 151852
rect 343928 150226 343956 155450
rect 344388 155446 344416 163200
rect 345020 157344 345072 157350
rect 345020 157286 345072 157292
rect 344376 155440 344428 155446
rect 344376 155382 344428 155388
rect 344560 152788 344612 152794
rect 344560 152730 344612 152736
rect 344572 150226 344600 152730
rect 345032 151814 345060 157286
rect 345216 155310 345244 163200
rect 346044 159662 346072 163200
rect 346308 159860 346360 159866
rect 346308 159802 346360 159808
rect 346032 159656 346084 159662
rect 346032 159598 346084 159604
rect 346320 155854 346348 159802
rect 346872 157146 346900 163200
rect 347792 157214 347820 163200
rect 347780 157208 347832 157214
rect 347780 157150 347832 157156
rect 346860 157140 346912 157146
rect 346860 157082 346912 157088
rect 348620 156806 348648 163200
rect 347780 156800 347832 156806
rect 347780 156742 347832 156748
rect 348608 156800 348660 156806
rect 348608 156742 348660 156748
rect 346492 156460 346544 156466
rect 346492 156402 346544 156408
rect 346308 155848 346360 155854
rect 346308 155790 346360 155796
rect 345848 155576 345900 155582
rect 345848 155518 345900 155524
rect 345204 155304 345256 155310
rect 345204 155246 345256 155252
rect 345032 151786 345244 151814
rect 345216 150226 345244 151786
rect 345860 150226 345888 155518
rect 346504 150226 346532 156402
rect 347136 151904 347188 151910
rect 347136 151846 347188 151852
rect 347148 150226 347176 151846
rect 347792 150226 347820 156742
rect 349252 156596 349304 156602
rect 349252 156538 349304 156544
rect 348424 155372 348476 155378
rect 348424 155314 348476 155320
rect 348436 150226 348464 155314
rect 349068 154012 349120 154018
rect 349068 153954 349120 153960
rect 349080 150226 349108 153954
rect 332462 150146 332514 150152
rect 332474 149940 332502 150146
rect 333118 149940 333146 150198
rect 333762 149940 333790 150198
rect 334406 149940 334434 150198
rect 334958 149940 334986 150198
rect 335602 149940 335630 150198
rect 336246 149940 336274 150198
rect 336890 149940 336918 150198
rect 337534 149940 337562 150198
rect 338178 149940 338206 150198
rect 338822 149940 338850 150198
rect 339466 149940 339494 150198
rect 339592 150204 339644 150210
rect 340064 150198 340138 150226
rect 339592 150146 339644 150152
rect 340110 149940 340138 150198
rect 340742 150204 340794 150210
rect 341352 150198 341426 150226
rect 341996 150198 342070 150226
rect 342640 150198 342714 150226
rect 343284 150198 343358 150226
rect 343928 150198 344002 150226
rect 344572 150198 344646 150226
rect 345216 150198 345290 150226
rect 345860 150198 345934 150226
rect 346504 150198 346578 150226
rect 347148 150198 347222 150226
rect 347792 150198 347866 150226
rect 348436 150198 348510 150226
rect 349080 150198 349154 150226
rect 349264 150210 349292 156538
rect 349448 152454 349476 163200
rect 350276 158574 350304 163200
rect 350264 158568 350316 158574
rect 350264 158510 350316 158516
rect 351104 158098 351132 163200
rect 351932 158642 351960 163200
rect 352760 159730 352788 163200
rect 352748 159724 352800 159730
rect 352748 159666 352800 159672
rect 352012 159316 352064 159322
rect 352012 159258 352064 159264
rect 351920 158636 351972 158642
rect 351920 158578 351972 158584
rect 351092 158092 351144 158098
rect 351092 158034 351144 158040
rect 350540 157888 350592 157894
rect 350540 157830 350592 157836
rect 349712 152516 349764 152522
rect 349712 152458 349764 152464
rect 349436 152448 349488 152454
rect 349436 152390 349488 152396
rect 349724 150226 349752 152458
rect 340742 150146 340794 150152
rect 340754 149940 340782 150146
rect 341398 149940 341426 150198
rect 342042 149940 342070 150198
rect 342686 149940 342714 150198
rect 343330 149940 343358 150198
rect 343974 149940 344002 150198
rect 344618 149940 344646 150198
rect 345262 149940 345290 150198
rect 345906 149940 345934 150198
rect 346550 149940 346578 150198
rect 347194 149940 347222 150198
rect 347838 149940 347866 150198
rect 348482 149940 348510 150198
rect 349126 149940 349154 150198
rect 349252 150204 349304 150210
rect 349724 150198 349798 150226
rect 350552 150210 350580 157830
rect 352024 157282 352052 159258
rect 353300 158160 353352 158166
rect 353300 158102 353352 158108
rect 352012 157276 352064 157282
rect 352012 157218 352064 157224
rect 351920 156868 351972 156874
rect 351920 156810 351972 156816
rect 351000 156664 351052 156670
rect 351000 156606 351052 156612
rect 351012 150226 351040 156606
rect 349252 150146 349304 150152
rect 349770 149940 349798 150198
rect 350402 150204 350454 150210
rect 350402 150146 350454 150152
rect 350540 150204 350592 150210
rect 351012 150198 351086 150226
rect 351932 150210 351960 156810
rect 352288 155848 352340 155854
rect 352288 155790 352340 155796
rect 352300 150226 352328 155790
rect 353312 151814 353340 158102
rect 353680 155514 353708 163200
rect 354220 156528 354272 156534
rect 354220 156470 354272 156476
rect 353668 155508 353720 155514
rect 353668 155450 353720 155456
rect 353312 151786 353616 151814
rect 353588 150226 353616 151786
rect 354232 150226 354260 156470
rect 354508 155378 354536 163200
rect 355232 159452 355284 159458
rect 355232 159394 355284 159400
rect 354496 155372 354548 155378
rect 354496 155314 354548 155320
rect 355244 153202 355272 159394
rect 355336 154018 355364 163200
rect 356164 157350 356192 163200
rect 356992 163146 357020 163200
rect 357084 163146 357112 163254
rect 356992 163118 357112 163146
rect 356152 157344 356204 157350
rect 356152 157286 356204 157292
rect 356152 156936 356204 156942
rect 356152 156878 356204 156884
rect 355324 154012 355376 154018
rect 355324 153954 355376 153960
rect 355508 153944 355560 153950
rect 355508 153886 355560 153892
rect 355232 153196 355284 153202
rect 355232 153138 355284 153144
rect 354864 152584 354916 152590
rect 354864 152526 354916 152532
rect 354876 150226 354904 152526
rect 355520 150226 355548 153886
rect 356164 150226 356192 156878
rect 356796 155168 356848 155174
rect 356796 155110 356848 155116
rect 356808 150226 356836 155110
rect 357360 154018 357388 163254
rect 357806 163200 357862 164400
rect 358634 163200 358690 164400
rect 359554 163200 359610 164400
rect 360382 163200 360438 164400
rect 361210 163200 361266 164400
rect 362038 163200 362094 164400
rect 362866 163200 362922 164400
rect 363694 163200 363750 164400
rect 364522 163200 364578 164400
rect 365442 163200 365498 164400
rect 366270 163200 366326 164400
rect 367098 163200 367154 164400
rect 367926 163200 367982 164400
rect 368032 163254 368336 163282
rect 357624 158228 357676 158234
rect 357624 158170 357676 158176
rect 357348 154012 357400 154018
rect 357348 153954 357400 153960
rect 357440 153196 357492 153202
rect 357440 153138 357492 153144
rect 357452 150226 357480 153138
rect 350540 150146 350592 150152
rect 350414 149940 350442 150146
rect 351058 149940 351086 150198
rect 351690 150204 351742 150210
rect 351690 150146 351742 150152
rect 351920 150204 351972 150210
rect 352300 150198 352374 150226
rect 351920 150146 351972 150152
rect 351702 149940 351730 150146
rect 352346 149940 352374 150198
rect 352978 150204 353030 150210
rect 353588 150198 353662 150226
rect 354232 150198 354306 150226
rect 354876 150198 354950 150226
rect 355520 150198 355594 150226
rect 356164 150198 356238 150226
rect 356808 150198 356882 150226
rect 357452 150198 357526 150226
rect 357636 150210 357664 158170
rect 357820 156670 357848 163200
rect 358648 158166 358676 163200
rect 359568 159458 359596 163200
rect 359556 159452 359608 159458
rect 359556 159394 359608 159400
rect 360200 158364 360252 158370
rect 360200 158306 360252 158312
rect 358636 158160 358688 158166
rect 358636 158102 358688 158108
rect 359464 157956 359516 157962
rect 359464 157898 359516 157904
rect 358820 157344 358872 157350
rect 358820 157286 358872 157292
rect 357808 156664 357860 156670
rect 357808 156606 357860 156612
rect 358084 154148 358136 154154
rect 358084 154090 358136 154096
rect 358096 150226 358124 154090
rect 358832 152794 358860 157286
rect 358820 152788 358872 152794
rect 358820 152730 358872 152736
rect 359372 152652 359424 152658
rect 359372 152594 359424 152600
rect 359384 150226 359412 152594
rect 359476 151910 359504 157898
rect 360016 153060 360068 153066
rect 360016 153002 360068 153008
rect 359464 151904 359516 151910
rect 359464 151846 359516 151852
rect 360028 150226 360056 153002
rect 352978 150146 353030 150152
rect 352990 149940 353018 150146
rect 353634 149940 353662 150198
rect 354278 149940 354306 150198
rect 354922 149940 354950 150198
rect 355566 149940 355594 150198
rect 356210 149940 356238 150198
rect 356854 149940 356882 150198
rect 357498 149940 357526 150198
rect 357624 150204 357676 150210
rect 358096 150198 358170 150226
rect 357624 150146 357676 150152
rect 358142 149940 358170 150198
rect 358774 150204 358826 150210
rect 359384 150198 359458 150226
rect 360028 150198 360102 150226
rect 360212 150210 360240 158306
rect 360396 154154 360424 163200
rect 361224 158234 361252 163200
rect 361580 159520 361632 159526
rect 361580 159462 361632 159468
rect 361212 158228 361264 158234
rect 361212 158170 361264 158176
rect 360660 154216 360712 154222
rect 360660 154158 360712 154164
rect 360384 154148 360436 154154
rect 360384 154090 360436 154096
rect 360672 150226 360700 154158
rect 358774 150146 358826 150152
rect 358786 149940 358814 150146
rect 359430 149940 359458 150198
rect 360074 149940 360102 150198
rect 360200 150204 360252 150210
rect 360672 150198 360746 150226
rect 361592 150210 361620 159462
rect 362052 158982 362080 163200
rect 362132 159928 362184 159934
rect 362132 159870 362184 159876
rect 362040 158976 362092 158982
rect 362040 158918 362092 158924
rect 362144 155786 362172 159870
rect 362880 158794 362908 163200
rect 362880 158766 363000 158794
rect 361948 155780 362000 155786
rect 361948 155722 362000 155728
rect 362132 155780 362184 155786
rect 362132 155722 362184 155728
rect 361960 150226 361988 155722
rect 362972 152658 363000 158766
rect 363512 158296 363564 158302
rect 363512 158238 363564 158244
rect 363236 154488 363288 154494
rect 363236 154430 363288 154436
rect 362960 152652 363012 152658
rect 362960 152594 363012 152600
rect 363248 150226 363276 154430
rect 363524 151814 363552 158238
rect 363708 156874 363736 163200
rect 363696 156868 363748 156874
rect 363696 156810 363748 156816
rect 364536 155582 364564 163200
rect 364524 155576 364576 155582
rect 364524 155518 364576 155524
rect 365168 152856 365220 152862
rect 365168 152798 365220 152804
rect 364524 151904 364576 151910
rect 364524 151846 364576 151852
rect 363524 151786 363920 151814
rect 363892 150226 363920 151786
rect 364536 150226 364564 151846
rect 365180 150226 365208 152798
rect 365456 152590 365484 163200
rect 366284 159798 366312 163200
rect 366272 159792 366324 159798
rect 366272 159734 366324 159740
rect 366824 158976 366876 158982
rect 366824 158918 366876 158924
rect 365904 157276 365956 157282
rect 365904 157218 365956 157224
rect 365720 154284 365772 154290
rect 365720 154226 365772 154232
rect 365444 152584 365496 152590
rect 365444 152526 365496 152532
rect 365732 150226 365760 154226
rect 360200 150146 360252 150152
rect 360718 149940 360746 150198
rect 361350 150204 361402 150210
rect 361350 150146 361402 150152
rect 361580 150204 361632 150210
rect 361960 150198 362034 150226
rect 361580 150146 361632 150152
rect 361362 149940 361390 150146
rect 362006 149940 362034 150198
rect 362638 150204 362690 150210
rect 363248 150198 363322 150226
rect 363892 150198 363966 150226
rect 364536 150198 364610 150226
rect 365180 150198 365254 150226
rect 365732 150198 365806 150226
rect 365916 150210 365944 157218
rect 366272 155916 366324 155922
rect 366272 155858 366324 155864
rect 366284 151814 366312 155858
rect 366836 154494 366864 158918
rect 367112 158302 367140 163200
rect 367940 163146 367968 163200
rect 368032 163146 368060 163254
rect 367940 163118 368060 163146
rect 367100 158296 367152 158302
rect 367100 158238 367152 158244
rect 367652 155780 367704 155786
rect 367652 155722 367704 155728
rect 366824 154488 366876 154494
rect 366824 154430 366876 154436
rect 366284 151786 366404 151814
rect 366376 150226 366404 151786
rect 367664 150226 367692 155722
rect 368308 154222 368336 163254
rect 368754 163200 368810 164400
rect 369582 163200 369638 164400
rect 370410 163200 370466 164400
rect 371330 163200 371386 164400
rect 372158 163200 372214 164400
rect 372986 163200 373042 164400
rect 373814 163200 373870 164400
rect 374642 163200 374698 164400
rect 375470 163200 375526 164400
rect 376298 163200 376354 164400
rect 376404 163254 376708 163282
rect 368480 159996 368532 160002
rect 368480 159938 368532 159944
rect 368388 154352 368440 154358
rect 368388 154294 368440 154300
rect 368296 154216 368348 154222
rect 368296 154158 368348 154164
rect 368400 150226 368428 154294
rect 368492 153202 368520 159938
rect 368768 159526 368796 163200
rect 368756 159520 368808 159526
rect 368756 159462 368808 159468
rect 369596 155650 369624 163200
rect 370424 155786 370452 163200
rect 370872 158432 370924 158438
rect 370872 158374 370924 158380
rect 370412 155780 370464 155786
rect 370412 155722 370464 155728
rect 368940 155644 368992 155650
rect 368940 155586 368992 155592
rect 369584 155644 369636 155650
rect 369584 155586 369636 155592
rect 368480 153196 368532 153202
rect 368480 153138 368532 153144
rect 362638 150146 362690 150152
rect 362650 149940 362678 150146
rect 363294 149940 363322 150198
rect 363938 149940 363966 150198
rect 364582 149940 364610 150198
rect 365226 149940 365254 150198
rect 365778 149940 365806 150198
rect 365904 150204 365956 150210
rect 366376 150198 366450 150226
rect 365904 150146 365956 150152
rect 366422 149940 366450 150198
rect 367054 150204 367106 150210
rect 367664 150198 367738 150226
rect 367054 150146 367106 150152
rect 367066 149940 367094 150146
rect 367710 149940 367738 150198
rect 368354 150198 368428 150226
rect 368952 150226 368980 155586
rect 369584 152924 369636 152930
rect 369584 152866 369636 152872
rect 369596 150226 369624 152866
rect 370228 152720 370280 152726
rect 370228 152662 370280 152668
rect 370240 150226 370268 152662
rect 370884 150226 370912 158374
rect 371240 157004 371292 157010
rect 371240 156946 371292 156952
rect 371252 151814 371280 156946
rect 371344 154290 371372 163200
rect 372068 159384 372120 159390
rect 372068 159326 372120 159332
rect 371332 154284 371384 154290
rect 371332 154226 371384 154232
rect 372080 151814 372108 159326
rect 372172 158982 372200 163200
rect 372620 160064 372672 160070
rect 372620 160006 372672 160012
rect 372160 158976 372212 158982
rect 372160 158918 372212 158924
rect 372632 152930 372660 160006
rect 373000 159390 373028 163200
rect 372988 159384 373040 159390
rect 372988 159326 373040 159332
rect 373828 157010 373856 163200
rect 374276 158976 374328 158982
rect 374276 158918 374328 158924
rect 373816 157004 373868 157010
rect 373816 156946 373868 156952
rect 374092 155712 374144 155718
rect 374092 155654 374144 155660
rect 373448 153876 373500 153882
rect 373448 153818 373500 153824
rect 372804 153196 372856 153202
rect 372804 153138 372856 153144
rect 372620 152924 372672 152930
rect 372620 152866 372672 152872
rect 371252 151786 371556 151814
rect 372080 151786 372200 151814
rect 371528 150226 371556 151786
rect 372172 150226 372200 151786
rect 372816 150226 372844 153138
rect 373460 150226 373488 153818
rect 374104 150226 374132 155654
rect 374288 152862 374316 158918
rect 374656 156942 374684 163200
rect 375484 159866 375512 163200
rect 376312 163146 376340 163200
rect 376404 163146 376432 163254
rect 376312 163118 376432 163146
rect 375472 159860 375524 159866
rect 375472 159802 375524 159808
rect 376024 157072 376076 157078
rect 376024 157014 376076 157020
rect 374644 156936 374696 156942
rect 374644 156878 374696 156884
rect 374736 153128 374788 153134
rect 374736 153070 374788 153076
rect 374276 152856 374328 152862
rect 374276 152798 374328 152804
rect 374748 150226 374776 153070
rect 375380 152992 375432 152998
rect 375380 152934 375432 152940
rect 375392 150226 375420 152934
rect 376036 150226 376064 157014
rect 376576 154080 376628 154086
rect 376576 154022 376628 154028
rect 376588 151814 376616 154022
rect 376680 152726 376708 163254
rect 377218 163200 377274 164400
rect 378046 163200 378102 164400
rect 378874 163200 378930 164400
rect 379702 163200 379758 164400
rect 380530 163200 380586 164400
rect 380636 163254 380848 163282
rect 377232 158506 377260 163200
rect 377956 159588 378008 159594
rect 377956 159530 378008 159536
rect 376852 158500 376904 158506
rect 376852 158442 376904 158448
rect 377220 158500 377272 158506
rect 377220 158442 377272 158448
rect 376668 152720 376720 152726
rect 376668 152662 376720 152668
rect 376864 151814 376892 158442
rect 376588 151786 376708 151814
rect 376864 151786 377352 151814
rect 376680 150226 376708 151786
rect 377324 150226 377352 151786
rect 377968 150226 377996 159530
rect 378060 158370 378088 163200
rect 378140 159656 378192 159662
rect 378140 159598 378192 159604
rect 378048 158364 378100 158370
rect 378048 158306 378100 158312
rect 378152 155922 378180 159598
rect 378888 158778 378916 163200
rect 379716 159594 379744 163200
rect 380544 163146 380572 163200
rect 380636 163146 380664 163254
rect 380544 163118 380664 163146
rect 379704 159588 379756 159594
rect 379704 159530 379756 159536
rect 378876 158772 378928 158778
rect 378876 158714 378928 158720
rect 378600 158024 378652 158030
rect 378600 157966 378652 157972
rect 378140 155916 378192 155922
rect 378140 155858 378192 155864
rect 378612 150226 378640 157966
rect 379888 156732 379940 156738
rect 379888 156674 379940 156680
rect 379244 154420 379296 154426
rect 379244 154362 379296 154368
rect 379256 150226 379284 154362
rect 379900 150226 379928 156674
rect 380820 153882 380848 163254
rect 381358 163200 381414 164400
rect 382186 163200 382242 164400
rect 383106 163200 383162 164400
rect 383934 163200 383990 164400
rect 384762 163200 384818 164400
rect 385590 163200 385646 164400
rect 386418 163200 386474 164400
rect 387246 163200 387302 164400
rect 388074 163200 388130 164400
rect 388994 163200 389050 164400
rect 389822 163200 389878 164400
rect 390650 163200 390706 164400
rect 391478 163200 391534 164400
rect 391584 163254 391888 163282
rect 380992 158772 381044 158778
rect 380992 158714 381044 158720
rect 380900 155440 380952 155446
rect 380900 155382 380952 155388
rect 380808 153876 380860 153882
rect 380808 153818 380860 153824
rect 380532 152924 380584 152930
rect 380532 152866 380584 152872
rect 380544 150226 380572 152866
rect 368952 150198 369026 150226
rect 369596 150198 369670 150226
rect 370240 150198 370314 150226
rect 370884 150198 370958 150226
rect 371528 150198 371602 150226
rect 372172 150198 372246 150226
rect 372816 150198 372890 150226
rect 373460 150198 373534 150226
rect 374104 150198 374178 150226
rect 374748 150198 374822 150226
rect 375392 150198 375466 150226
rect 376036 150198 376110 150226
rect 376680 150198 376754 150226
rect 377324 150198 377398 150226
rect 377968 150198 378042 150226
rect 378612 150198 378686 150226
rect 379256 150198 379330 150226
rect 379900 150198 379974 150226
rect 380544 150198 380618 150226
rect 380912 150210 380940 155382
rect 381004 152930 381032 158714
rect 381372 155242 381400 163200
rect 382200 159662 382228 163200
rect 382188 159656 382240 159662
rect 382188 159598 382240 159604
rect 383120 157078 383148 163200
rect 383752 157140 383804 157146
rect 383752 157082 383804 157088
rect 383108 157072 383160 157078
rect 383108 157014 383160 157020
rect 382280 155916 382332 155922
rect 382280 155858 382332 155864
rect 381176 155236 381228 155242
rect 381176 155178 381228 155184
rect 381360 155236 381412 155242
rect 381360 155178 381412 155184
rect 380992 152924 381044 152930
rect 380992 152866 381044 152872
rect 381188 150226 381216 155178
rect 368354 149940 368382 150198
rect 368998 149940 369026 150198
rect 369642 149940 369670 150198
rect 370286 149940 370314 150198
rect 370930 149940 370958 150198
rect 371574 149940 371602 150198
rect 372218 149940 372246 150198
rect 372862 149940 372890 150198
rect 373506 149940 373534 150198
rect 374150 149940 374178 150198
rect 374794 149940 374822 150198
rect 375438 149940 375466 150198
rect 376082 149940 376110 150198
rect 376726 149940 376754 150198
rect 377370 149940 377398 150198
rect 378014 149940 378042 150198
rect 378658 149940 378686 150198
rect 379302 149940 379330 150198
rect 379946 149940 379974 150198
rect 380590 149940 380618 150198
rect 380900 150204 380952 150210
rect 381188 150198 381262 150226
rect 382292 150210 382320 155858
rect 382464 155304 382516 155310
rect 382464 155246 382516 155252
rect 382476 150226 382504 155246
rect 383764 150226 383792 157082
rect 383948 155310 383976 163200
rect 384396 157208 384448 157214
rect 384396 157150 384448 157156
rect 383936 155304 383988 155310
rect 383936 155246 383988 155252
rect 384408 150226 384436 157150
rect 384776 156738 384804 163200
rect 385604 158778 385632 163200
rect 386432 159934 386460 163200
rect 386420 159928 386472 159934
rect 386420 159870 386472 159876
rect 385960 159724 386012 159730
rect 385960 159666 386012 159672
rect 385592 158772 385644 158778
rect 385592 158714 385644 158720
rect 385224 158568 385276 158574
rect 385224 158510 385276 158516
rect 385040 156800 385092 156806
rect 385040 156742 385092 156748
rect 384764 156732 384816 156738
rect 384764 156674 384816 156680
rect 385052 150226 385080 156742
rect 380900 150146 380952 150152
rect 381234 149940 381262 150198
rect 381866 150204 381918 150210
rect 381866 150146 381918 150152
rect 382280 150204 382332 150210
rect 382476 150198 382550 150226
rect 382280 150146 382332 150152
rect 381878 149940 381906 150146
rect 382522 149940 382550 150198
rect 383154 150204 383206 150210
rect 383764 150198 383838 150226
rect 384408 150198 384482 150226
rect 385052 150198 385126 150226
rect 385236 150210 385264 158510
rect 385972 153202 386000 159666
rect 386512 158636 386564 158642
rect 386512 158578 386564 158584
rect 385960 153196 386012 153202
rect 385960 153138 386012 153144
rect 385592 152516 385644 152522
rect 385592 152458 385644 152464
rect 385604 151814 385632 152458
rect 385604 151786 385724 151814
rect 385696 150226 385724 151786
rect 383154 150146 383206 150152
rect 383166 149940 383194 150146
rect 383810 149940 383838 150198
rect 384454 149940 384482 150198
rect 385098 149940 385126 150198
rect 385224 150204 385276 150210
rect 385696 150198 385770 150226
rect 386524 150210 386552 158578
rect 386972 158092 387024 158098
rect 386972 158034 387024 158040
rect 386984 150226 387012 158034
rect 387260 156806 387288 163200
rect 388088 158030 388116 163200
rect 389008 159730 389036 163200
rect 388996 159724 389048 159730
rect 388996 159666 389048 159672
rect 389836 158778 389864 163200
rect 389088 158772 389140 158778
rect 389088 158714 389140 158720
rect 389824 158772 389876 158778
rect 389824 158714 389876 158720
rect 388076 158024 388128 158030
rect 388076 157966 388128 157972
rect 387248 156800 387300 156806
rect 387248 156742 387300 156748
rect 388352 155508 388404 155514
rect 388352 155450 388404 155456
rect 388260 153196 388312 153202
rect 388260 153138 388312 153144
rect 388272 150226 388300 153138
rect 388364 151814 388392 155450
rect 389100 152998 389128 158714
rect 389548 155372 389600 155378
rect 389548 155314 389600 155320
rect 389088 152992 389140 152998
rect 389088 152934 389140 152940
rect 388364 151786 388944 151814
rect 388916 150226 388944 151786
rect 389560 150226 389588 155314
rect 390664 153950 390692 163200
rect 391492 163146 391520 163200
rect 391584 163146 391612 163254
rect 391492 163118 391612 163146
rect 391572 158772 391624 158778
rect 391572 158714 391624 158720
rect 391480 154012 391532 154018
rect 391480 153954 391532 153960
rect 390192 153944 390244 153950
rect 390192 153886 390244 153892
rect 390652 153944 390704 153950
rect 390652 153886 390704 153892
rect 390204 150226 390232 153886
rect 390836 152788 390888 152794
rect 390836 152730 390888 152736
rect 390848 150226 390876 152730
rect 391492 150226 391520 153954
rect 391584 152794 391612 158714
rect 391860 154018 391888 163254
rect 392306 163200 392362 164400
rect 393134 163200 393190 164400
rect 393962 163200 394018 164400
rect 394882 163200 394938 164400
rect 395710 163200 395766 164400
rect 396538 163200 396594 164400
rect 397366 163200 397422 164400
rect 398194 163200 398250 164400
rect 399022 163200 399078 164400
rect 399850 163200 399906 164400
rect 400770 163200 400826 164400
rect 401598 163200 401654 164400
rect 402426 163200 402482 164400
rect 403254 163200 403310 164400
rect 404082 163200 404138 164400
rect 404910 163200 404966 164400
rect 405738 163200 405794 164400
rect 406658 163200 406714 164400
rect 407486 163200 407542 164400
rect 408314 163200 408370 164400
rect 409142 163200 409198 164400
rect 409970 163200 410026 164400
rect 410798 163200 410854 164400
rect 411626 163200 411682 164400
rect 412546 163200 412602 164400
rect 413374 163200 413430 164400
rect 414202 163200 414258 164400
rect 415030 163200 415086 164400
rect 415858 163200 415914 164400
rect 416686 163200 416742 164400
rect 417514 163200 417570 164400
rect 418434 163200 418490 164400
rect 419262 163200 419318 164400
rect 420090 163200 420146 164400
rect 420918 163200 420974 164400
rect 421746 163200 421802 164400
rect 422574 163200 422630 164400
rect 423402 163200 423458 164400
rect 424322 163200 424378 164400
rect 425150 163200 425206 164400
rect 425978 163200 426034 164400
rect 426806 163200 426862 164400
rect 427634 163200 427690 164400
rect 428462 163200 428518 164400
rect 429290 163200 429346 164400
rect 430210 163200 430266 164400
rect 431038 163200 431094 164400
rect 431866 163200 431922 164400
rect 432694 163200 432750 164400
rect 433522 163200 433578 164400
rect 434350 163200 434406 164400
rect 435178 163200 435234 164400
rect 436098 163200 436154 164400
rect 436926 163200 436982 164400
rect 437032 163254 437428 163282
rect 391940 158160 391992 158166
rect 391940 158102 391992 158108
rect 391848 154012 391900 154018
rect 391848 153954 391900 153960
rect 391572 152788 391624 152794
rect 391572 152730 391624 152736
rect 385224 150146 385276 150152
rect 385742 149940 385770 150198
rect 386374 150204 386426 150210
rect 386374 150146 386426 150152
rect 386512 150204 386564 150210
rect 386984 150198 387058 150226
rect 386512 150146 386564 150152
rect 386386 149940 386414 150146
rect 387030 149940 387058 150198
rect 387662 150204 387714 150210
rect 388272 150198 388346 150226
rect 388916 150198 388990 150226
rect 389560 150198 389634 150226
rect 390204 150198 390278 150226
rect 390848 150198 390922 150226
rect 391492 150198 391566 150226
rect 391952 150210 391980 158102
rect 392124 156664 392176 156670
rect 392124 156606 392176 156612
rect 392136 150226 392164 156606
rect 392320 152522 392348 163200
rect 393148 160002 393176 163200
rect 393136 159996 393188 160002
rect 393136 159938 393188 159944
rect 393412 159452 393464 159458
rect 393412 159394 393464 159400
rect 392308 152516 392360 152522
rect 392308 152458 392360 152464
rect 393424 150226 393452 159394
rect 393976 158098 394004 163200
rect 394700 158228 394752 158234
rect 394700 158170 394752 158176
rect 393964 158092 394016 158098
rect 393964 158034 394016 158040
rect 394056 154148 394108 154154
rect 394056 154090 394108 154096
rect 394068 150226 394096 154090
rect 394712 150226 394740 158170
rect 394896 155446 394924 163200
rect 395724 159458 395752 163200
rect 396552 161474 396580 163200
rect 396552 161446 396672 161474
rect 395712 159452 395764 159458
rect 395712 159394 395764 159400
rect 396540 156868 396592 156874
rect 396540 156810 396592 156816
rect 396172 155576 396224 155582
rect 396172 155518 396224 155524
rect 394884 155440 394936 155446
rect 394884 155382 394936 155388
rect 395344 154488 395396 154494
rect 395344 154430 395396 154436
rect 395356 150226 395384 154430
rect 395988 152652 396040 152658
rect 395988 152594 396040 152600
rect 396000 150226 396028 152594
rect 387662 150146 387714 150152
rect 387674 149940 387702 150146
rect 388318 149940 388346 150198
rect 388962 149940 388990 150198
rect 389606 149940 389634 150198
rect 390250 149940 390278 150198
rect 390894 149940 390922 150198
rect 391538 149940 391566 150198
rect 391940 150204 391992 150210
rect 392136 150198 392210 150226
rect 391940 150146 391992 150152
rect 392182 149940 392210 150198
rect 392814 150204 392866 150210
rect 393424 150198 393498 150226
rect 394068 150198 394142 150226
rect 394712 150198 394786 150226
rect 395356 150198 395430 150226
rect 396000 150198 396074 150226
rect 396184 150210 396212 155518
rect 396552 150226 396580 156810
rect 396644 152658 396672 161446
rect 397380 155378 397408 163200
rect 397368 155372 397420 155378
rect 397368 155314 397420 155320
rect 398208 154086 398236 163200
rect 398472 159792 398524 159798
rect 398472 159734 398524 159740
rect 398196 154080 398248 154086
rect 398196 154022 398248 154028
rect 396632 152652 396684 152658
rect 396632 152594 396684 152600
rect 397828 152584 397880 152590
rect 397828 152526 397880 152532
rect 397840 150226 397868 152526
rect 398484 150226 398512 159734
rect 399036 153066 399064 163200
rect 399864 159798 399892 163200
rect 399852 159792 399904 159798
rect 399852 159734 399904 159740
rect 400404 159520 400456 159526
rect 400404 159462 400456 159468
rect 399116 158296 399168 158302
rect 399116 158238 399168 158244
rect 399024 153060 399076 153066
rect 399024 153002 399076 153008
rect 399128 150226 399156 158238
rect 400220 155644 400272 155650
rect 400220 155586 400272 155592
rect 399760 154216 399812 154222
rect 399760 154158 399812 154164
rect 399772 150226 399800 154158
rect 392814 150146 392866 150152
rect 392826 149940 392854 150146
rect 393470 149940 393498 150198
rect 394114 149940 394142 150198
rect 394758 149940 394786 150198
rect 395402 149940 395430 150198
rect 396046 149940 396074 150198
rect 396172 150204 396224 150210
rect 396552 150198 396626 150226
rect 396172 150146 396224 150152
rect 396598 149940 396626 150198
rect 397230 150204 397282 150210
rect 397840 150198 397914 150226
rect 398484 150198 398558 150226
rect 399128 150198 399202 150226
rect 399772 150198 399846 150226
rect 400232 150210 400260 155586
rect 400416 150226 400444 159462
rect 400784 156670 400812 163200
rect 401612 156874 401640 163200
rect 402440 159526 402468 163200
rect 402428 159520 402480 159526
rect 402428 159462 402480 159468
rect 403164 159384 403216 159390
rect 403164 159326 403216 159332
rect 401600 156868 401652 156874
rect 401600 156810 401652 156816
rect 400772 156664 400824 156670
rect 400772 156606 400824 156612
rect 401692 155780 401744 155786
rect 401692 155722 401744 155728
rect 401704 150226 401732 155722
rect 402336 154284 402388 154290
rect 402336 154226 402388 154232
rect 402348 150226 402376 154226
rect 402980 152856 403032 152862
rect 402980 152798 403032 152804
rect 402992 150226 403020 152798
rect 403176 151814 403204 159326
rect 403268 152590 403296 163200
rect 404096 158234 404124 163200
rect 404084 158228 404136 158234
rect 404084 158170 404136 158176
rect 404924 158166 404952 163200
rect 405556 159860 405608 159866
rect 405556 159802 405608 159808
rect 404912 158160 404964 158166
rect 404912 158102 404964 158108
rect 404084 157004 404136 157010
rect 404084 156946 404136 156952
rect 403256 152584 403308 152590
rect 403256 152526 403308 152532
rect 404096 151814 404124 156946
rect 404452 156936 404504 156942
rect 404452 156878 404504 156884
rect 404464 151814 404492 156878
rect 403176 151786 403664 151814
rect 404096 151786 404308 151814
rect 404464 151786 404952 151814
rect 403636 150226 403664 151786
rect 404280 150226 404308 151786
rect 404924 150226 404952 151786
rect 405568 150226 405596 159802
rect 405752 158982 405780 163200
rect 406672 159866 406700 163200
rect 406660 159860 406712 159866
rect 406660 159802 406712 159808
rect 405740 158976 405792 158982
rect 405740 158918 405792 158924
rect 407028 158976 407080 158982
rect 407028 158918 407080 158924
rect 406844 158500 406896 158506
rect 406844 158442 406896 158448
rect 406200 152720 406252 152726
rect 406200 152662 406252 152668
rect 406212 150226 406240 152662
rect 406856 150226 406884 158442
rect 407040 152726 407068 158918
rect 407396 158364 407448 158370
rect 407396 158306 407448 158312
rect 407028 152720 407080 152726
rect 407028 152662 407080 152668
rect 407408 151814 407436 158306
rect 407500 154154 407528 163200
rect 408328 155514 408356 163200
rect 409156 160070 409184 163200
rect 409144 160064 409196 160070
rect 409144 160006 409196 160012
rect 408500 159656 408552 159662
rect 408500 159598 408552 159604
rect 408316 155508 408368 155514
rect 408316 155450 408368 155456
rect 407488 154148 407540 154154
rect 407488 154090 407540 154096
rect 408512 153202 408540 159598
rect 408776 159588 408828 159594
rect 408776 159530 408828 159536
rect 408500 153196 408552 153202
rect 408500 153138 408552 153144
rect 408132 152924 408184 152930
rect 408132 152866 408184 152872
rect 407408 151786 407528 151814
rect 407500 150226 407528 151786
rect 408144 150226 408172 152866
rect 408788 150226 408816 159530
rect 409420 153876 409472 153882
rect 409420 153818 409472 153824
rect 409432 150226 409460 153818
rect 409984 152930 410012 163200
rect 410812 155242 410840 163200
rect 411352 157072 411404 157078
rect 411352 157014 411404 157020
rect 410064 155236 410116 155242
rect 410064 155178 410116 155184
rect 410800 155236 410852 155242
rect 410800 155178 410852 155184
rect 409972 152924 410024 152930
rect 409972 152866 410024 152872
rect 410076 150226 410104 155178
rect 410708 153196 410760 153202
rect 410708 153138 410760 153144
rect 410720 150226 410748 153138
rect 411364 150226 411392 157014
rect 411640 156942 411668 163200
rect 411628 156936 411680 156942
rect 411628 156878 411680 156884
rect 411996 155304 412048 155310
rect 411996 155246 412048 155252
rect 412008 150226 412036 155246
rect 412560 152862 412588 163200
rect 412824 159928 412876 159934
rect 412824 159870 412876 159876
rect 412640 156732 412692 156738
rect 412640 156674 412692 156680
rect 412548 152856 412600 152862
rect 412548 152798 412600 152804
rect 412652 150226 412680 156674
rect 397230 150146 397282 150152
rect 397242 149940 397270 150146
rect 397886 149940 397914 150198
rect 398530 149940 398558 150198
rect 399174 149940 399202 150198
rect 399818 149940 399846 150198
rect 400220 150204 400272 150210
rect 400416 150198 400490 150226
rect 400220 150146 400272 150152
rect 400462 149940 400490 150198
rect 401094 150204 401146 150210
rect 401704 150198 401778 150226
rect 402348 150198 402422 150226
rect 402992 150198 403066 150226
rect 403636 150198 403710 150226
rect 404280 150198 404354 150226
rect 404924 150198 404998 150226
rect 405568 150198 405642 150226
rect 406212 150198 406286 150226
rect 406856 150198 406930 150226
rect 407500 150198 407574 150226
rect 408144 150198 408218 150226
rect 408788 150198 408862 150226
rect 409432 150198 409506 150226
rect 410076 150198 410150 150226
rect 410720 150198 410794 150226
rect 411364 150198 411438 150226
rect 412008 150198 412082 150226
rect 412652 150198 412726 150226
rect 412836 150210 412864 159870
rect 413388 159662 413416 163200
rect 413376 159656 413428 159662
rect 413376 159598 413428 159604
rect 414216 156806 414244 163200
rect 414296 159724 414348 159730
rect 414296 159666 414348 159672
rect 414112 156800 414164 156806
rect 414112 156742 414164 156748
rect 414204 156800 414256 156806
rect 414204 156742 414256 156748
rect 413284 152992 413336 152998
rect 413284 152934 413336 152940
rect 413296 150226 413324 152934
rect 414124 151814 414152 156742
rect 414308 152454 414336 159666
rect 415044 158030 415072 163200
rect 414572 158024 414624 158030
rect 414572 157966 414624 157972
rect 415032 158024 415084 158030
rect 415032 157966 415084 157972
rect 414296 152448 414348 152454
rect 414296 152390 414348 152396
rect 414584 151814 414612 157966
rect 415872 152998 415900 163200
rect 415860 152992 415912 152998
rect 415860 152934 415912 152940
rect 416700 152794 416728 163200
rect 417148 153944 417200 153950
rect 417148 153886 417200 153892
rect 416504 152788 416556 152794
rect 416504 152730 416556 152736
rect 416688 152788 416740 152794
rect 416688 152730 416740 152736
rect 415860 152448 415912 152454
rect 415860 152390 415912 152396
rect 414124 151786 414520 151814
rect 414584 151786 415256 151814
rect 414492 150226 414520 151786
rect 415228 150226 415256 151786
rect 415872 150226 415900 152390
rect 416516 150226 416544 152730
rect 417160 150226 417188 153886
rect 417528 153882 417556 163200
rect 417792 154012 417844 154018
rect 417792 153954 417844 153960
rect 417516 153876 417568 153882
rect 417516 153818 417568 153824
rect 417804 150226 417832 153954
rect 418448 153950 418476 163200
rect 419080 159996 419132 160002
rect 419080 159938 419132 159944
rect 418436 153944 418488 153950
rect 418436 153886 418488 153892
rect 418436 152516 418488 152522
rect 418436 152458 418488 152464
rect 418448 150226 418476 152458
rect 419092 150226 419120 159938
rect 419276 156738 419304 163200
rect 420104 159730 420132 163200
rect 420092 159724 420144 159730
rect 420092 159666 420144 159672
rect 420932 158098 420960 163200
rect 421104 159452 421156 159458
rect 421104 159394 421156 159400
rect 419540 158092 419592 158098
rect 419540 158034 419592 158040
rect 420920 158092 420972 158098
rect 420920 158034 420972 158040
rect 419264 156732 419316 156738
rect 419264 156674 419316 156680
rect 419552 151814 419580 158034
rect 420368 155440 420420 155446
rect 420368 155382 420420 155388
rect 419552 151786 419764 151814
rect 419736 150226 419764 151786
rect 420380 150226 420408 155382
rect 421116 150226 421144 159394
rect 421760 155310 421788 163200
rect 422300 155372 422352 155378
rect 422300 155314 422352 155320
rect 421748 155304 421800 155310
rect 421748 155246 421800 155252
rect 421656 152652 421708 152658
rect 421656 152594 421708 152600
rect 401094 150146 401146 150152
rect 401106 149940 401134 150146
rect 401750 149940 401778 150198
rect 402394 149940 402422 150198
rect 403038 149940 403066 150198
rect 403682 149940 403710 150198
rect 404326 149940 404354 150198
rect 404970 149940 404998 150198
rect 405614 149940 405642 150198
rect 406258 149940 406286 150198
rect 406902 149940 406930 150198
rect 407546 149940 407574 150198
rect 408190 149940 408218 150198
rect 408834 149940 408862 150198
rect 409478 149940 409506 150198
rect 410122 149940 410150 150198
rect 410766 149940 410794 150198
rect 411410 149940 411438 150198
rect 412054 149940 412082 150198
rect 412698 149940 412726 150198
rect 412824 150204 412876 150210
rect 413296 150198 413370 150226
rect 412824 150146 412876 150152
rect 413342 149940 413370 150198
rect 413974 150204 414026 150210
rect 414492 150198 414658 150226
rect 415228 150198 415302 150226
rect 415872 150198 415946 150226
rect 416516 150198 416590 150226
rect 417160 150198 417234 150226
rect 417804 150198 417878 150226
rect 418448 150198 418522 150226
rect 419092 150198 419166 150226
rect 419736 150198 419810 150226
rect 420380 150198 420454 150226
rect 413974 150146 414026 150152
rect 413986 149940 414014 150146
rect 414630 149940 414658 150198
rect 415274 149940 415302 150198
rect 415918 149940 415946 150198
rect 416562 149940 416590 150198
rect 417206 149940 417234 150198
rect 417850 149940 417878 150198
rect 418494 149940 418522 150198
rect 419138 149940 419166 150198
rect 419782 149940 419810 150198
rect 420426 149940 420454 150198
rect 421070 150198 421144 150226
rect 421668 150226 421696 152594
rect 422312 150226 422340 155314
rect 422588 154222 422616 163200
rect 423416 157010 423444 163200
rect 424232 159792 424284 159798
rect 424232 159734 424284 159740
rect 423404 157004 423456 157010
rect 423404 156946 423456 156952
rect 423772 156664 423824 156670
rect 423772 156606 423824 156612
rect 422576 154216 422628 154222
rect 422576 154158 422628 154164
rect 422944 154080 422996 154086
rect 422944 154022 422996 154028
rect 422956 150226 422984 154022
rect 423588 153060 423640 153066
rect 423588 153002 423640 153008
rect 423600 150226 423628 153002
rect 421668 150198 421742 150226
rect 422312 150198 422386 150226
rect 422956 150198 423030 150226
rect 423600 150198 423674 150226
rect 423784 150210 423812 156606
rect 424244 150226 424272 159734
rect 424336 155378 424364 163200
rect 425164 161474 425192 163200
rect 425164 161446 425284 161474
rect 425152 156868 425204 156874
rect 425152 156810 425204 156816
rect 424324 155372 424376 155378
rect 424324 155314 424376 155320
rect 425164 151814 425192 156810
rect 425256 154018 425284 161446
rect 425992 160002 426020 163200
rect 425980 159996 426032 160002
rect 425980 159938 426032 159944
rect 426440 159996 426492 160002
rect 426440 159938 426492 159944
rect 426164 159520 426216 159526
rect 426164 159462 426216 159468
rect 425244 154012 425296 154018
rect 425244 153954 425296 153960
rect 425164 151786 425560 151814
rect 425532 150226 425560 151786
rect 426176 150226 426204 159462
rect 426452 158234 426480 159938
rect 426820 159390 426848 163200
rect 426808 159384 426860 159390
rect 426808 159326 426860 159332
rect 427360 158364 427412 158370
rect 427360 158306 427412 158312
rect 426440 158228 426492 158234
rect 426440 158170 426492 158176
rect 426808 152584 426860 152590
rect 426808 152526 426860 152532
rect 426820 150226 426848 152526
rect 427372 150226 427400 158306
rect 427648 156670 427676 163200
rect 428476 158166 428504 163200
rect 428004 158160 428056 158166
rect 428004 158102 428056 158108
rect 428464 158160 428516 158166
rect 428464 158102 428516 158108
rect 427636 156664 427688 156670
rect 427636 156606 427688 156612
rect 428016 150226 428044 158102
rect 429304 155446 429332 163200
rect 430224 160002 430252 163200
rect 430212 159996 430264 160002
rect 430212 159938 430264 159944
rect 429384 159860 429436 159866
rect 429384 159802 429436 159808
rect 429292 155440 429344 155446
rect 429292 155382 429344 155388
rect 428648 152720 428700 152726
rect 428648 152662 428700 152668
rect 428660 150226 428688 152662
rect 429396 150226 429424 159802
rect 430580 155508 430632 155514
rect 430580 155450 430632 155456
rect 429936 154148 429988 154154
rect 429936 154090 429988 154096
rect 421070 149940 421098 150198
rect 421714 149940 421742 150198
rect 422358 149940 422386 150198
rect 423002 149940 423030 150198
rect 423646 149940 423674 150198
rect 423772 150204 423824 150210
rect 424244 150198 424318 150226
rect 423772 150146 423824 150152
rect 424290 149940 424318 150198
rect 424922 150204 424974 150210
rect 425532 150198 425606 150226
rect 426176 150198 426250 150226
rect 426820 150198 426894 150226
rect 427372 150198 427446 150226
rect 428016 150198 428090 150226
rect 428660 150198 428734 150226
rect 424922 150146 424974 150152
rect 424934 149940 424962 150146
rect 425578 149940 425606 150198
rect 426222 149940 426250 150198
rect 426866 149940 426894 150198
rect 427418 149940 427446 150198
rect 428062 149940 428090 150198
rect 428706 149940 428734 150198
rect 429350 150198 429424 150226
rect 429948 150226 429976 154090
rect 430592 150226 430620 155450
rect 431052 154154 431080 163200
rect 431224 160064 431276 160070
rect 431224 160006 431276 160012
rect 431040 154148 431092 154154
rect 431040 154090 431092 154096
rect 431236 150226 431264 160006
rect 431880 159594 431908 163200
rect 431868 159588 431920 159594
rect 431868 159530 431920 159536
rect 432708 159458 432736 163200
rect 433064 159996 433116 160002
rect 433064 159938 433116 159944
rect 432696 159452 432748 159458
rect 432696 159394 432748 159400
rect 433076 156874 433104 159938
rect 433536 159526 433564 163200
rect 433524 159520 433576 159526
rect 433524 159462 433576 159468
rect 434364 159390 434392 163200
rect 434444 159656 434496 159662
rect 434444 159598 434496 159604
rect 433248 159384 433300 159390
rect 433248 159326 433300 159332
rect 434352 159384 434404 159390
rect 434352 159326 434404 159332
rect 433156 156936 433208 156942
rect 433156 156878 433208 156884
rect 433064 156868 433116 156874
rect 433064 156810 433116 156816
rect 432052 155236 432104 155242
rect 432052 155178 432104 155184
rect 431868 152924 431920 152930
rect 431868 152866 431920 152872
rect 431880 150226 431908 152866
rect 432064 151814 432092 155178
rect 432064 151786 432552 151814
rect 432524 150226 432552 151786
rect 433168 150226 433196 156878
rect 433260 155514 433288 159326
rect 433248 155508 433300 155514
rect 433248 155450 433300 155456
rect 433800 152856 433852 152862
rect 433800 152798 433852 152804
rect 433812 150226 433840 152798
rect 434456 150226 434484 159598
rect 435192 158030 435220 163200
rect 435824 159724 435876 159730
rect 435824 159666 435876 159672
rect 434720 158024 434772 158030
rect 434720 157966 434772 157972
rect 435180 158024 435232 158030
rect 435180 157966 435232 157972
rect 429948 150198 430022 150226
rect 430592 150198 430666 150226
rect 431236 150198 431310 150226
rect 431880 150198 431954 150226
rect 432524 150198 432598 150226
rect 433168 150198 433242 150226
rect 433812 150198 433886 150226
rect 434456 150198 434530 150226
rect 434732 150210 434760 157966
rect 435088 156800 435140 156806
rect 435088 156742 435140 156748
rect 435100 150226 435128 156742
rect 435836 153202 435864 159666
rect 436112 158846 436140 163200
rect 436940 163146 436968 163200
rect 437032 163146 437060 163254
rect 436940 163118 437060 163146
rect 436376 159588 436428 159594
rect 436376 159530 436428 159536
rect 436100 158840 436152 158846
rect 436100 158782 436152 158788
rect 436388 156806 436416 159530
rect 436376 156800 436428 156806
rect 436376 156742 436428 156748
rect 435824 153196 435876 153202
rect 435824 153138 435876 153144
rect 436376 152992 436428 152998
rect 436376 152934 436428 152940
rect 436388 150226 436416 152934
rect 437020 152788 437072 152794
rect 437020 152730 437072 152736
rect 437032 150226 437060 152730
rect 437400 152522 437428 163254
rect 437754 163200 437810 164400
rect 438582 163200 438638 164400
rect 439410 163200 439466 164400
rect 440238 163200 440294 164400
rect 441066 163200 441122 164400
rect 441986 163200 442042 164400
rect 442814 163200 442870 164400
rect 443642 163200 443698 164400
rect 444470 163200 444526 164400
rect 445298 163200 445354 164400
rect 446126 163200 446182 164400
rect 446954 163200 447010 164400
rect 447874 163200 447930 164400
rect 448702 163200 448758 164400
rect 449530 163200 449586 164400
rect 450358 163200 450414 164400
rect 451186 163200 451242 164400
rect 452014 163200 452070 164400
rect 452842 163200 452898 164400
rect 453762 163200 453818 164400
rect 454590 163200 454646 164400
rect 455418 163200 455474 164400
rect 456246 163200 456302 164400
rect 457074 163200 457130 164400
rect 457902 163200 457958 164400
rect 458730 163200 458786 164400
rect 459650 163200 459706 164400
rect 460478 163200 460534 164400
rect 461306 163200 461362 164400
rect 462134 163200 462190 164400
rect 462962 163200 463018 164400
rect 463790 163200 463846 164400
rect 464618 163200 464674 164400
rect 465538 163200 465594 164400
rect 466366 163200 466422 164400
rect 467194 163200 467250 164400
rect 468022 163200 468078 164400
rect 468850 163200 468906 164400
rect 469678 163200 469734 164400
rect 470506 163200 470562 164400
rect 471426 163200 471482 164400
rect 472254 163200 472310 164400
rect 473082 163200 473138 164400
rect 473910 163200 473966 164400
rect 474738 163200 474794 164400
rect 475566 163200 475622 164400
rect 476394 163200 476450 164400
rect 477314 163200 477370 164400
rect 478142 163200 478198 164400
rect 478970 163200 479026 164400
rect 479798 163200 479854 164400
rect 480626 163200 480682 164400
rect 481454 163200 481510 164400
rect 482282 163200 482338 164400
rect 483202 163200 483258 164400
rect 484030 163200 484086 164400
rect 484136 163254 484348 163282
rect 437768 158982 437796 163200
rect 437756 158976 437808 158982
rect 437756 158918 437808 158924
rect 438308 153944 438360 153950
rect 438308 153886 438360 153892
rect 437664 153876 437716 153882
rect 437664 153818 437716 153824
rect 437388 152516 437440 152522
rect 437388 152458 437440 152464
rect 437676 150226 437704 153818
rect 438320 150226 438348 153886
rect 438596 153882 438624 163200
rect 438860 158840 438912 158846
rect 438860 158782 438912 158788
rect 438872 154222 438900 158782
rect 439424 158302 439452 163200
rect 439412 158296 439464 158302
rect 439412 158238 439464 158244
rect 438952 156732 439004 156738
rect 438952 156674 439004 156680
rect 438860 154216 438912 154222
rect 438860 154158 438912 154164
rect 438584 153876 438636 153882
rect 438584 153818 438636 153824
rect 438964 150226 438992 156674
rect 440252 153950 440280 163200
rect 441080 159662 441108 163200
rect 441068 159656 441120 159662
rect 441068 159598 441120 159604
rect 440332 158092 440384 158098
rect 440332 158034 440384 158040
rect 440240 153944 440292 153950
rect 440240 153886 440292 153892
rect 439596 153196 439648 153202
rect 439596 153138 439648 153144
rect 439608 150226 439636 153138
rect 440344 150226 440372 158034
rect 441712 155372 441764 155378
rect 441712 155314 441764 155320
rect 440884 155304 440936 155310
rect 440884 155246 440936 155252
rect 429350 149940 429378 150198
rect 429994 149940 430022 150198
rect 430638 149940 430666 150198
rect 431282 149940 431310 150198
rect 431926 149940 431954 150198
rect 432570 149940 432598 150198
rect 433214 149940 433242 150198
rect 433858 149940 433886 150198
rect 434502 149940 434530 150198
rect 434720 150204 434772 150210
rect 435100 150198 435174 150226
rect 434720 150146 434772 150152
rect 435146 149940 435174 150198
rect 435778 150204 435830 150210
rect 436388 150198 436462 150226
rect 437032 150198 437106 150226
rect 437676 150198 437750 150226
rect 438320 150198 438394 150226
rect 438964 150198 439038 150226
rect 439608 150198 439682 150226
rect 435778 150146 435830 150152
rect 435790 149940 435818 150146
rect 436434 149940 436462 150198
rect 437078 149940 437106 150198
rect 437722 149940 437750 150198
rect 438366 149940 438394 150198
rect 439010 149940 439038 150198
rect 439654 149940 439682 150198
rect 440298 150198 440372 150226
rect 440896 150226 440924 155246
rect 441436 154080 441488 154086
rect 441436 154022 441488 154028
rect 441448 151814 441476 154022
rect 441448 151786 441568 151814
rect 441540 150226 441568 151786
rect 440896 150198 440970 150226
rect 441540 150198 441614 150226
rect 441724 150210 441752 155314
rect 442000 155310 442028 163200
rect 442172 157004 442224 157010
rect 442172 156946 442224 156952
rect 441988 155304 442040 155310
rect 441988 155246 442040 155252
rect 442184 150226 442212 156946
rect 442828 155242 442856 163200
rect 443000 158228 443052 158234
rect 443000 158170 443052 158176
rect 442816 155236 442868 155242
rect 442816 155178 442868 155184
rect 440298 149940 440326 150198
rect 440942 149940 440970 150198
rect 441586 149940 441614 150198
rect 441712 150204 441764 150210
rect 442184 150198 442258 150226
rect 443012 150210 443040 158170
rect 443656 158098 443684 163200
rect 444288 158976 444340 158982
rect 444288 158918 444340 158924
rect 443644 158092 443696 158098
rect 443644 158034 443696 158040
rect 443460 154012 443512 154018
rect 443460 153954 443512 153960
rect 443472 150226 443500 153954
rect 444300 152726 444328 158918
rect 444380 156664 444432 156670
rect 444380 156606 444432 156612
rect 444288 152720 444340 152726
rect 444288 152662 444340 152668
rect 441712 150146 441764 150152
rect 442230 149940 442258 150198
rect 442862 150204 442914 150210
rect 442862 150146 442914 150152
rect 443000 150204 443052 150210
rect 443472 150198 443546 150226
rect 444392 150210 444420 156606
rect 444484 155378 444512 163200
rect 445312 156670 445340 163200
rect 445668 159656 445720 159662
rect 445668 159598 445720 159604
rect 445300 156664 445352 156670
rect 445300 156606 445352 156612
rect 444748 155508 444800 155514
rect 444748 155450 444800 155456
rect 444472 155372 444524 155378
rect 444472 155314 444524 155320
rect 444760 150226 444788 155450
rect 445680 152658 445708 159598
rect 446140 159186 446168 163200
rect 446128 159180 446180 159186
rect 446128 159122 446180 159128
rect 445760 158160 445812 158166
rect 445760 158102 445812 158108
rect 445668 152652 445720 152658
rect 445668 152594 445720 152600
rect 445772 151814 445800 158102
rect 446680 155440 446732 155446
rect 446680 155382 446732 155388
rect 445772 151786 446076 151814
rect 446048 150226 446076 151786
rect 446692 150226 446720 155382
rect 446968 152590 446996 163200
rect 447888 159662 447916 163200
rect 447876 159656 447928 159662
rect 447876 159598 447928 159604
rect 448716 159458 448744 163200
rect 449544 159594 449572 163200
rect 450372 160002 450400 163200
rect 450360 159996 450412 160002
rect 450360 159938 450412 159944
rect 451200 159798 451228 163200
rect 451188 159792 451240 159798
rect 451188 159734 451240 159740
rect 449532 159588 449584 159594
rect 449532 159530 449584 159536
rect 449808 159520 449860 159526
rect 449808 159462 449860 159468
rect 447140 159452 447192 159458
rect 447140 159394 447192 159400
rect 448704 159452 448756 159458
rect 448704 159394 448756 159400
rect 447152 153202 447180 159394
rect 447324 156868 447376 156874
rect 447324 156810 447376 156816
rect 447140 153196 447192 153202
rect 447140 153138 447192 153144
rect 446956 152584 447008 152590
rect 446956 152526 447008 152532
rect 447336 150226 447364 156810
rect 448612 156800 448664 156806
rect 448612 156742 448664 156748
rect 447968 154148 448020 154154
rect 447968 154090 448020 154096
rect 447980 150226 448008 154090
rect 448624 150226 448652 156742
rect 449256 153196 449308 153202
rect 449256 153138 449308 153144
rect 449268 150226 449296 153138
rect 449820 151814 449848 159462
rect 452028 159390 452056 163200
rect 450084 159384 450136 159390
rect 450084 159326 450136 159332
rect 452016 159384 452068 159390
rect 452016 159326 452068 159332
rect 450096 151814 450124 159326
rect 452856 158778 452884 163200
rect 453776 159526 453804 163200
rect 453764 159520 453816 159526
rect 453764 159462 453816 159468
rect 454604 158982 454632 163200
rect 455432 159050 455460 163200
rect 456064 159996 456116 160002
rect 456064 159938 456116 159944
rect 455420 159044 455472 159050
rect 455420 158986 455472 158992
rect 454592 158976 454644 158982
rect 454592 158918 454644 158924
rect 452844 158772 452896 158778
rect 452844 158714 452896 158720
rect 454408 158296 454460 158302
rect 454408 158238 454460 158244
rect 451188 158024 451240 158030
rect 451188 157966 451240 157972
rect 449820 151786 449940 151814
rect 450096 151786 450584 151814
rect 449912 150226 449940 151786
rect 450556 150226 450584 151786
rect 451200 150226 451228 157966
rect 451832 154216 451884 154222
rect 451832 154158 451884 154164
rect 451844 150226 451872 154158
rect 453764 153876 453816 153882
rect 453764 153818 453816 153824
rect 453120 152720 453172 152726
rect 453120 152662 453172 152668
rect 452476 152516 452528 152522
rect 452476 152458 452528 152464
rect 452488 150226 452516 152458
rect 453132 150226 453160 152662
rect 453776 150226 453804 153818
rect 454420 150226 454448 158238
rect 455972 155304 456024 155310
rect 455972 155246 456024 155252
rect 455052 153944 455104 153950
rect 455052 153886 455104 153892
rect 455064 150226 455092 153886
rect 455696 152652 455748 152658
rect 455696 152594 455748 152600
rect 455708 150226 455736 152594
rect 455984 151814 456012 155246
rect 456076 151910 456104 159938
rect 456260 158914 456288 163200
rect 457088 160070 457116 163200
rect 457076 160064 457128 160070
rect 457076 160006 457128 160012
rect 457916 160002 457944 163200
rect 457904 159996 457956 160002
rect 457904 159938 457956 159944
rect 458744 159730 458772 163200
rect 458732 159724 458784 159730
rect 458732 159666 458784 159672
rect 458364 159180 458416 159186
rect 458364 159122 458416 159128
rect 456248 158908 456300 158914
rect 456248 158850 456300 158856
rect 456800 158092 456852 158098
rect 456800 158034 456852 158040
rect 456064 151904 456116 151910
rect 456064 151846 456116 151852
rect 455984 151786 456380 151814
rect 456352 150226 456380 151786
rect 443000 150146 443052 150152
rect 442874 149940 442902 150146
rect 443518 149940 443546 150198
rect 444150 150204 444202 150210
rect 444150 150146 444202 150152
rect 444380 150204 444432 150210
rect 444760 150198 444834 150226
rect 444380 150146 444432 150152
rect 444162 149940 444190 150146
rect 444806 149940 444834 150198
rect 445438 150204 445490 150210
rect 446048 150198 446122 150226
rect 446692 150198 446766 150226
rect 447336 150198 447410 150226
rect 447980 150198 448054 150226
rect 448624 150198 448698 150226
rect 449268 150198 449342 150226
rect 449912 150198 449986 150226
rect 450556 150198 450630 150226
rect 451200 150198 451274 150226
rect 451844 150198 451918 150226
rect 452488 150198 452562 150226
rect 453132 150198 453206 150226
rect 453776 150198 453850 150226
rect 454420 150198 454494 150226
rect 455064 150198 455138 150226
rect 455708 150198 455782 150226
rect 456352 150198 456426 150226
rect 456812 150210 456840 158034
rect 458180 155372 458232 155378
rect 458180 155314 458232 155320
rect 456984 155236 457036 155242
rect 456984 155178 457036 155184
rect 456996 150226 457024 155178
rect 458192 150226 458220 155314
rect 445438 150146 445490 150152
rect 445450 149940 445478 150146
rect 446094 149940 446122 150198
rect 446738 149940 446766 150198
rect 447382 149940 447410 150198
rect 448026 149940 448054 150198
rect 448670 149940 448698 150198
rect 449314 149940 449342 150198
rect 449958 149940 449986 150198
rect 450602 149940 450630 150198
rect 451246 149940 451274 150198
rect 451890 149940 451918 150198
rect 452534 149940 452562 150198
rect 453178 149940 453206 150198
rect 453822 149940 453850 150198
rect 454466 149940 454494 150198
rect 455110 149940 455138 150198
rect 455754 149940 455782 150198
rect 456398 149940 456426 150198
rect 456800 150204 456852 150210
rect 456996 150198 457070 150226
rect 456800 150146 456852 150152
rect 457042 149940 457070 150198
rect 457674 150204 457726 150210
rect 458192 150198 458266 150226
rect 458376 150210 458404 159122
rect 459664 159118 459692 163200
rect 460204 159656 460256 159662
rect 460204 159598 460256 159604
rect 459652 159112 459704 159118
rect 459652 159054 459704 159060
rect 460112 158772 460164 158778
rect 460112 158714 460164 158720
rect 458824 156664 458876 156670
rect 458824 156606 458876 156612
rect 458836 150226 458864 156606
rect 460124 152590 460152 158714
rect 460020 152584 460072 152590
rect 460020 152526 460072 152532
rect 460112 152584 460164 152590
rect 460112 152526 460164 152532
rect 460032 151814 460060 152526
rect 460216 151814 460244 159598
rect 460492 159254 460520 163200
rect 460940 159452 460992 159458
rect 460940 159394 460992 159400
rect 460480 159248 460532 159254
rect 460480 159190 460532 159196
rect 460952 151814 460980 159394
rect 461320 159322 461348 163200
rect 461492 159588 461544 159594
rect 461492 159530 461544 159536
rect 461308 159316 461360 159322
rect 461308 159258 461360 159264
rect 461504 151814 461532 159530
rect 461584 158976 461636 158982
rect 461584 158918 461636 158924
rect 461596 153202 461624 158918
rect 462148 158778 462176 163200
rect 462872 159792 462924 159798
rect 462872 159734 462924 159740
rect 462136 158772 462188 158778
rect 462136 158714 462188 158720
rect 461584 153196 461636 153202
rect 461584 153138 461636 153144
rect 462688 151904 462740 151910
rect 462688 151846 462740 151852
rect 460032 151786 460152 151814
rect 460216 151786 460796 151814
rect 460952 151786 461440 151814
rect 461504 151786 462084 151814
rect 460124 150226 460152 151786
rect 460768 150226 460796 151786
rect 461412 150226 461440 151786
rect 462056 150226 462084 151786
rect 462700 150226 462728 151846
rect 462884 151814 462912 159734
rect 462976 159186 463004 163200
rect 463804 159798 463832 163200
rect 464344 160064 464396 160070
rect 464344 160006 464396 160012
rect 463792 159792 463844 159798
rect 463792 159734 463844 159740
rect 463976 159384 464028 159390
rect 463976 159326 464028 159332
rect 462964 159180 463016 159186
rect 462964 159122 463016 159128
rect 462964 159044 463016 159050
rect 462964 158986 463016 158992
rect 462976 153066 463004 158986
rect 463148 158908 463200 158914
rect 463148 158850 463200 158856
rect 463160 153134 463188 158850
rect 463148 153128 463200 153134
rect 463148 153070 463200 153076
rect 462964 153060 463016 153066
rect 462964 153002 463016 153008
rect 462884 151786 463372 151814
rect 463344 150226 463372 151786
rect 463988 150226 464016 159326
rect 464356 151910 464384 160006
rect 464632 158846 464660 163200
rect 464712 159996 464764 160002
rect 464712 159938 464764 159944
rect 464620 158840 464672 158846
rect 464620 158782 464672 158788
rect 464724 152930 464752 159938
rect 465080 159724 465132 159730
rect 465080 159666 465132 159672
rect 465092 152998 465120 159666
rect 465264 159520 465316 159526
rect 465264 159462 465316 159468
rect 465080 152992 465132 152998
rect 465080 152934 465132 152940
rect 464712 152924 464764 152930
rect 464712 152866 464764 152872
rect 464620 152584 464672 152590
rect 464620 152526 464672 152532
rect 464344 151904 464396 151910
rect 464344 151846 464396 151852
rect 464632 150226 464660 152526
rect 465276 150226 465304 159462
rect 465552 158914 465580 163200
rect 466380 158982 466408 163200
rect 467208 159526 467236 163200
rect 468036 159662 468064 163200
rect 468024 159656 468076 159662
rect 468024 159598 468076 159604
rect 467196 159520 467248 159526
rect 467196 159462 467248 159468
rect 468864 159458 468892 163200
rect 468852 159452 468904 159458
rect 468852 159394 468904 159400
rect 469692 159390 469720 163200
rect 470520 159594 470548 163200
rect 470508 159588 470560 159594
rect 470508 159530 470560 159536
rect 469680 159384 469732 159390
rect 469680 159326 469732 159332
rect 467932 159316 467984 159322
rect 467932 159258 467984 159264
rect 466644 159248 466696 159254
rect 466644 159190 466696 159196
rect 466460 159112 466512 159118
rect 466460 159054 466512 159060
rect 466368 158976 466420 158982
rect 466368 158918 466420 158924
rect 465540 158908 465592 158914
rect 465540 158850 465592 158856
rect 466472 153202 466500 159054
rect 465908 153196 465960 153202
rect 465908 153138 465960 153144
rect 466460 153196 466512 153202
rect 466460 153138 466512 153144
rect 465920 150226 465948 153138
rect 466656 153066 466684 159190
rect 467840 158772 467892 158778
rect 467840 158714 467892 158720
rect 467196 153128 467248 153134
rect 467196 153070 467248 153076
rect 466552 153060 466604 153066
rect 466552 153002 466604 153008
rect 466644 153060 466696 153066
rect 466644 153002 466696 153008
rect 466564 150226 466592 153002
rect 467208 150226 467236 153070
rect 467852 152046 467880 158714
rect 467840 152040 467892 152046
rect 467840 151982 467892 151988
rect 467944 151910 467972 159258
rect 469220 159180 469272 159186
rect 469220 159122 469272 159128
rect 469128 152992 469180 152998
rect 469128 152934 469180 152940
rect 468392 152924 468444 152930
rect 468392 152866 468444 152872
rect 467840 151904 467892 151910
rect 467840 151846 467892 151852
rect 467932 151904 467984 151910
rect 467932 151846 467984 151852
rect 467852 150226 467880 151846
rect 468404 151814 468432 152866
rect 468404 151786 468524 151814
rect 468496 150226 468524 151786
rect 469140 150226 469168 152934
rect 469232 151978 469260 159122
rect 471440 159118 471468 163200
rect 472268 159866 472296 163200
rect 472256 159860 472308 159866
rect 472256 159802 472308 159808
rect 471796 159792 471848 159798
rect 471796 159734 471848 159740
rect 471428 159112 471480 159118
rect 471428 159054 471480 159060
rect 471612 158840 471664 158846
rect 471612 158782 471664 158788
rect 471624 153202 471652 158782
rect 469772 153196 469824 153202
rect 469772 153138 469824 153144
rect 471612 153196 471664 153202
rect 471612 153138 471664 153144
rect 469220 151972 469272 151978
rect 469220 151914 469272 151920
rect 469784 150226 469812 153138
rect 470416 153060 470468 153066
rect 470416 153002 470468 153008
rect 470428 150226 470456 153002
rect 471808 152998 471836 159734
rect 472808 158976 472860 158982
rect 472808 158918 472860 158924
rect 471980 158908 472032 158914
rect 471980 158850 472032 158856
rect 471992 153134 472020 158850
rect 471980 153128 472032 153134
rect 471980 153070 472032 153076
rect 472820 153066 472848 158918
rect 473096 158778 473124 163200
rect 473360 159520 473412 159526
rect 473360 159462 473412 159468
rect 473084 158772 473136 158778
rect 473084 158714 473136 158720
rect 472808 153060 472860 153066
rect 472808 153002 472860 153008
rect 473372 152998 473400 159462
rect 473924 159050 473952 163200
rect 473912 159044 473964 159050
rect 473912 158986 473964 158992
rect 474752 158914 474780 163200
rect 474832 159452 474884 159458
rect 474832 159394 474884 159400
rect 474740 158908 474792 158914
rect 474740 158850 474792 158856
rect 474844 153202 474872 159394
rect 475580 158982 475608 163200
rect 476028 159656 476080 159662
rect 476028 159598 476080 159604
rect 475568 158976 475620 158982
rect 475568 158918 475620 158924
rect 473636 153196 473688 153202
rect 473636 153138 473688 153144
rect 474832 153196 474884 153202
rect 474832 153138 474884 153144
rect 471796 152992 471848 152998
rect 471796 152934 471848 152940
rect 472992 152992 473044 152998
rect 472992 152934 473044 152940
rect 473360 152992 473412 152998
rect 473360 152934 473412 152940
rect 471704 152040 471756 152046
rect 471704 151982 471756 151988
rect 471060 151904 471112 151910
rect 471060 151846 471112 151852
rect 471072 150226 471100 151846
rect 471716 150226 471744 151982
rect 472348 151972 472400 151978
rect 472348 151914 472400 151920
rect 472360 150226 472388 151914
rect 473004 150226 473032 152934
rect 473648 150226 473676 153138
rect 474280 153128 474332 153134
rect 474280 153070 474332 153076
rect 474292 150226 474320 153070
rect 474924 153060 474976 153066
rect 474924 153002 474976 153008
rect 474936 150226 474964 153002
rect 475568 152992 475620 152998
rect 475568 152934 475620 152940
rect 475580 150226 475608 152934
rect 476040 151814 476068 159598
rect 476120 159588 476172 159594
rect 476120 159530 476172 159536
rect 476132 153134 476160 159530
rect 476408 158846 476436 163200
rect 477328 159458 477356 163200
rect 477316 159452 477368 159458
rect 477316 159394 477368 159400
rect 478156 159390 478184 163200
rect 478984 159798 479012 163200
rect 479812 159866 479840 163200
rect 479432 159860 479484 159866
rect 479432 159802 479484 159808
rect 479800 159860 479852 159866
rect 479800 159802 479852 159808
rect 478972 159792 479024 159798
rect 478972 159734 479024 159740
rect 477408 159384 477460 159390
rect 477408 159326 477460 159332
rect 478144 159384 478196 159390
rect 478144 159326 478196 159332
rect 476396 158840 476448 158846
rect 476396 158782 476448 158788
rect 476948 153196 477000 153202
rect 476948 153138 477000 153144
rect 476120 153128 476172 153134
rect 476120 153070 476172 153076
rect 476040 151786 476252 151814
rect 476224 150226 476252 151786
rect 476960 150226 476988 153138
rect 477420 151814 477448 159326
rect 477684 159112 477736 159118
rect 477684 159054 477736 159060
rect 477420 151786 477540 151814
rect 457674 150146 457726 150152
rect 457686 149940 457714 150146
rect 458238 149940 458266 150198
rect 458364 150204 458416 150210
rect 458836 150198 458910 150226
rect 458364 150146 458416 150152
rect 458882 149940 458910 150198
rect 459514 150204 459566 150210
rect 460124 150198 460198 150226
rect 460768 150198 460842 150226
rect 461412 150198 461486 150226
rect 462056 150198 462130 150226
rect 462700 150198 462774 150226
rect 463344 150198 463418 150226
rect 463988 150198 464062 150226
rect 464632 150198 464706 150226
rect 465276 150198 465350 150226
rect 465920 150198 465994 150226
rect 466564 150198 466638 150226
rect 467208 150198 467282 150226
rect 467852 150198 467926 150226
rect 468496 150198 468570 150226
rect 469140 150198 469214 150226
rect 469784 150198 469858 150226
rect 470428 150198 470502 150226
rect 471072 150198 471146 150226
rect 471716 150198 471790 150226
rect 472360 150198 472434 150226
rect 473004 150198 473078 150226
rect 473648 150198 473722 150226
rect 474292 150198 474366 150226
rect 474936 150198 475010 150226
rect 475580 150198 475654 150226
rect 476224 150198 476298 150226
rect 459514 150146 459566 150152
rect 459526 149940 459554 150146
rect 460170 149940 460198 150198
rect 460814 149940 460842 150198
rect 461458 149940 461486 150198
rect 462102 149940 462130 150198
rect 462746 149940 462774 150198
rect 463390 149940 463418 150198
rect 464034 149940 464062 150198
rect 464678 149940 464706 150198
rect 465322 149940 465350 150198
rect 465966 149940 465994 150198
rect 466610 149940 466638 150198
rect 467254 149940 467282 150198
rect 467898 149940 467926 150198
rect 468542 149940 468570 150198
rect 469186 149940 469214 150198
rect 469830 149940 469858 150198
rect 470474 149940 470502 150198
rect 471118 149940 471146 150198
rect 471762 149940 471790 150198
rect 472406 149940 472434 150198
rect 473050 149940 473078 150198
rect 473694 149940 473722 150198
rect 474338 149940 474366 150198
rect 474982 149940 475010 150198
rect 475626 149940 475654 150198
rect 476270 149940 476298 150198
rect 476914 150198 476988 150226
rect 477512 150226 477540 151786
rect 477512 150198 477586 150226
rect 477696 150210 477724 159054
rect 478972 158772 479024 158778
rect 478972 158714 479024 158720
rect 478144 153128 478196 153134
rect 478144 153070 478196 153076
rect 478156 150226 478184 153070
rect 476914 149940 476942 150198
rect 477558 149940 477586 150198
rect 477684 150204 477736 150210
rect 478156 150198 478230 150226
rect 478984 150210 479012 158714
rect 479444 150226 479472 159802
rect 480640 158914 480668 163200
rect 480720 159044 480772 159050
rect 480720 158986 480772 158992
rect 480260 158908 480312 158914
rect 480260 158850 480312 158856
rect 480628 158908 480680 158914
rect 480628 158850 480680 158856
rect 477684 150146 477736 150152
rect 478202 149940 478230 150198
rect 478834 150204 478886 150210
rect 478834 150146 478886 150152
rect 478972 150204 479024 150210
rect 479444 150198 479518 150226
rect 480272 150210 480300 158850
rect 480732 150226 480760 158986
rect 481468 158778 481496 163200
rect 482296 159526 482324 163200
rect 482284 159520 482336 159526
rect 482284 159462 482336 159468
rect 482008 158976 482060 158982
rect 482008 158918 482060 158924
rect 481640 158840 481692 158846
rect 481640 158782 481692 158788
rect 481456 158772 481508 158778
rect 481456 158714 481508 158720
rect 478972 150146 479024 150152
rect 478846 149940 478874 150146
rect 479490 149940 479518 150198
rect 480122 150204 480174 150210
rect 480122 150146 480174 150152
rect 480260 150204 480312 150210
rect 480732 150198 480806 150226
rect 481652 150210 481680 158782
rect 482020 150226 482048 158918
rect 483216 152998 483244 163200
rect 484044 163146 484072 163200
rect 484136 163146 484164 163254
rect 484044 163118 484164 163146
rect 483296 159452 483348 159458
rect 483296 159394 483348 159400
rect 483204 152992 483256 152998
rect 483204 152934 483256 152940
rect 483308 150226 483336 159394
rect 483940 159384 483992 159390
rect 483940 159326 483992 159332
rect 483952 150226 483980 159326
rect 484320 153066 484348 163254
rect 484858 163200 484914 164400
rect 485686 163200 485742 164400
rect 486514 163200 486570 164400
rect 487342 163200 487398 164400
rect 488170 163200 488226 164400
rect 489090 163200 489146 164400
rect 489918 163200 489974 164400
rect 490746 163200 490802 164400
rect 491574 163200 491630 164400
rect 492402 163200 492458 164400
rect 493230 163200 493286 164400
rect 494058 163200 494114 164400
rect 494978 163200 495034 164400
rect 495084 163254 495296 163282
rect 484584 159792 484636 159798
rect 484584 159734 484636 159740
rect 484308 153060 484360 153066
rect 484308 153002 484360 153008
rect 484596 150226 484624 159734
rect 484872 153134 484900 163200
rect 485228 159860 485280 159866
rect 485228 159802 485280 159808
rect 484860 153128 484912 153134
rect 484860 153070 484912 153076
rect 485240 150226 485268 159802
rect 485700 153202 485728 163200
rect 485964 158908 486016 158914
rect 485964 158850 486016 158856
rect 485688 153196 485740 153202
rect 485688 153138 485740 153144
rect 485976 150226 486004 158850
rect 486424 158772 486476 158778
rect 486424 158714 486476 158720
rect 486436 151814 486464 158714
rect 486528 151910 486556 163200
rect 487252 159520 487304 159526
rect 487252 159462 487304 159468
rect 486516 151904 486568 151910
rect 486516 151846 486568 151852
rect 486436 151786 486556 151814
rect 480260 150146 480312 150152
rect 480134 149940 480162 150146
rect 480778 149940 480806 150198
rect 481410 150204 481462 150210
rect 481410 150146 481462 150152
rect 481640 150204 481692 150210
rect 482020 150198 482094 150226
rect 481640 150146 481692 150152
rect 481422 149940 481450 150146
rect 482066 149940 482094 150198
rect 482698 150204 482750 150210
rect 483308 150198 483382 150226
rect 483952 150198 484026 150226
rect 484596 150198 484670 150226
rect 485240 150198 485314 150226
rect 482698 150146 482750 150152
rect 482710 149940 482738 150146
rect 483354 149940 483382 150198
rect 483998 149940 484026 150198
rect 484642 149940 484670 150198
rect 485286 149940 485314 150198
rect 485930 150198 486004 150226
rect 486528 150226 486556 151786
rect 487264 150226 487292 159462
rect 487356 151978 487384 163200
rect 487804 152992 487856 152998
rect 487804 152934 487856 152940
rect 487344 151972 487396 151978
rect 487344 151914 487396 151920
rect 486528 150198 486602 150226
rect 485930 149940 485958 150198
rect 486574 149940 486602 150198
rect 487218 150198 487292 150226
rect 487816 150226 487844 152934
rect 488184 152046 488212 163200
rect 489000 153128 489052 153134
rect 489000 153070 489052 153076
rect 488264 153060 488316 153066
rect 488264 153002 488316 153008
rect 488172 152040 488224 152046
rect 488172 151982 488224 151988
rect 488276 151814 488304 153002
rect 488276 151786 488488 151814
rect 488460 150226 488488 151786
rect 489012 150226 489040 153070
rect 489104 151910 489132 163200
rect 489644 153196 489696 153202
rect 489644 153138 489696 153144
rect 489092 151904 489144 151910
rect 489092 151846 489144 151852
rect 489656 150226 489684 153138
rect 489932 153134 489960 163200
rect 490760 153202 490788 163200
rect 490748 153196 490800 153202
rect 490748 153138 490800 153144
rect 489920 153128 489972 153134
rect 489920 153070 489972 153076
rect 491588 152998 491616 163200
rect 492416 153066 492444 163200
rect 493244 153134 493272 163200
rect 494072 153202 494100 163200
rect 494992 163146 495020 163200
rect 495084 163146 495112 163254
rect 494992 163118 495112 163146
rect 493508 153196 493560 153202
rect 493508 153138 493560 153144
rect 494060 153196 494112 153202
rect 494060 153138 494112 153144
rect 492864 153128 492916 153134
rect 492864 153070 492916 153076
rect 493232 153128 493284 153134
rect 493232 153070 493284 153076
rect 492404 153060 492456 153066
rect 492404 153002 492456 153008
rect 491576 152992 491628 152998
rect 491576 152934 491628 152940
rect 491576 152040 491628 152046
rect 491576 151982 491628 151988
rect 490932 151972 490984 151978
rect 490932 151914 490984 151920
rect 490288 151836 490340 151842
rect 490288 151778 490340 151784
rect 490300 150226 490328 151778
rect 490944 150226 490972 151914
rect 491588 150226 491616 151982
rect 492220 151904 492272 151910
rect 492220 151846 492272 151852
rect 492232 150226 492260 151846
rect 492876 150226 492904 153070
rect 493520 150226 493548 153138
rect 495268 153066 495296 163254
rect 495806 163200 495862 164400
rect 496634 163200 496690 164400
rect 497462 163200 497518 164400
rect 498290 163200 498346 164400
rect 499118 163200 499174 164400
rect 499224 163254 499528 163282
rect 495820 153134 495848 163200
rect 496648 153202 496676 163200
rect 496084 153196 496136 153202
rect 496084 153138 496136 153144
rect 496636 153196 496688 153202
rect 496636 153138 496688 153144
rect 495440 153128 495492 153134
rect 495440 153070 495492 153076
rect 495808 153128 495860 153134
rect 495808 153070 495860 153076
rect 494796 153060 494848 153066
rect 494796 153002 494848 153008
rect 495256 153060 495308 153066
rect 495256 153002 495308 153008
rect 494152 152992 494204 152998
rect 494152 152934 494204 152940
rect 494164 150226 494192 152934
rect 494808 150226 494836 153002
rect 495452 150226 495480 153070
rect 496096 150226 496124 153138
rect 497476 153134 497504 163200
rect 498304 153202 498332 163200
rect 499132 163146 499160 163200
rect 499224 163146 499252 163254
rect 499132 163118 499252 163146
rect 498016 153196 498068 153202
rect 498016 153138 498068 153144
rect 498292 153196 498344 153202
rect 498292 153138 498344 153144
rect 499304 153196 499356 153202
rect 499304 153138 499356 153144
rect 497372 153128 497424 153134
rect 497372 153070 497424 153076
rect 497464 153128 497516 153134
rect 497464 153070 497516 153076
rect 496728 153060 496780 153066
rect 496728 153002 496780 153008
rect 496740 150226 496768 153002
rect 497384 150226 497412 153070
rect 498028 150226 498056 153138
rect 498660 153128 498712 153134
rect 498660 153070 498712 153076
rect 498672 150226 498700 153070
rect 499316 150226 499344 153138
rect 499500 151910 499528 163254
rect 499946 163200 500002 164400
rect 500866 163200 500922 164400
rect 500972 163254 501644 163282
rect 499960 158846 499988 163200
rect 499948 158840 500000 158846
rect 499948 158782 500000 158788
rect 500592 158840 500644 158846
rect 500592 158782 500644 158788
rect 499488 151904 499540 151910
rect 499488 151846 499540 151852
rect 499948 151904 500000 151910
rect 499948 151846 500000 151852
rect 499960 150226 499988 151846
rect 500604 150226 500632 158782
rect 500880 151814 500908 163200
rect 500972 153202 501000 163254
rect 501616 163146 501644 163254
rect 501694 163200 501750 164400
rect 502522 163200 502578 164400
rect 503350 163200 503406 164400
rect 503824 163254 504128 163282
rect 501708 163146 501736 163200
rect 501616 163118 501736 163146
rect 500960 153196 501012 153202
rect 500960 153138 501012 153144
rect 501880 153196 501932 153202
rect 501880 153138 501932 153144
rect 500880 151786 501276 151814
rect 501248 150226 501276 151786
rect 501892 150226 501920 153138
rect 502536 150226 502564 163200
rect 503364 151814 503392 163200
rect 503272 151786 503392 151814
rect 503272 150226 503300 151786
rect 487816 150198 487890 150226
rect 488460 150198 488534 150226
rect 489012 150198 489086 150226
rect 489656 150198 489730 150226
rect 490300 150198 490374 150226
rect 490944 150198 491018 150226
rect 491588 150198 491662 150226
rect 492232 150198 492306 150226
rect 492876 150198 492950 150226
rect 493520 150198 493594 150226
rect 494164 150198 494238 150226
rect 494808 150198 494882 150226
rect 495452 150198 495526 150226
rect 496096 150198 496170 150226
rect 496740 150198 496814 150226
rect 497384 150198 497458 150226
rect 498028 150198 498102 150226
rect 498672 150198 498746 150226
rect 499316 150198 499390 150226
rect 499960 150198 500034 150226
rect 500604 150198 500678 150226
rect 501248 150198 501322 150226
rect 501892 150198 501966 150226
rect 502536 150198 502610 150226
rect 487218 149940 487246 150198
rect 487862 149940 487890 150198
rect 488506 149940 488534 150198
rect 489058 149940 489086 150198
rect 489702 149940 489730 150198
rect 490346 149940 490374 150198
rect 490990 149940 491018 150198
rect 491634 149940 491662 150198
rect 492278 149940 492306 150198
rect 492922 149940 492950 150198
rect 493566 149940 493594 150198
rect 494210 149940 494238 150198
rect 494854 149940 494882 150198
rect 495498 149940 495526 150198
rect 496142 149940 496170 150198
rect 496786 149940 496814 150198
rect 497430 149940 497458 150198
rect 498074 149940 498102 150198
rect 498718 149940 498746 150198
rect 499362 149940 499390 150198
rect 500006 149940 500034 150198
rect 500650 149940 500678 150198
rect 501294 149940 501322 150198
rect 501938 149940 501966 150198
rect 502582 149940 502610 150198
rect 503226 150198 503300 150226
rect 503824 150226 503852 163254
rect 504100 163146 504128 163254
rect 504178 163200 504234 164400
rect 505006 163200 505062 164400
rect 505112 163254 505784 163282
rect 504192 163146 504220 163200
rect 504100 163118 504220 163146
rect 505020 158778 505048 163200
rect 504456 158772 504508 158778
rect 504456 158714 504508 158720
rect 505008 158772 505060 158778
rect 505008 158714 505060 158720
rect 504468 150226 504496 158714
rect 505112 150226 505140 163254
rect 505756 163146 505784 163254
rect 505834 163200 505890 164400
rect 506754 163200 506810 164400
rect 507582 163200 507638 164400
rect 508410 163200 508466 164400
rect 509238 163200 509294 164400
rect 510066 163200 510122 164400
rect 510894 163200 510950 164400
rect 511722 163200 511778 164400
rect 512012 163254 512592 163282
rect 505848 163146 505876 163200
rect 505756 163118 505876 163146
rect 506388 158840 506440 158846
rect 506388 158782 506440 158788
rect 505836 158772 505888 158778
rect 505836 158714 505888 158720
rect 505848 150226 505876 158714
rect 503824 150198 503898 150226
rect 504468 150198 504542 150226
rect 505112 150198 505186 150226
rect 503226 149940 503254 150198
rect 503870 149940 503898 150198
rect 504514 149940 504542 150198
rect 505158 149940 505186 150198
rect 505802 150198 505876 150226
rect 506400 150226 506428 158782
rect 506768 158778 506796 163200
rect 507124 159044 507176 159050
rect 507124 158986 507176 158992
rect 506756 158772 506808 158778
rect 506756 158714 506808 158720
rect 507136 150226 507164 158986
rect 507596 158846 507624 163200
rect 508424 159050 508452 163200
rect 508412 159044 508464 159050
rect 508412 158986 508464 158992
rect 508412 158908 508464 158914
rect 508412 158850 508464 158856
rect 507584 158840 507636 158846
rect 507584 158782 507636 158788
rect 507676 151972 507728 151978
rect 507676 151914 507728 151920
rect 506400 150198 506474 150226
rect 505802 149940 505830 150198
rect 506446 149940 506474 150198
rect 507090 150198 507164 150226
rect 507688 150226 507716 151914
rect 508424 150226 508452 158850
rect 509252 151978 509280 163200
rect 510080 158914 510108 163200
rect 510068 158908 510120 158914
rect 510068 158850 510120 158856
rect 509700 158772 509752 158778
rect 509700 158714 509752 158720
rect 509240 151972 509292 151978
rect 509240 151914 509292 151920
rect 509056 151836 509108 151842
rect 509056 151778 509108 151784
rect 509068 150226 509096 151778
rect 509712 150226 509740 158714
rect 510344 152856 510396 152862
rect 510344 152798 510396 152804
rect 510356 150226 510384 152798
rect 510908 151842 510936 163200
rect 511736 158778 511764 163200
rect 511724 158772 511776 158778
rect 511724 158714 511776 158720
rect 510988 153196 511040 153202
rect 510988 153138 511040 153144
rect 510896 151836 510948 151842
rect 510896 151778 510948 151784
rect 511000 150226 511028 153138
rect 512012 152862 512040 163254
rect 512564 163146 512592 163254
rect 512642 163200 512698 164400
rect 513470 163200 513526 164400
rect 513576 163254 514248 163282
rect 512656 163146 512684 163200
rect 512564 163118 512684 163146
rect 513484 153202 513512 163200
rect 513472 153196 513524 153202
rect 513472 153138 513524 153144
rect 512920 153128 512972 153134
rect 512920 153070 512972 153076
rect 512276 152992 512328 152998
rect 512276 152934 512328 152940
rect 512000 152856 512052 152862
rect 512000 152798 512052 152804
rect 511632 152380 511684 152386
rect 511632 152322 511684 152328
rect 511644 150226 511672 152322
rect 512288 150226 512316 152934
rect 512932 150226 512960 153070
rect 513576 152386 513604 163254
rect 514220 163146 514248 163254
rect 514298 163200 514354 164400
rect 514772 163254 515076 163282
rect 514312 163146 514340 163200
rect 514220 163118 514340 163146
rect 514208 153196 514260 153202
rect 514208 153138 514260 153144
rect 513564 152380 513616 152386
rect 513564 152322 513616 152328
rect 513564 152244 513616 152250
rect 513564 152186 513616 152192
rect 513576 150226 513604 152186
rect 514220 150226 514248 153138
rect 514772 152998 514800 163254
rect 515048 163146 515076 163254
rect 515126 163200 515182 164400
rect 515324 163254 515904 163282
rect 515140 163146 515168 163200
rect 515048 163118 515168 163146
rect 514852 158772 514904 158778
rect 514852 158714 514904 158720
rect 514760 152992 514812 152998
rect 514760 152934 514812 152940
rect 514864 150226 514892 158714
rect 515324 153134 515352 163254
rect 515876 163146 515904 163254
rect 515954 163200 516010 164400
rect 516152 163254 516732 163282
rect 515968 163146 515996 163200
rect 515876 163118 515996 163146
rect 515312 153128 515364 153134
rect 515312 153070 515364 153076
rect 516152 152250 516180 163254
rect 516704 163146 516732 163254
rect 516782 163200 516838 164400
rect 517610 163200 517666 164400
rect 518530 163200 518586 164400
rect 518912 163254 519308 163282
rect 516796 163146 516824 163200
rect 516704 163118 516824 163146
rect 517624 161474 517652 163200
rect 517532 161446 517652 161474
rect 517532 158794 517560 161446
rect 518072 159452 518124 159458
rect 518072 159394 518124 159400
rect 517440 158766 517560 158794
rect 517440 153202 517468 158766
rect 517428 153196 517480 153202
rect 517428 153138 517480 153144
rect 516140 152244 516192 152250
rect 516140 152186 516192 152192
rect 516692 152176 516744 152182
rect 516692 152118 516744 152124
rect 515496 152108 515548 152114
rect 515496 152050 515548 152056
rect 515508 150226 515536 152050
rect 515956 152040 516008 152046
rect 515956 151982 516008 151988
rect 515968 151814 515996 151982
rect 515968 151786 516088 151814
rect 507688 150198 507762 150226
rect 507090 149940 507118 150198
rect 507734 149940 507762 150198
rect 508378 150198 508452 150226
rect 509022 150198 509096 150226
rect 509666 150198 509740 150226
rect 510310 150198 510384 150226
rect 510954 150198 511028 150226
rect 511598 150198 511672 150226
rect 512242 150198 512316 150226
rect 512886 150198 512960 150226
rect 513530 150198 513604 150226
rect 514174 150198 514248 150226
rect 514818 150198 514892 150226
rect 515462 150198 515536 150226
rect 516060 150226 516088 151786
rect 516704 150226 516732 152118
rect 517428 151972 517480 151978
rect 517428 151914 517480 151920
rect 517440 150226 517468 151914
rect 518084 150226 518112 159394
rect 518544 158778 518572 163200
rect 518716 159384 518768 159390
rect 518716 159326 518768 159332
rect 518532 158772 518584 158778
rect 518532 158714 518584 158720
rect 518728 150226 518756 159326
rect 518912 152114 518940 163254
rect 519280 163146 519308 163254
rect 519358 163200 519414 164400
rect 519464 163254 520136 163282
rect 519372 163146 519400 163200
rect 519280 163118 519400 163146
rect 519358 158672 519414 158681
rect 519358 158607 519414 158616
rect 518900 152108 518952 152114
rect 518900 152050 518952 152056
rect 516060 150198 516134 150226
rect 516704 150198 516778 150226
rect 508378 149940 508406 150198
rect 509022 149940 509050 150198
rect 509666 149940 509694 150198
rect 510310 149940 510338 150198
rect 510954 149940 510982 150198
rect 511598 149940 511626 150198
rect 512242 149940 512270 150198
rect 512886 149940 512914 150198
rect 513530 149940 513558 150198
rect 514174 149940 514202 150198
rect 514818 149940 514846 150198
rect 515462 149940 515490 150198
rect 516106 149940 516134 150198
rect 516750 149940 516778 150198
rect 517394 150198 517468 150226
rect 518038 150198 518112 150226
rect 518682 150198 518756 150226
rect 517394 149940 517422 150198
rect 518038 149940 518066 150198
rect 518682 149940 518710 150198
rect 117228 149874 117280 149880
rect 117136 149864 117188 149870
rect 117136 149806 117188 149812
rect 117044 145580 117096 145586
rect 117044 145522 117096 145528
rect 116950 108760 117006 108769
rect 116950 108695 117006 108704
rect 117056 106865 117084 145522
rect 117148 110673 117176 149806
rect 117240 133657 117268 149874
rect 519372 145217 519400 158607
rect 519464 152046 519492 163254
rect 519726 163160 519782 163169
rect 520108 163146 520136 163254
rect 520186 163200 520242 164400
rect 520292 163254 520964 163282
rect 520200 163146 520228 163200
rect 520108 163118 520228 163146
rect 519726 163095 519782 163104
rect 519542 161664 519598 161673
rect 519542 161599 519598 161608
rect 519452 152040 519504 152046
rect 519452 151982 519504 151988
rect 519556 147937 519584 161599
rect 519634 160168 519690 160177
rect 519634 160103 519690 160112
rect 519542 147928 519598 147937
rect 519542 147863 519598 147872
rect 519648 146577 519676 160103
rect 519740 149297 519768 163095
rect 520094 157176 520150 157185
rect 520094 157111 520150 157120
rect 519910 154048 519966 154057
rect 519910 153983 519966 153992
rect 519818 151056 519874 151065
rect 519818 150991 519874 151000
rect 519726 149288 519782 149297
rect 519726 149223 519782 149232
rect 519726 148064 519782 148073
rect 519726 147999 519782 148008
rect 519634 146568 519690 146577
rect 519634 146503 519690 146512
rect 519358 145208 519414 145217
rect 519358 145143 519414 145152
rect 519542 144936 519598 144945
rect 519542 144871 519598 144880
rect 519266 143440 519322 143449
rect 519266 143375 519322 143384
rect 117226 133648 117282 133657
rect 117226 133583 117282 133592
rect 519280 131481 519308 143375
rect 519358 141944 519414 141953
rect 519358 141879 519414 141888
rect 519266 131472 519322 131481
rect 519266 131407 519322 131416
rect 519372 130121 519400 141879
rect 519450 140448 519506 140457
rect 519450 140383 519506 140392
rect 519358 130112 519414 130121
rect 519358 130047 519414 130056
rect 519464 128761 519492 140383
rect 519556 132977 519584 144871
rect 519740 135697 519768 147999
rect 519832 138417 519860 150991
rect 519924 141137 519952 153983
rect 520002 149560 520058 149569
rect 520002 149495 520058 149504
rect 519910 141128 519966 141137
rect 519910 141063 519966 141072
rect 519818 138408 519874 138417
rect 519818 138343 519874 138352
rect 520016 137057 520044 149495
rect 520108 143857 520136 157111
rect 520186 155680 520242 155689
rect 520186 155615 520242 155624
rect 520094 143848 520150 143857
rect 520094 143783 520150 143792
rect 520200 142497 520228 155615
rect 520292 152182 520320 163254
rect 520936 163146 520964 163254
rect 521014 163200 521070 164400
rect 521842 163200 521898 164400
rect 522670 163200 522726 164400
rect 523498 163200 523554 164400
rect 521028 163146 521056 163200
rect 520936 163118 521056 163146
rect 521856 161474 521884 163200
rect 521672 161446 521884 161474
rect 521672 158794 521700 161446
rect 522684 159458 522712 163200
rect 522672 159452 522724 159458
rect 522672 159394 522724 159400
rect 523512 159390 523540 163200
rect 523500 159384 523552 159390
rect 523500 159326 523552 159332
rect 521580 158766 521700 158794
rect 521014 152552 521070 152561
rect 521014 152487 521070 152496
rect 520280 152176 520332 152182
rect 520280 152118 520332 152124
rect 520922 146568 520978 146577
rect 520922 146503 520978 146512
rect 520186 142488 520242 142497
rect 520186 142423 520242 142432
rect 520094 138952 520150 138961
rect 520094 138887 520150 138896
rect 520002 137048 520058 137057
rect 520002 136983 520058 136992
rect 519910 135824 519966 135833
rect 519910 135759 519966 135768
rect 519726 135688 519782 135697
rect 519726 135623 519782 135632
rect 519634 134328 519690 134337
rect 519634 134263 519690 134272
rect 519542 132968 519598 132977
rect 519542 132903 519598 132912
rect 519542 131336 519598 131345
rect 519542 131271 519598 131280
rect 519450 128752 519506 128761
rect 519450 128687 519506 128696
rect 519450 128344 519506 128353
rect 519450 128279 519506 128288
rect 519358 123720 519414 123729
rect 519358 123655 519414 123664
rect 519266 119096 519322 119105
rect 519266 119031 519322 119040
rect 117134 110664 117190 110673
rect 117134 110599 117190 110608
rect 519280 109585 519308 119031
rect 519372 113801 519400 123655
rect 519464 117881 519492 128279
rect 519556 120601 519584 131271
rect 519648 123321 519676 134263
rect 519726 132832 519782 132841
rect 519726 132767 519782 132776
rect 519634 123312 519690 123321
rect 519634 123247 519690 123256
rect 519740 121961 519768 132767
rect 519818 129840 519874 129849
rect 519818 129775 519874 129784
rect 519726 121952 519782 121961
rect 519726 121887 519782 121896
rect 519542 120592 519598 120601
rect 519542 120527 519598 120536
rect 519832 119241 519860 129775
rect 519924 124681 519952 135759
rect 520108 127401 520136 138887
rect 520186 137456 520242 137465
rect 520186 137391 520242 137400
rect 520094 127392 520150 127401
rect 520094 127327 520150 127336
rect 520002 126712 520058 126721
rect 520002 126647 520058 126656
rect 519910 124672 519966 124681
rect 519910 124607 519966 124616
rect 519910 122224 519966 122233
rect 519910 122159 519966 122168
rect 519818 119232 519874 119241
rect 519818 119167 519874 119176
rect 519450 117872 519506 117881
rect 519450 117807 519506 117816
rect 519726 117600 519782 117609
rect 519726 117535 519782 117544
rect 519634 116104 519690 116113
rect 519634 116039 519690 116048
rect 519542 114608 519598 114617
rect 519542 114543 519598 114552
rect 519358 113792 519414 113801
rect 519358 113727 519414 113736
rect 519266 109576 519322 109585
rect 519266 109511 519322 109520
rect 117042 106856 117098 106865
rect 117042 106791 117098 106800
rect 519556 105505 519584 114543
rect 519648 106865 519676 116039
rect 519740 108225 519768 117535
rect 519924 112305 519952 122159
rect 520016 116521 520044 126647
rect 520200 126041 520228 137391
rect 520936 134473 520964 146503
rect 521028 139777 521056 152487
rect 521580 151978 521608 158766
rect 521568 151972 521620 151978
rect 521568 151914 521620 151920
rect 521014 139768 521070 139777
rect 521014 139703 521070 139712
rect 520922 134464 520978 134473
rect 520922 134399 520978 134408
rect 520186 126032 520242 126041
rect 520186 125967 520242 125976
rect 520094 125216 520150 125225
rect 520094 125151 520150 125160
rect 520002 116512 520058 116521
rect 520002 116447 520058 116456
rect 520108 115161 520136 125151
rect 520186 120728 520242 120737
rect 520186 120663 520242 120672
rect 520094 115152 520150 115161
rect 520094 115087 520150 115096
rect 519910 112296 519966 112305
rect 519910 112231 519966 112240
rect 520200 110945 520228 120663
rect 521198 113112 521254 113121
rect 521198 113047 521254 113056
rect 520186 110936 520242 110945
rect 520186 110871 520242 110880
rect 521106 110120 521162 110129
rect 521106 110055 521162 110064
rect 521014 108488 521070 108497
rect 521014 108423 521070 108432
rect 519726 108216 519782 108225
rect 519726 108151 519782 108160
rect 520922 106992 520978 107001
rect 520922 106927 520978 106936
rect 519634 106856 519690 106865
rect 519634 106791 519690 106800
rect 519542 105496 519598 105505
rect 519542 105431 519598 105440
rect 520278 105496 520334 105505
rect 520278 105431 520334 105440
rect 116858 102912 116914 102921
rect 116858 102847 116914 102856
rect 116766 101008 116822 101017
rect 116766 100943 116822 100952
rect 519542 99376 519598 99385
rect 519542 99311 519598 99320
rect 116768 96892 116820 96898
rect 116768 96834 116820 96840
rect 116674 95296 116730 95305
rect 116674 95231 116730 95240
rect 116492 93628 116544 93634
rect 116492 93570 116544 93576
rect 116504 93401 116532 93570
rect 116490 93392 116546 93401
rect 116490 93327 116546 93336
rect 116124 92472 116176 92478
rect 116124 92414 116176 92420
rect 116136 91361 116164 92414
rect 116122 91352 116178 91361
rect 116122 91287 116178 91296
rect 116676 87236 116728 87242
rect 116676 87178 116728 87184
rect 116216 86964 116268 86970
rect 116216 86906 116268 86912
rect 116228 85649 116256 86906
rect 116214 85640 116270 85649
rect 116214 85575 116270 85584
rect 115386 81832 115442 81841
rect 115386 81767 115442 81776
rect 116688 78033 116716 87178
rect 116780 79937 116808 96834
rect 519266 94888 519322 94897
rect 519266 94823 519322 94832
rect 116860 91656 116912 91662
rect 116860 91598 116912 91604
rect 116872 87553 116900 91598
rect 519280 87689 519308 94823
rect 519450 91896 519506 91905
rect 519450 91831 519506 91840
rect 519266 87680 519322 87689
rect 519266 87615 519322 87624
rect 116858 87544 116914 87553
rect 116858 87479 116914 87488
rect 519082 85776 519138 85785
rect 519082 85711 519138 85720
rect 116766 79928 116822 79937
rect 116766 79863 116822 79872
rect 519096 79529 519124 85711
rect 519464 84969 519492 91831
rect 519556 91769 519584 99311
rect 520186 97880 520242 97889
rect 520186 97815 520242 97824
rect 520002 96384 520058 96393
rect 520002 96319 520058 96328
rect 519542 91760 519598 91769
rect 519542 91695 519598 91704
rect 519818 90264 519874 90273
rect 519818 90199 519874 90208
rect 519726 88768 519782 88777
rect 519726 88703 519782 88712
rect 519450 84960 519506 84969
rect 519450 84895 519506 84904
rect 519266 84280 519322 84289
rect 519266 84215 519322 84224
rect 519082 79520 519138 79529
rect 519082 79455 519138 79464
rect 519280 78169 519308 84215
rect 519450 82784 519506 82793
rect 519450 82719 519506 82728
rect 519266 78160 519322 78169
rect 519266 78095 519322 78104
rect 116674 78024 116730 78033
rect 116674 77959 116730 77968
rect 519464 76809 519492 82719
rect 519740 82249 519768 88703
rect 519832 83609 519860 90199
rect 520016 89049 520044 96319
rect 520094 93392 520150 93401
rect 520094 93327 520150 93336
rect 520002 89040 520058 89049
rect 520002 88975 520058 88984
rect 520002 87272 520058 87281
rect 520002 87207 520058 87216
rect 519818 83600 519874 83609
rect 519818 83535 519874 83544
rect 519726 82240 519782 82249
rect 519726 82175 519782 82184
rect 519634 81152 519690 81161
rect 519634 81087 519690 81096
rect 519450 76800 519506 76809
rect 519450 76735 519506 76744
rect 519082 76664 519138 76673
rect 519082 76599 519138 76608
rect 116582 74080 116638 74089
rect 116582 74015 116638 74024
rect 116490 72176 116546 72185
rect 116490 72111 116546 72120
rect 116504 71806 116532 72111
rect 113916 71800 113968 71806
rect 113916 71742 113968 71748
rect 116492 71800 116544 71806
rect 116492 71742 116544 71748
rect 113548 64796 113600 64802
rect 113548 64738 113600 64744
rect 113560 64569 113588 64738
rect 113546 64560 113602 64569
rect 113546 64495 113602 64504
rect 112444 62144 112496 62150
rect 112444 62086 112496 62092
rect 111064 46980 111116 46986
rect 111064 46922 111116 46928
rect 109684 4956 109736 4962
rect 109684 4898 109736 4904
rect 109592 4548 109644 4554
rect 109592 4490 109644 4496
rect 109604 2666 109632 4490
rect 32496 2644 32548 2650
rect 32496 2586 32548 2592
rect 98276 2644 98328 2650
rect 109342 2638 109632 2666
rect 98276 2586 98328 2592
rect 29550 2136 29606 2145
rect 2700 746 2728 2108
rect 6012 1737 6040 2108
rect 5998 1728 6054 1737
rect 5998 1663 6054 1672
rect 9324 1601 9352 2108
rect 9310 1592 9366 1601
rect 9310 1527 9366 1536
rect 12636 1426 12664 2108
rect 15948 1494 15976 2108
rect 19352 1873 19380 2108
rect 19338 1864 19394 1873
rect 19338 1799 19394 1808
rect 15936 1488 15988 1494
rect 15936 1430 15988 1436
rect 12624 1420 12676 1426
rect 12624 1362 12676 1368
rect 22664 1290 22692 2108
rect 25990 2094 26096 2122
rect 29302 2094 29550 2122
rect 26068 2009 26096 2094
rect 29550 2071 29606 2080
rect 26054 2000 26110 2009
rect 26054 1935 26110 1944
rect 22652 1284 22704 1290
rect 22652 1226 22704 1232
rect 32508 762 32536 2586
rect 33046 2272 33102 2281
rect 32706 2230 33046 2258
rect 33046 2207 33102 2216
rect 96344 2168 96396 2174
rect 36004 1630 36032 2108
rect 35992 1624 36044 1630
rect 35992 1566 36044 1572
rect 39316 1562 39344 2108
rect 39304 1556 39356 1562
rect 39304 1498 39356 1504
rect 42628 1222 42656 2108
rect 46032 1698 46060 2108
rect 49344 1766 49372 2108
rect 49332 1760 49384 1766
rect 49332 1702 49384 1708
rect 46020 1692 46072 1698
rect 46020 1634 46072 1640
rect 42616 1216 42668 1222
rect 42616 1158 42668 1164
rect 52656 1154 52684 2108
rect 55968 1465 55996 2108
rect 59372 1834 59400 2108
rect 62684 1902 62712 2108
rect 62672 1896 62724 1902
rect 62672 1838 62724 1844
rect 59360 1828 59412 1834
rect 59360 1770 59412 1776
rect 55954 1456 56010 1465
rect 55954 1391 56010 1400
rect 52644 1148 52696 1154
rect 52644 1090 52696 1096
rect 65996 1086 66024 2108
rect 65984 1080 66036 1086
rect 65984 1022 66036 1028
rect 69308 1018 69336 2108
rect 69296 1012 69348 1018
rect 69296 954 69348 960
rect 72712 950 72740 2108
rect 76024 1970 76052 2108
rect 76012 1964 76064 1970
rect 76012 1906 76064 1912
rect 72700 944 72752 950
rect 32692 870 32812 898
rect 72700 886 72752 892
rect 79336 882 79364 2108
rect 82662 2094 82768 2122
rect 82740 2038 82768 2094
rect 82728 2032 82780 2038
rect 82728 1974 82780 1980
rect 32692 762 32720 870
rect 32784 800 32812 870
rect 79324 876 79376 882
rect 79324 818 79376 824
rect 86052 814 86080 2108
rect 89378 2106 89668 2122
rect 96002 2116 96344 2122
rect 96002 2110 96396 2116
rect 89378 2100 89680 2106
rect 89378 2094 89628 2100
rect 89628 2042 89680 2048
rect 92676 1358 92704 2108
rect 96002 2094 96384 2110
rect 92664 1352 92716 1358
rect 92664 1294 92716 1300
rect 86040 808 86092 814
rect 2688 740 2740 746
rect 32508 734 32720 762
rect 2688 682 2740 688
rect 32770 -400 32826 800
rect 98288 800 98316 2586
rect 106030 2378 106228 2394
rect 106030 2372 106240 2378
rect 106030 2366 106188 2372
rect 106188 2314 106240 2320
rect 102968 2304 103020 2310
rect 99406 2242 99696 2258
rect 102718 2252 102968 2258
rect 102718 2246 103020 2252
rect 99406 2236 99708 2242
rect 99406 2230 99656 2236
rect 102718 2230 103008 2246
rect 99656 2178 99708 2184
rect 109696 2145 109724 4898
rect 109868 4888 109920 4894
rect 109868 4830 109920 4836
rect 109776 4820 109828 4826
rect 109776 4762 109828 4768
rect 109682 2136 109738 2145
rect 109682 2071 109738 2080
rect 109788 1970 109816 4762
rect 109880 2009 109908 4830
rect 109960 4208 110012 4214
rect 109960 4150 110012 4156
rect 109866 2000 109922 2009
rect 109776 1964 109828 1970
rect 109866 1935 109922 1944
rect 109776 1906 109828 1912
rect 109972 1737 110000 4150
rect 110052 2984 110104 2990
rect 110052 2926 110104 2932
rect 109958 1728 110014 1737
rect 109958 1663 110014 1672
rect 110064 1494 110092 2926
rect 110420 2916 110472 2922
rect 110420 2858 110472 2864
rect 98644 1488 98696 1494
rect 98644 1430 98696 1436
rect 110052 1488 110104 1494
rect 110052 1430 110104 1436
rect 98656 1193 98684 1430
rect 110432 1426 110460 2858
rect 111076 2038 111104 46922
rect 111156 29028 111208 29034
rect 111156 28970 111208 28976
rect 111064 2032 111116 2038
rect 111064 1974 111116 1980
rect 111168 1766 111196 28970
rect 111248 27668 111300 27674
rect 111248 27610 111300 27616
rect 111156 1760 111208 1766
rect 111156 1702 111208 1708
rect 111260 1698 111288 27610
rect 111340 19372 111392 19378
rect 111340 19314 111392 19320
rect 111352 2281 111380 19314
rect 112456 4554 112484 62086
rect 113928 53145 113956 71742
rect 116306 70272 116362 70281
rect 116306 70207 116362 70216
rect 116320 69086 116348 70207
rect 114100 69080 114152 69086
rect 114100 69022 114152 69028
rect 116308 69080 116360 69086
rect 116308 69022 116360 69028
rect 113914 53136 113970 53145
rect 113914 53071 113970 53080
rect 113824 52488 113876 52494
rect 113824 52430 113876 52436
rect 113640 44192 113692 44198
rect 113640 44134 113692 44140
rect 112536 24880 112588 24886
rect 112536 24822 112588 24828
rect 112444 4548 112496 4554
rect 112444 4490 112496 4496
rect 111338 2272 111394 2281
rect 111338 2207 111394 2216
rect 111248 1692 111300 1698
rect 111248 1634 111300 1640
rect 100760 1420 100812 1426
rect 100760 1362 100812 1368
rect 110420 1420 110472 1426
rect 110420 1362 110472 1368
rect 100772 1329 100800 1362
rect 100758 1320 100814 1329
rect 100758 1255 100814 1264
rect 112548 1222 112576 24822
rect 113652 19009 113680 44134
rect 113732 33176 113784 33182
rect 113732 33118 113784 33124
rect 113638 19000 113694 19009
rect 113638 18935 113694 18944
rect 113548 13864 113600 13870
rect 113548 13806 113600 13812
rect 113560 6914 113588 13806
rect 113640 8288 113692 8294
rect 113640 8230 113692 8236
rect 113652 7721 113680 8230
rect 113638 7712 113694 7721
rect 113638 7647 113694 7656
rect 113560 6886 113680 6914
rect 113652 1290 113680 6886
rect 113744 1834 113772 33118
rect 113732 1828 113784 1834
rect 113732 1770 113784 1776
rect 113836 1358 113864 52430
rect 113916 48340 113968 48346
rect 113916 48282 113968 48288
rect 113824 1352 113876 1358
rect 113824 1294 113876 1300
rect 113640 1284 113692 1290
rect 113640 1226 113692 1232
rect 112536 1216 112588 1222
rect 98642 1184 98698 1193
rect 112536 1158 112588 1164
rect 98642 1119 98698 1128
rect 113928 814 113956 48282
rect 114112 41857 114140 69022
rect 116214 68368 116270 68377
rect 116214 68303 116270 68312
rect 116228 67658 116256 68303
rect 114192 67652 114244 67658
rect 114192 67594 114244 67600
rect 116216 67652 116268 67658
rect 116216 67594 116268 67600
rect 114098 41848 114154 41857
rect 114098 41783 114154 41792
rect 114008 41472 114060 41478
rect 114008 41414 114060 41420
rect 114020 950 114048 41414
rect 114100 38684 114152 38690
rect 114100 38626 114152 38632
rect 114112 1018 114140 38626
rect 114204 30433 114232 67594
rect 116596 64802 116624 74015
rect 519096 71233 519124 76599
rect 519648 75313 519676 81087
rect 520016 80889 520044 87207
rect 520108 86329 520136 93327
rect 520200 90409 520228 97815
rect 520292 97345 520320 105431
rect 520738 102504 520794 102513
rect 520738 102439 520794 102448
rect 520278 97336 520334 97345
rect 520278 97271 520334 97280
rect 520752 94489 520780 102439
rect 520936 98705 520964 106927
rect 521028 100065 521056 108423
rect 521120 101425 521148 110055
rect 521212 104145 521240 113047
rect 521566 111616 521622 111625
rect 521566 111551 521622 111560
rect 521198 104136 521254 104145
rect 521198 104071 521254 104080
rect 521198 104000 521254 104009
rect 521198 103935 521254 103944
rect 521106 101416 521162 101425
rect 521106 101351 521162 101360
rect 521014 100056 521070 100065
rect 521014 99991 521070 100000
rect 520922 98696 520978 98705
rect 520922 98631 520978 98640
rect 521212 95985 521240 103935
rect 521580 102785 521608 111551
rect 521566 102776 521622 102785
rect 521566 102711 521622 102720
rect 521382 101008 521438 101017
rect 521382 100943 521438 100952
rect 521198 95976 521254 95985
rect 521198 95911 521254 95920
rect 520738 94480 520794 94489
rect 520738 94415 520794 94424
rect 521396 93129 521424 100943
rect 521382 93120 521438 93129
rect 521382 93055 521438 93064
rect 520186 90400 520242 90409
rect 520186 90335 520242 90344
rect 520094 86320 520150 86329
rect 520094 86255 520150 86264
rect 520002 80880 520058 80889
rect 520002 80815 520058 80824
rect 520002 79656 520058 79665
rect 520002 79591 520058 79600
rect 519726 78160 519782 78169
rect 519726 78095 519782 78104
rect 519634 75304 519690 75313
rect 519634 75239 519690 75248
rect 519266 73672 519322 73681
rect 519266 73607 519322 73616
rect 519082 71224 519138 71233
rect 519082 71159 519138 71168
rect 519280 68513 519308 73607
rect 519740 72593 519768 78095
rect 519910 75168 519966 75177
rect 519910 75103 519966 75112
rect 519726 72584 519782 72593
rect 519726 72519 519782 72528
rect 519924 69873 519952 75103
rect 520016 73953 520044 79591
rect 520002 73944 520058 73953
rect 520002 73879 520058 73888
rect 520094 72040 520150 72049
rect 520094 71975 520150 71984
rect 519910 69864 519966 69873
rect 519910 69799 519966 69808
rect 519634 69048 519690 69057
rect 519634 68983 519690 68992
rect 519266 68504 519322 68513
rect 519266 68439 519322 68448
rect 117134 66464 117190 66473
rect 117134 66399 117190 66408
rect 116584 64796 116636 64802
rect 116584 64738 116636 64744
rect 115202 64560 115258 64569
rect 115202 64495 115258 64504
rect 114284 37324 114336 37330
rect 114284 37266 114336 37272
rect 114190 30424 114246 30433
rect 114190 30359 114246 30368
rect 114192 22160 114244 22166
rect 114192 22102 114244 22108
rect 114204 1630 114232 22102
rect 114192 1624 114244 1630
rect 114192 1566 114244 1572
rect 114296 1086 114324 37266
rect 114376 34536 114428 34542
rect 114376 34478 114428 34484
rect 114388 1902 114416 34478
rect 114468 31816 114520 31822
rect 114468 31758 114520 31764
rect 114376 1896 114428 1902
rect 114376 1838 114428 1844
rect 114480 1154 114508 31758
rect 115216 8294 115244 64495
rect 116122 62656 116178 62665
rect 116122 62591 116178 62600
rect 116136 62150 116164 62591
rect 116124 62144 116176 62150
rect 116124 62086 116176 62092
rect 116582 60616 116638 60625
rect 116582 60551 116638 60560
rect 116398 53000 116454 53009
rect 116398 52935 116454 52944
rect 116412 52494 116440 52935
rect 116400 52488 116452 52494
rect 116400 52430 116452 52436
rect 115938 49192 115994 49201
rect 115938 49127 115994 49136
rect 115952 48346 115980 49127
rect 115940 48340 115992 48346
rect 115940 48282 115992 48288
rect 116030 47152 116086 47161
rect 116030 47087 116086 47096
rect 116044 46986 116072 47087
rect 116032 46980 116084 46986
rect 116032 46922 116084 46928
rect 115940 41472 115992 41478
rect 115938 41440 115940 41449
rect 115992 41440 115994 41449
rect 115938 41375 115994 41384
rect 115938 39536 115994 39545
rect 115938 39471 115994 39480
rect 115952 38690 115980 39471
rect 115940 38684 115992 38690
rect 115940 38626 115992 38632
rect 116398 37632 116454 37641
rect 116398 37567 116454 37576
rect 116412 37330 116440 37567
rect 116400 37324 116452 37330
rect 116400 37266 116452 37272
rect 115938 35728 115994 35737
rect 115938 35663 115994 35672
rect 115952 34542 115980 35663
rect 115940 34536 115992 34542
rect 115940 34478 115992 34484
rect 116398 33824 116454 33833
rect 116398 33759 116454 33768
rect 116412 33182 116440 33759
rect 116400 33176 116452 33182
rect 116400 33118 116452 33124
rect 115940 31816 115992 31822
rect 115938 31784 115940 31793
rect 115992 31784 115994 31793
rect 115938 31719 115994 31728
rect 116122 29880 116178 29889
rect 116122 29815 116178 29824
rect 116136 29034 116164 29815
rect 116124 29028 116176 29034
rect 116124 28970 116176 28976
rect 116122 27976 116178 27985
rect 116122 27911 116178 27920
rect 116136 27674 116164 27911
rect 116124 27668 116176 27674
rect 116124 27610 116176 27616
rect 116122 26072 116178 26081
rect 116122 26007 116178 26016
rect 116136 24886 116164 26007
rect 116124 24880 116176 24886
rect 116124 24822 116176 24828
rect 115938 22264 115994 22273
rect 115938 22199 115994 22208
rect 115952 22166 115980 22199
rect 115940 22160 115992 22166
rect 115940 22102 115992 22108
rect 116122 20360 116178 20369
rect 116122 20295 116178 20304
rect 116136 19378 116164 20295
rect 116124 19372 116176 19378
rect 116124 19314 116176 19320
rect 116306 18456 116362 18465
rect 116306 18391 116362 18400
rect 116320 16574 116348 18391
rect 116320 16546 116532 16574
rect 116398 16416 116454 16425
rect 116398 16351 116454 16360
rect 116214 14512 116270 14521
rect 116214 14447 116270 14456
rect 116228 13870 116256 14447
rect 116216 13864 116268 13870
rect 116216 13806 116268 13812
rect 115204 8288 115256 8294
rect 115204 8230 115256 8236
rect 116122 4992 116178 5001
rect 116122 4927 116178 4936
rect 116136 4214 116164 4927
rect 116412 4894 116440 16351
rect 116504 4962 116532 16546
rect 116492 4956 116544 4962
rect 116492 4898 116544 4904
rect 116400 4888 116452 4894
rect 116400 4830 116452 4836
rect 116124 4208 116176 4214
rect 116124 4150 116176 4156
rect 116122 3088 116178 3097
rect 116122 3023 116178 3032
rect 114468 1148 114520 1154
rect 114468 1090 114520 1096
rect 114284 1080 114336 1086
rect 114284 1022 114336 1028
rect 114100 1012 114152 1018
rect 114100 954 114152 960
rect 114008 944 114060 950
rect 114008 886 114060 892
rect 113916 808 113968 814
rect 86040 750 86092 756
rect 98274 -400 98330 800
rect 113916 750 113968 756
rect 116136 746 116164 3023
rect 116596 2378 116624 60551
rect 116674 58712 116730 58721
rect 116674 58647 116730 58656
rect 116584 2372 116636 2378
rect 116584 2314 116636 2320
rect 116688 2310 116716 58647
rect 116766 56808 116822 56817
rect 116766 56743 116822 56752
rect 116676 2304 116728 2310
rect 116676 2246 116728 2252
rect 116780 2242 116808 56743
rect 116858 54904 116914 54913
rect 116858 54839 116914 54848
rect 116768 2236 116820 2242
rect 116768 2178 116820 2184
rect 116872 2174 116900 54839
rect 116950 51096 117006 51105
rect 116950 51031 117006 51040
rect 116860 2168 116912 2174
rect 116860 2110 116912 2116
rect 116964 2106 116992 51031
rect 117042 45248 117098 45257
rect 117042 45183 117098 45192
rect 116952 2100 117004 2106
rect 116952 2042 117004 2048
rect 117056 882 117084 45183
rect 117148 44198 117176 66399
rect 519648 64433 519676 68983
rect 520108 67153 520136 71975
rect 520186 70544 520242 70553
rect 520186 70479 520242 70488
rect 520094 67144 520150 67153
rect 520094 67079 520150 67088
rect 520200 65793 520228 70479
rect 520462 67552 520518 67561
rect 520462 67487 520518 67496
rect 520370 66056 520426 66065
rect 520370 65991 520426 66000
rect 520186 65784 520242 65793
rect 520186 65719 520242 65728
rect 519634 64424 519690 64433
rect 519634 64359 519690 64368
rect 520384 61713 520412 65991
rect 520476 63073 520504 67487
rect 520738 64560 520794 64569
rect 520738 64495 520794 64504
rect 520462 63064 520518 63073
rect 520462 62999 520518 63008
rect 520370 61704 520426 61713
rect 520370 61639 520426 61648
rect 520752 60353 520780 64495
rect 521014 62928 521070 62937
rect 521014 62863 521070 62872
rect 520738 60344 520794 60353
rect 520738 60279 520794 60288
rect 520738 59936 520794 59945
rect 520738 59871 520794 59880
rect 520370 56944 520426 56953
rect 520370 56879 520426 56888
rect 520278 55448 520334 55457
rect 520278 55383 520334 55392
rect 519082 53816 519138 53825
rect 519082 53751 519138 53760
rect 519096 50697 519124 53751
rect 519910 52320 519966 52329
rect 519910 52255 519966 52264
rect 519082 50688 519138 50697
rect 519082 50623 519138 50632
rect 519924 49337 519952 52255
rect 520292 52057 520320 55383
rect 520384 53417 520412 56879
rect 520752 56137 520780 59871
rect 521028 58993 521056 62863
rect 521106 61432 521162 61441
rect 521106 61367 521162 61376
rect 521014 58984 521070 58993
rect 521014 58919 521070 58928
rect 521120 57497 521148 61367
rect 521290 58440 521346 58449
rect 521290 58375 521346 58384
rect 521106 57488 521162 57497
rect 521106 57423 521162 57432
rect 520738 56128 520794 56137
rect 520738 56063 520794 56072
rect 521304 54777 521332 58375
rect 521290 54768 521346 54777
rect 521290 54703 521346 54712
rect 520370 53408 520426 53417
rect 520370 53343 520426 53352
rect 520278 52048 520334 52057
rect 520278 51983 520334 51992
rect 520002 50824 520058 50833
rect 520002 50759 520058 50768
rect 519910 49328 519966 49337
rect 519910 49263 519966 49272
rect 520016 47977 520044 50759
rect 520186 49328 520242 49337
rect 520186 49263 520242 49272
rect 520002 47968 520058 47977
rect 520002 47903 520058 47912
rect 519266 47832 519322 47841
rect 519266 47767 519322 47776
rect 519280 45257 519308 47767
rect 520200 46617 520228 49263
rect 520186 46608 520242 46617
rect 520186 46543 520242 46552
rect 519910 46336 519966 46345
rect 519910 46271 519966 46280
rect 519266 45248 519322 45257
rect 519266 45183 519322 45192
rect 519818 44704 519874 44713
rect 519818 44639 519874 44648
rect 117136 44192 117188 44198
rect 117136 44134 117188 44140
rect 117134 43344 117190 43353
rect 117134 43279 117190 43288
rect 117148 4826 117176 43279
rect 519832 42537 519860 44639
rect 519924 43897 519952 46271
rect 519910 43888 519966 43897
rect 519910 43823 519966 43832
rect 520094 43208 520150 43217
rect 520094 43143 520150 43152
rect 519818 42528 519874 42537
rect 519818 42463 519874 42472
rect 520108 41177 520136 43143
rect 520186 41712 520242 41721
rect 520186 41647 520242 41656
rect 520094 41168 520150 41177
rect 520094 41103 520150 41112
rect 519818 40216 519874 40225
rect 519818 40151 519874 40160
rect 519832 38321 519860 40151
rect 520200 39817 520228 41647
rect 520186 39808 520242 39817
rect 520186 39743 520242 39752
rect 520186 38720 520242 38729
rect 520186 38655 520242 38664
rect 519818 38312 519874 38321
rect 519818 38247 519874 38256
rect 520200 36961 520228 38655
rect 521106 37224 521162 37233
rect 521106 37159 521162 37168
rect 520186 36952 520242 36961
rect 520186 36887 520242 36896
rect 521120 36009 521148 37159
rect 521106 36000 521162 36009
rect 521106 35935 521162 35944
rect 520922 35592 520978 35601
rect 520922 35527 520978 35536
rect 520936 34649 520964 35527
rect 520922 34640 520978 34649
rect 520922 34575 520978 34584
rect 520830 34096 520886 34105
rect 520830 34031 520886 34040
rect 520844 33289 520872 34031
rect 520830 33280 520886 33289
rect 520830 33215 520886 33224
rect 521106 32600 521162 32609
rect 521106 32535 521162 32544
rect 521120 31793 521148 32535
rect 521106 31784 521162 31793
rect 521106 31719 521162 31728
rect 521106 31104 521162 31113
rect 521106 31039 521162 31048
rect 521120 30433 521148 31039
rect 521106 30424 521162 30433
rect 521106 30359 521162 30368
rect 521106 29608 521162 29617
rect 521106 29543 521162 29552
rect 521120 28801 521148 29543
rect 521106 28792 521162 28801
rect 521106 28727 521162 28736
rect 117226 24168 117282 24177
rect 117226 24103 117282 24112
rect 117136 4820 117188 4826
rect 117136 4762 117188 4768
rect 117240 1562 117268 24103
rect 521106 20496 521162 20505
rect 521106 20431 521162 20440
rect 521120 19825 521148 20431
rect 521106 19816 521162 19825
rect 521106 19751 521162 19760
rect 521106 15056 521162 15065
rect 521106 14991 521162 15000
rect 521120 14385 521148 14991
rect 521106 14376 521162 14385
rect 521106 14311 521162 14320
rect 521106 13696 521162 13705
rect 521106 13631 521162 13640
rect 521120 12889 521148 13631
rect 521106 12880 521162 12889
rect 521106 12815 521162 12824
rect 519634 12336 519690 12345
rect 519634 12271 519690 12280
rect 519648 11393 519676 12271
rect 519634 11384 519690 11393
rect 519634 11319 519690 11328
rect 521106 10976 521162 10985
rect 521106 10911 521162 10920
rect 521120 9897 521148 10911
rect 521106 9888 521162 9897
rect 521106 9823 521162 9832
rect 521106 9616 521162 9625
rect 521106 9551 521162 9560
rect 521120 8265 521148 9551
rect 520370 8256 520426 8265
rect 520370 8191 520426 8200
rect 521106 8256 521162 8265
rect 521106 8191 521162 8200
rect 520384 6769 520412 8191
rect 521106 6896 521162 6905
rect 521106 6831 521162 6840
rect 520370 6760 520426 6769
rect 520370 6695 520426 6704
rect 521014 5536 521070 5545
rect 521014 5471 521070 5480
rect 521028 3777 521056 5471
rect 521120 5273 521148 6831
rect 521106 5264 521162 5273
rect 521106 5199 521162 5208
rect 521106 4176 521162 4185
rect 521106 4111 521162 4120
rect 521014 3768 521070 3777
rect 521014 3703 521070 3712
rect 520002 2816 520058 2825
rect 520002 2751 520058 2760
rect 143644 2094 143980 2122
rect 193600 2094 193936 2122
rect 243648 2094 243984 2122
rect 293604 2094 293940 2122
rect 343652 2094 343988 2122
rect 393608 2094 393944 2122
rect 443656 2094 443992 2122
rect 117228 1556 117280 1562
rect 117228 1498 117280 1504
rect 143644 1494 143672 2094
rect 163778 1592 163834 1601
rect 163778 1527 163834 1536
rect 143632 1488 143684 1494
rect 143632 1430 143684 1436
rect 117044 876 117096 882
rect 117044 818 117096 824
rect 163792 800 163820 1527
rect 193600 1426 193628 2094
rect 229282 1728 229338 1737
rect 229282 1663 229338 1672
rect 193588 1420 193640 1426
rect 193588 1362 193640 1368
rect 229296 800 229324 1663
rect 243648 1601 243676 2094
rect 293604 1737 293632 2094
rect 293590 1728 293646 1737
rect 293590 1663 293646 1672
rect 243634 1592 243690 1601
rect 243634 1527 243690 1536
rect 343652 1465 343680 2094
rect 393608 1465 393636 2094
rect 443656 1465 443684 2094
rect 493934 1902 493962 2108
rect 491300 1896 491352 1902
rect 491300 1838 491352 1844
rect 493922 1896 493974 1902
rect 493922 1838 493974 1844
rect 294786 1456 294842 1465
rect 294786 1391 294842 1400
rect 343638 1456 343694 1465
rect 343638 1391 343694 1400
rect 360290 1456 360346 1465
rect 360290 1391 360346 1400
rect 393594 1456 393650 1465
rect 393594 1391 393650 1400
rect 425794 1456 425850 1465
rect 425794 1391 425850 1400
rect 443642 1456 443698 1465
rect 443642 1391 443698 1400
rect 294800 800 294828 1391
rect 360304 800 360332 1391
rect 425808 800 425836 1391
rect 491312 800 491340 1838
rect 116124 740 116176 746
rect 116124 682 116176 688
rect 163778 -400 163834 800
rect 229282 -400 229338 800
rect 294786 -400 294842 800
rect 360290 -400 360346 800
rect 425794 -400 425850 800
rect 491298 -400 491354 800
rect 520016 785 520044 2751
rect 521120 2281 521148 4111
rect 521106 2272 521162 2281
rect 521106 2207 521162 2216
rect 520002 776 520058 785
rect 520002 711 520058 720
<< via2 >>
rect 7930 156576 7986 156632
rect 7102 153720 7158 153776
rect 12162 157936 12218 157992
rect 10414 153856 10470 153912
rect 19706 159296 19762 159352
rect 28078 156712 28134 156768
rect 27250 155216 27306 155272
rect 16302 152496 16358 152552
rect 9586 152360 9642 152416
rect 23294 152224 23350 152280
rect 12990 152088 13046 152144
rect 9494 151952 9550 152008
rect 2686 151816 2742 151872
rect 2042 151000 2098 151056
rect 19798 150456 19854 150512
rect 33138 159432 33194 159488
rect 32310 158072 32366 158128
rect 30654 155352 30710 155408
rect 29826 152632 29882 152688
rect 38474 153992 38530 154048
rect 28906 151136 28962 151192
rect 42430 158208 42486 158264
rect 37002 150592 37058 150648
rect 44086 151272 44142 151328
rect 70122 159568 70178 159624
rect 74354 160656 74410 160712
rect 71686 151408 71742 151464
rect 82818 156848 82874 156904
rect 85302 155488 85358 155544
rect 87786 160792 87842 160848
rect 85486 151544 85542 151600
rect 109222 152768 109278 152824
rect 110050 152224 110106 152280
rect 106922 149640 106978 149696
rect 6366 149368 6422 149424
rect 16486 149368 16542 149424
rect 30286 149368 30342 149424
rect 116214 152088 116270 152144
rect 113822 151952 113878 152008
rect 111798 149640 111854 149696
rect 113730 144200 113786 144256
rect 113546 110064 113602 110120
rect 114006 150456 114062 150512
rect 113914 149096 113970 149152
rect 114190 149368 114246 149424
rect 114098 132776 114154 132832
rect 116122 148996 116124 149016
rect 116124 148996 116176 149016
rect 116176 148996 116178 149016
rect 116122 148960 116178 148996
rect 116122 147056 116178 147112
rect 116030 145152 116086 145208
rect 114282 121352 114338 121408
rect 114466 98640 114522 98696
rect 116122 143248 116178 143304
rect 116582 149232 116638 149288
rect 116490 141344 116546 141400
rect 116490 139440 116546 139496
rect 116398 137536 116454 137592
rect 116306 135496 116362 135552
rect 116122 131688 116178 131744
rect 115938 129784 115994 129840
rect 116122 127880 116178 127936
rect 116122 125976 116178 126032
rect 116122 124108 116124 124128
rect 116124 124108 116176 124128
rect 116176 124108 116178 124128
rect 116122 124072 116178 124108
rect 115938 122168 115994 122224
rect 116122 120128 116178 120184
rect 114466 87236 114522 87272
rect 114466 87216 114468 87236
rect 114468 87216 114520 87236
rect 114520 87216 114522 87236
rect 116122 118224 116178 118280
rect 116122 116320 116178 116376
rect 116122 114452 116124 114472
rect 116124 114452 116176 114472
rect 116176 114452 116178 114472
rect 116122 114416 116178 114452
rect 116122 112512 116178 112568
rect 115294 83680 115350 83736
rect 115938 104796 115940 104816
rect 115940 104796 115992 104816
rect 115992 104796 115994 104816
rect 115938 104760 115994 104796
rect 116490 99048 116546 99104
rect 116582 97144 116638 97200
rect 118974 151000 119030 151056
rect 116950 150592 117006 150648
rect 124770 156576 124826 156632
rect 124310 153720 124366 153776
rect 125506 153720 125562 153776
rect 127622 159296 127678 159352
rect 127070 157936 127126 157992
rect 126886 153856 126942 153912
rect 126334 152360 126390 152416
rect 131394 152496 131450 152552
rect 136362 159432 136418 159488
rect 137466 159432 137522 159488
rect 139398 156712 139454 156768
rect 142342 155352 142398 155408
rect 139766 155216 139822 155272
rect 141698 152632 141754 152688
rect 141054 151136 141110 151192
rect 142526 155216 142582 155272
rect 145930 159568 145986 159624
rect 143630 158072 143686 158128
rect 146114 157936 146170 157992
rect 145930 153856 145986 153912
rect 148138 153992 148194 154048
rect 150530 158208 150586 158264
rect 152554 151272 152610 151328
rect 157062 152768 157118 152824
rect 159362 159296 159418 159352
rect 161386 152360 161442 152416
rect 162674 156576 162730 156632
rect 172518 153856 172574 153912
rect 175462 160656 175518 160712
rect 173162 151408 173218 151464
rect 178682 153856 178738 153912
rect 180982 156848 181038 156904
rect 182914 156712 182970 156768
rect 183374 151544 183430 151600
rect 184018 155488 184074 155544
rect 185950 160792 186006 160848
rect 189630 155352 189686 155408
rect 195242 152496 195298 152552
rect 201314 159432 201370 159488
rect 203338 157936 203394 157992
rect 204718 159432 204774 159488
rect 207294 157936 207350 157992
rect 209778 153720 209834 153776
rect 218702 152496 218758 152552
rect 222106 152496 222162 152552
rect 223486 153720 223542 153776
rect 227718 155216 227774 155272
rect 227902 155216 227958 155272
rect 235998 159296 236054 159352
rect 235906 158072 235962 158128
rect 241886 152360 241942 152416
rect 243082 156576 243138 156632
rect 247038 156576 247094 156632
rect 255318 153856 255374 153912
rect 255502 153856 255558 153912
rect 258538 156712 258594 156768
rect 263690 155352 263746 155408
rect 265070 159432 265126 159488
rect 263874 155352 263930 155408
rect 276018 157936 276074 157992
rect 277766 152496 277822 152552
rect 284850 153720 284906 153776
rect 287426 155216 287482 155272
rect 292578 156576 292634 156632
rect 298650 158072 298706 158128
rect 297730 153856 297786 153912
rect 302882 155352 302938 155408
rect 519358 158616 519414 158672
rect 116950 108704 117006 108760
rect 519726 163104 519782 163160
rect 519542 161608 519598 161664
rect 519634 160112 519690 160168
rect 519542 147872 519598 147928
rect 520094 157120 520150 157176
rect 519910 153992 519966 154048
rect 519818 151000 519874 151056
rect 519726 149232 519782 149288
rect 519726 148008 519782 148064
rect 519634 146512 519690 146568
rect 519358 145152 519414 145208
rect 519542 144880 519598 144936
rect 519266 143384 519322 143440
rect 117226 133592 117282 133648
rect 519358 141888 519414 141944
rect 519266 131416 519322 131472
rect 519450 140392 519506 140448
rect 519358 130056 519414 130112
rect 520002 149504 520058 149560
rect 519910 141072 519966 141128
rect 519818 138352 519874 138408
rect 520186 155624 520242 155680
rect 520094 143792 520150 143848
rect 521014 152496 521070 152552
rect 520922 146512 520978 146568
rect 520186 142432 520242 142488
rect 520094 138896 520150 138952
rect 520002 136992 520058 137048
rect 519910 135768 519966 135824
rect 519726 135632 519782 135688
rect 519634 134272 519690 134328
rect 519542 132912 519598 132968
rect 519542 131280 519598 131336
rect 519450 128696 519506 128752
rect 519450 128288 519506 128344
rect 519358 123664 519414 123720
rect 519266 119040 519322 119096
rect 117134 110608 117190 110664
rect 519726 132776 519782 132832
rect 519634 123256 519690 123312
rect 519818 129784 519874 129840
rect 519726 121896 519782 121952
rect 519542 120536 519598 120592
rect 520186 137400 520242 137456
rect 520094 127336 520150 127392
rect 520002 126656 520058 126712
rect 519910 124616 519966 124672
rect 519910 122168 519966 122224
rect 519818 119176 519874 119232
rect 519450 117816 519506 117872
rect 519726 117544 519782 117600
rect 519634 116048 519690 116104
rect 519542 114552 519598 114608
rect 519358 113736 519414 113792
rect 519266 109520 519322 109576
rect 117042 106800 117098 106856
rect 521014 139712 521070 139768
rect 520922 134408 520978 134464
rect 520186 125976 520242 126032
rect 520094 125160 520150 125216
rect 520002 116456 520058 116512
rect 520186 120672 520242 120728
rect 520094 115096 520150 115152
rect 519910 112240 519966 112296
rect 521198 113056 521254 113112
rect 520186 110880 520242 110936
rect 521106 110064 521162 110120
rect 521014 108432 521070 108488
rect 519726 108160 519782 108216
rect 520922 106936 520978 106992
rect 519634 106800 519690 106856
rect 519542 105440 519598 105496
rect 520278 105440 520334 105496
rect 116858 102856 116914 102912
rect 116766 100952 116822 101008
rect 519542 99320 519598 99376
rect 116674 95240 116730 95296
rect 116490 93336 116546 93392
rect 116122 91296 116178 91352
rect 116214 85584 116270 85640
rect 115386 81776 115442 81832
rect 519266 94832 519322 94888
rect 519450 91840 519506 91896
rect 519266 87624 519322 87680
rect 116858 87488 116914 87544
rect 519082 85720 519138 85776
rect 116766 79872 116822 79928
rect 520186 97824 520242 97880
rect 520002 96328 520058 96384
rect 519542 91704 519598 91760
rect 519818 90208 519874 90264
rect 519726 88712 519782 88768
rect 519450 84904 519506 84960
rect 519266 84224 519322 84280
rect 519082 79464 519138 79520
rect 519450 82728 519506 82784
rect 519266 78104 519322 78160
rect 116674 77968 116730 78024
rect 520094 93336 520150 93392
rect 520002 88984 520058 89040
rect 520002 87216 520058 87272
rect 519818 83544 519874 83600
rect 519726 82184 519782 82240
rect 519634 81096 519690 81152
rect 519450 76744 519506 76800
rect 519082 76608 519138 76664
rect 116582 74024 116638 74080
rect 116490 72120 116546 72176
rect 113546 64504 113602 64560
rect 5998 1672 6054 1728
rect 9310 1536 9366 1592
rect 19338 1808 19394 1864
rect 29550 2080 29606 2136
rect 26054 1944 26110 2000
rect 33046 2216 33102 2272
rect 55954 1400 56010 1456
rect 109682 2080 109738 2136
rect 109866 1944 109922 2000
rect 109958 1672 110014 1728
rect 116306 70216 116362 70272
rect 113914 53080 113970 53136
rect 111338 2216 111394 2272
rect 100758 1264 100814 1320
rect 113638 18944 113694 19000
rect 113638 7656 113694 7712
rect 98642 1128 98698 1184
rect 116214 68312 116270 68368
rect 114098 41792 114154 41848
rect 520738 102448 520794 102504
rect 520278 97280 520334 97336
rect 521566 111560 521622 111616
rect 521198 104080 521254 104136
rect 521198 103944 521254 104000
rect 521106 101360 521162 101416
rect 521014 100000 521070 100056
rect 520922 98640 520978 98696
rect 521566 102720 521622 102776
rect 521382 100952 521438 101008
rect 521198 95920 521254 95976
rect 520738 94424 520794 94480
rect 521382 93064 521438 93120
rect 520186 90344 520242 90400
rect 520094 86264 520150 86320
rect 520002 80824 520058 80880
rect 520002 79600 520058 79656
rect 519726 78104 519782 78160
rect 519634 75248 519690 75304
rect 519266 73616 519322 73672
rect 519082 71168 519138 71224
rect 519910 75112 519966 75168
rect 519726 72528 519782 72584
rect 520002 73888 520058 73944
rect 520094 71984 520150 72040
rect 519910 69808 519966 69864
rect 519634 68992 519690 69048
rect 519266 68448 519322 68504
rect 117134 66408 117190 66464
rect 115202 64504 115258 64560
rect 114190 30368 114246 30424
rect 116122 62600 116178 62656
rect 116582 60560 116638 60616
rect 116398 52944 116454 53000
rect 115938 49136 115994 49192
rect 116030 47096 116086 47152
rect 115938 41420 115940 41440
rect 115940 41420 115992 41440
rect 115992 41420 115994 41440
rect 115938 41384 115994 41420
rect 115938 39480 115994 39536
rect 116398 37576 116454 37632
rect 115938 35672 115994 35728
rect 116398 33768 116454 33824
rect 115938 31764 115940 31784
rect 115940 31764 115992 31784
rect 115992 31764 115994 31784
rect 115938 31728 115994 31764
rect 116122 29824 116178 29880
rect 116122 27920 116178 27976
rect 116122 26016 116178 26072
rect 115938 22208 115994 22264
rect 116122 20304 116178 20360
rect 116306 18400 116362 18456
rect 116398 16360 116454 16416
rect 116214 14456 116270 14512
rect 116122 4936 116178 4992
rect 116122 3032 116178 3088
rect 116674 58656 116730 58712
rect 116766 56752 116822 56808
rect 116858 54848 116914 54904
rect 116950 51040 117006 51096
rect 117042 45192 117098 45248
rect 520186 70488 520242 70544
rect 520094 67088 520150 67144
rect 520462 67496 520518 67552
rect 520370 66000 520426 66056
rect 520186 65728 520242 65784
rect 519634 64368 519690 64424
rect 520738 64504 520794 64560
rect 520462 63008 520518 63064
rect 520370 61648 520426 61704
rect 521014 62872 521070 62928
rect 520738 60288 520794 60344
rect 520738 59880 520794 59936
rect 520370 56888 520426 56944
rect 520278 55392 520334 55448
rect 519082 53760 519138 53816
rect 519910 52264 519966 52320
rect 519082 50632 519138 50688
rect 521106 61376 521162 61432
rect 521014 58928 521070 58984
rect 521290 58384 521346 58440
rect 521106 57432 521162 57488
rect 520738 56072 520794 56128
rect 521290 54712 521346 54768
rect 520370 53352 520426 53408
rect 520278 51992 520334 52048
rect 520002 50768 520058 50824
rect 519910 49272 519966 49328
rect 520186 49272 520242 49328
rect 520002 47912 520058 47968
rect 519266 47776 519322 47832
rect 520186 46552 520242 46608
rect 519910 46280 519966 46336
rect 519266 45192 519322 45248
rect 519818 44648 519874 44704
rect 117134 43288 117190 43344
rect 519910 43832 519966 43888
rect 520094 43152 520150 43208
rect 519818 42472 519874 42528
rect 520186 41656 520242 41712
rect 520094 41112 520150 41168
rect 519818 40160 519874 40216
rect 520186 39752 520242 39808
rect 520186 38664 520242 38720
rect 519818 38256 519874 38312
rect 521106 37168 521162 37224
rect 520186 36896 520242 36952
rect 521106 35944 521162 36000
rect 520922 35536 520978 35592
rect 520922 34584 520978 34640
rect 520830 34040 520886 34096
rect 520830 33224 520886 33280
rect 521106 32544 521162 32600
rect 521106 31728 521162 31784
rect 521106 31048 521162 31104
rect 521106 30368 521162 30424
rect 521106 29552 521162 29608
rect 521106 28736 521162 28792
rect 117226 24112 117282 24168
rect 521106 20440 521162 20496
rect 521106 19760 521162 19816
rect 521106 15000 521162 15056
rect 521106 14320 521162 14376
rect 521106 13640 521162 13696
rect 521106 12824 521162 12880
rect 519634 12280 519690 12336
rect 519634 11328 519690 11384
rect 521106 10920 521162 10976
rect 521106 9832 521162 9888
rect 521106 9560 521162 9616
rect 520370 8200 520426 8256
rect 521106 8200 521162 8256
rect 521106 6840 521162 6896
rect 520370 6704 520426 6760
rect 521014 5480 521070 5536
rect 521106 5208 521162 5264
rect 521106 4120 521162 4176
rect 521014 3712 521070 3768
rect 520002 2760 520058 2816
rect 163778 1536 163834 1592
rect 229282 1672 229338 1728
rect 293590 1672 293646 1728
rect 243634 1536 243690 1592
rect 294786 1400 294842 1456
rect 343638 1400 343694 1456
rect 360290 1400 360346 1456
rect 393594 1400 393650 1456
rect 425794 1400 425850 1456
rect 443642 1400 443698 1456
rect 521106 2216 521162 2272
rect 520002 720 520058 776
<< metal3 >>
rect 519721 163162 519787 163165
rect 523200 163162 524400 163192
rect 519721 163160 524400 163162
rect 519721 163104 519726 163160
rect 519782 163104 524400 163160
rect 519721 163102 524400 163104
rect 519721 163099 519787 163102
rect 523200 163072 524400 163102
rect 519537 161666 519603 161669
rect 523200 161666 524400 161696
rect 519537 161664 524400 161666
rect 519537 161608 519542 161664
rect 519598 161608 524400 161664
rect 519537 161606 524400 161608
rect 519537 161603 519603 161606
rect 523200 161576 524400 161606
rect 87781 160850 87847 160853
rect 185945 160850 186011 160853
rect 87781 160848 186011 160850
rect 87781 160792 87786 160848
rect 87842 160792 185950 160848
rect 186006 160792 186011 160848
rect 87781 160790 186011 160792
rect 87781 160787 87847 160790
rect 185945 160787 186011 160790
rect 74349 160714 74415 160717
rect 175457 160714 175523 160717
rect 74349 160712 175523 160714
rect 74349 160656 74354 160712
rect 74410 160656 175462 160712
rect 175518 160656 175523 160712
rect 74349 160654 175523 160656
rect 74349 160651 74415 160654
rect 175457 160651 175523 160654
rect 519629 160170 519695 160173
rect 523200 160170 524400 160200
rect 519629 160168 524400 160170
rect 519629 160112 519634 160168
rect 519690 160112 524400 160168
rect 519629 160110 524400 160112
rect 519629 160107 519695 160110
rect 523200 160080 524400 160110
rect 70117 159626 70183 159629
rect 145925 159626 145991 159629
rect 70117 159624 145991 159626
rect 70117 159568 70122 159624
rect 70178 159568 145930 159624
rect 145986 159568 145991 159624
rect 70117 159566 145991 159568
rect 70117 159563 70183 159566
rect 145925 159563 145991 159566
rect 33133 159490 33199 159493
rect 136357 159490 136423 159493
rect 33133 159488 136423 159490
rect 33133 159432 33138 159488
rect 33194 159432 136362 159488
rect 136418 159432 136423 159488
rect 33133 159430 136423 159432
rect 33133 159427 33199 159430
rect 136357 159427 136423 159430
rect 137461 159490 137527 159493
rect 201309 159490 201375 159493
rect 137461 159488 201375 159490
rect 137461 159432 137466 159488
rect 137522 159432 201314 159488
rect 201370 159432 201375 159488
rect 137461 159430 201375 159432
rect 137461 159427 137527 159430
rect 201309 159427 201375 159430
rect 204713 159490 204779 159493
rect 265065 159490 265131 159493
rect 204713 159488 265131 159490
rect 204713 159432 204718 159488
rect 204774 159432 265070 159488
rect 265126 159432 265131 159488
rect 204713 159430 265131 159432
rect 204713 159427 204779 159430
rect 265065 159427 265131 159430
rect 19701 159354 19767 159357
rect 127617 159354 127683 159357
rect 19701 159352 127683 159354
rect 19701 159296 19706 159352
rect 19762 159296 127622 159352
rect 127678 159296 127683 159352
rect 19701 159294 127683 159296
rect 19701 159291 19767 159294
rect 127617 159291 127683 159294
rect 159357 159354 159423 159357
rect 235993 159354 236059 159357
rect 159357 159352 236059 159354
rect 159357 159296 159362 159352
rect 159418 159296 235998 159352
rect 236054 159296 236059 159352
rect 159357 159294 236059 159296
rect 159357 159291 159423 159294
rect 235993 159291 236059 159294
rect 519353 158674 519419 158677
rect 523200 158674 524400 158704
rect 519353 158672 524400 158674
rect 519353 158616 519358 158672
rect 519414 158616 524400 158672
rect 519353 158614 524400 158616
rect 519353 158611 519419 158614
rect 523200 158584 524400 158614
rect 42425 158266 42491 158269
rect 150525 158266 150591 158269
rect 42425 158264 150591 158266
rect 42425 158208 42430 158264
rect 42486 158208 150530 158264
rect 150586 158208 150591 158264
rect 42425 158206 150591 158208
rect 42425 158203 42491 158206
rect 150525 158203 150591 158206
rect 32305 158130 32371 158133
rect 143625 158130 143691 158133
rect 32305 158128 143691 158130
rect 32305 158072 32310 158128
rect 32366 158072 143630 158128
rect 143686 158072 143691 158128
rect 32305 158070 143691 158072
rect 32305 158067 32371 158070
rect 143625 158067 143691 158070
rect 235901 158130 235967 158133
rect 298645 158130 298711 158133
rect 235901 158128 298711 158130
rect 235901 158072 235906 158128
rect 235962 158072 298650 158128
rect 298706 158072 298711 158128
rect 235901 158070 298711 158072
rect 235901 158067 235967 158070
rect 298645 158067 298711 158070
rect 12157 157994 12223 157997
rect 127065 157994 127131 157997
rect 12157 157992 127131 157994
rect 12157 157936 12162 157992
rect 12218 157936 127070 157992
rect 127126 157936 127131 157992
rect 12157 157934 127131 157936
rect 12157 157931 12223 157934
rect 127065 157931 127131 157934
rect 146109 157994 146175 157997
rect 203333 157994 203399 157997
rect 146109 157992 203399 157994
rect 146109 157936 146114 157992
rect 146170 157936 203338 157992
rect 203394 157936 203399 157992
rect 146109 157934 203399 157936
rect 146109 157931 146175 157934
rect 203333 157931 203399 157934
rect 207289 157994 207355 157997
rect 276013 157994 276079 157997
rect 207289 157992 276079 157994
rect 207289 157936 207294 157992
rect 207350 157936 276018 157992
rect 276074 157936 276079 157992
rect 207289 157934 276079 157936
rect 207289 157931 207355 157934
rect 276013 157931 276079 157934
rect 520089 157178 520155 157181
rect 523200 157178 524400 157208
rect 520089 157176 524400 157178
rect 520089 157120 520094 157176
rect 520150 157120 524400 157176
rect 520089 157118 524400 157120
rect 520089 157115 520155 157118
rect 523200 157088 524400 157118
rect 82813 156906 82879 156909
rect 180977 156906 181043 156909
rect 82813 156904 181043 156906
rect 82813 156848 82818 156904
rect 82874 156848 180982 156904
rect 181038 156848 181043 156904
rect 82813 156846 181043 156848
rect 82813 156843 82879 156846
rect 180977 156843 181043 156846
rect 28073 156770 28139 156773
rect 139393 156770 139459 156773
rect 28073 156768 139459 156770
rect 28073 156712 28078 156768
rect 28134 156712 139398 156768
rect 139454 156712 139459 156768
rect 28073 156710 139459 156712
rect 28073 156707 28139 156710
rect 139393 156707 139459 156710
rect 182909 156770 182975 156773
rect 258533 156770 258599 156773
rect 182909 156768 258599 156770
rect 182909 156712 182914 156768
rect 182970 156712 258538 156768
rect 258594 156712 258599 156768
rect 182909 156710 258599 156712
rect 182909 156707 182975 156710
rect 258533 156707 258599 156710
rect 7925 156634 7991 156637
rect 124765 156634 124831 156637
rect 7925 156632 124831 156634
rect 7925 156576 7930 156632
rect 7986 156576 124770 156632
rect 124826 156576 124831 156632
rect 7925 156574 124831 156576
rect 7925 156571 7991 156574
rect 124765 156571 124831 156574
rect 162669 156634 162735 156637
rect 243077 156634 243143 156637
rect 162669 156632 243143 156634
rect 162669 156576 162674 156632
rect 162730 156576 243082 156632
rect 243138 156576 243143 156632
rect 162669 156574 243143 156576
rect 162669 156571 162735 156574
rect 243077 156571 243143 156574
rect 247033 156634 247099 156637
rect 292573 156634 292639 156637
rect 247033 156632 292639 156634
rect 247033 156576 247038 156632
rect 247094 156576 292578 156632
rect 292634 156576 292639 156632
rect 247033 156574 292639 156576
rect 247033 156571 247099 156574
rect 292573 156571 292639 156574
rect 520181 155682 520247 155685
rect 523200 155682 524400 155712
rect 520181 155680 524400 155682
rect 520181 155624 520186 155680
rect 520242 155624 524400 155680
rect 520181 155622 524400 155624
rect 520181 155619 520247 155622
rect 523200 155592 524400 155622
rect 85297 155546 85363 155549
rect 184013 155546 184079 155549
rect 85297 155544 184079 155546
rect 85297 155488 85302 155544
rect 85358 155488 184018 155544
rect 184074 155488 184079 155544
rect 85297 155486 184079 155488
rect 85297 155483 85363 155486
rect 184013 155483 184079 155486
rect 30649 155410 30715 155413
rect 142337 155410 142403 155413
rect 30649 155408 142403 155410
rect 30649 155352 30654 155408
rect 30710 155352 142342 155408
rect 142398 155352 142403 155408
rect 30649 155350 142403 155352
rect 30649 155347 30715 155350
rect 142337 155347 142403 155350
rect 189625 155410 189691 155413
rect 263685 155410 263751 155413
rect 189625 155408 263751 155410
rect 189625 155352 189630 155408
rect 189686 155352 263690 155408
rect 263746 155352 263751 155408
rect 189625 155350 263751 155352
rect 189625 155347 189691 155350
rect 263685 155347 263751 155350
rect 263869 155410 263935 155413
rect 302877 155410 302943 155413
rect 263869 155408 302943 155410
rect 263869 155352 263874 155408
rect 263930 155352 302882 155408
rect 302938 155352 302943 155408
rect 263869 155350 302943 155352
rect 263869 155347 263935 155350
rect 302877 155347 302943 155350
rect 27245 155274 27311 155277
rect 139761 155274 139827 155277
rect 27245 155272 139827 155274
rect 27245 155216 27250 155272
rect 27306 155216 139766 155272
rect 139822 155216 139827 155272
rect 27245 155214 139827 155216
rect 27245 155211 27311 155214
rect 139761 155211 139827 155214
rect 142521 155274 142587 155277
rect 227713 155274 227779 155277
rect 142521 155272 227779 155274
rect 142521 155216 142526 155272
rect 142582 155216 227718 155272
rect 227774 155216 227779 155272
rect 142521 155214 227779 155216
rect 142521 155211 142587 155214
rect 227713 155211 227779 155214
rect 227897 155274 227963 155277
rect 287421 155274 287487 155277
rect 227897 155272 287487 155274
rect 227897 155216 227902 155272
rect 227958 155216 287426 155272
rect 287482 155216 287487 155272
rect 227897 155214 287487 155216
rect 227897 155211 227963 155214
rect 287421 155211 287487 155214
rect 38469 154050 38535 154053
rect 148133 154050 148199 154053
rect 38469 154048 148199 154050
rect 38469 153992 38474 154048
rect 38530 153992 148138 154048
rect 148194 153992 148199 154048
rect 38469 153990 148199 153992
rect 38469 153987 38535 153990
rect 148133 153987 148199 153990
rect 519905 154050 519971 154053
rect 523200 154050 524400 154080
rect 519905 154048 524400 154050
rect 519905 153992 519910 154048
rect 519966 153992 524400 154048
rect 519905 153990 524400 153992
rect 519905 153987 519971 153990
rect 523200 153960 524400 153990
rect 10409 153914 10475 153917
rect 126881 153914 126947 153917
rect 10409 153912 126947 153914
rect 10409 153856 10414 153912
rect 10470 153856 126886 153912
rect 126942 153856 126947 153912
rect 10409 153854 126947 153856
rect 10409 153851 10475 153854
rect 126881 153851 126947 153854
rect 145925 153914 145991 153917
rect 172513 153914 172579 153917
rect 145925 153912 172579 153914
rect 145925 153856 145930 153912
rect 145986 153856 172518 153912
rect 172574 153856 172579 153912
rect 145925 153854 172579 153856
rect 145925 153851 145991 153854
rect 172513 153851 172579 153854
rect 178677 153914 178743 153917
rect 255313 153914 255379 153917
rect 178677 153912 255379 153914
rect 178677 153856 178682 153912
rect 178738 153856 255318 153912
rect 255374 153856 255379 153912
rect 178677 153854 255379 153856
rect 178677 153851 178743 153854
rect 255313 153851 255379 153854
rect 255497 153914 255563 153917
rect 297725 153914 297791 153917
rect 255497 153912 297791 153914
rect 255497 153856 255502 153912
rect 255558 153856 297730 153912
rect 297786 153856 297791 153912
rect 255497 153854 297791 153856
rect 255497 153851 255563 153854
rect 297725 153851 297791 153854
rect 7097 153778 7163 153781
rect 124305 153778 124371 153781
rect 7097 153776 124371 153778
rect 7097 153720 7102 153776
rect 7158 153720 124310 153776
rect 124366 153720 124371 153776
rect 7097 153718 124371 153720
rect 7097 153715 7163 153718
rect 124305 153715 124371 153718
rect 125501 153778 125567 153781
rect 209773 153778 209839 153781
rect 125501 153776 209839 153778
rect 125501 153720 125506 153776
rect 125562 153720 209778 153776
rect 209834 153720 209839 153776
rect 125501 153718 209839 153720
rect 125501 153715 125567 153718
rect 209773 153715 209839 153718
rect 223481 153778 223547 153781
rect 284845 153778 284911 153781
rect 223481 153776 284911 153778
rect 223481 153720 223486 153776
rect 223542 153720 284850 153776
rect 284906 153720 284911 153776
rect 223481 153718 284911 153720
rect 223481 153715 223547 153718
rect 284845 153715 284911 153718
rect 109217 152826 109283 152829
rect 157057 152826 157123 152829
rect 109217 152824 157123 152826
rect 109217 152768 109222 152824
rect 109278 152768 157062 152824
rect 157118 152768 157123 152824
rect 109217 152766 157123 152768
rect 109217 152763 109283 152766
rect 157057 152763 157123 152766
rect 29821 152690 29887 152693
rect 141693 152690 141759 152693
rect 29821 152688 141759 152690
rect 29821 152632 29826 152688
rect 29882 152632 141698 152688
rect 141754 152632 141759 152688
rect 29821 152630 141759 152632
rect 29821 152627 29887 152630
rect 141693 152627 141759 152630
rect 16297 152554 16363 152557
rect 131389 152554 131455 152557
rect 16297 152552 131455 152554
rect 16297 152496 16302 152552
rect 16358 152496 131394 152552
rect 131450 152496 131455 152552
rect 16297 152494 131455 152496
rect 16297 152491 16363 152494
rect 131389 152491 131455 152494
rect 195237 152554 195303 152557
rect 218697 152554 218763 152557
rect 195237 152552 218763 152554
rect 195237 152496 195242 152552
rect 195298 152496 218702 152552
rect 218758 152496 218763 152552
rect 195237 152494 218763 152496
rect 195237 152491 195303 152494
rect 218697 152491 218763 152494
rect 222101 152554 222167 152557
rect 277761 152554 277827 152557
rect 222101 152552 277827 152554
rect 222101 152496 222106 152552
rect 222162 152496 277766 152552
rect 277822 152496 277827 152552
rect 222101 152494 277827 152496
rect 222101 152491 222167 152494
rect 277761 152491 277827 152494
rect 521009 152554 521075 152557
rect 523200 152554 524400 152584
rect 521009 152552 524400 152554
rect 521009 152496 521014 152552
rect 521070 152496 524400 152552
rect 521009 152494 524400 152496
rect 521009 152491 521075 152494
rect 523200 152464 524400 152494
rect 9581 152418 9647 152421
rect 126329 152418 126395 152421
rect 9581 152416 126395 152418
rect 9581 152360 9586 152416
rect 9642 152360 126334 152416
rect 126390 152360 126395 152416
rect 9581 152358 126395 152360
rect 9581 152355 9647 152358
rect 126329 152355 126395 152358
rect 161381 152418 161447 152421
rect 241881 152418 241947 152421
rect 161381 152416 241947 152418
rect 161381 152360 161386 152416
rect 161442 152360 241886 152416
rect 241942 152360 241947 152416
rect 161381 152358 241947 152360
rect 161381 152355 161447 152358
rect 241881 152355 241947 152358
rect 23289 152282 23355 152285
rect 110045 152282 110111 152285
rect 23289 152280 110111 152282
rect 23289 152224 23294 152280
rect 23350 152224 110050 152280
rect 110106 152224 110111 152280
rect 23289 152222 110111 152224
rect 23289 152219 23355 152222
rect 110045 152219 110111 152222
rect 12985 152146 13051 152149
rect 116209 152146 116275 152149
rect 12985 152144 116275 152146
rect 12985 152088 12990 152144
rect 13046 152088 116214 152144
rect 116270 152088 116275 152144
rect 12985 152086 116275 152088
rect 12985 152083 13051 152086
rect 116209 152083 116275 152086
rect 9489 152010 9555 152013
rect 113817 152010 113883 152013
rect 9489 152008 113883 152010
rect 9489 151952 9494 152008
rect 9550 151952 113822 152008
rect 113878 151952 113883 152008
rect 9489 151950 113883 151952
rect 9489 151947 9555 151950
rect 113817 151947 113883 151950
rect 2681 151874 2747 151877
rect 116526 151874 116532 151876
rect 2681 151872 116532 151874
rect 2681 151816 2686 151872
rect 2742 151816 116532 151872
rect 2681 151814 116532 151816
rect 2681 151811 2747 151814
rect 116526 151812 116532 151814
rect 116596 151812 116602 151876
rect 85481 151602 85547 151605
rect 183369 151602 183435 151605
rect 85481 151600 183435 151602
rect 85481 151544 85486 151600
rect 85542 151544 183374 151600
rect 183430 151544 183435 151600
rect 85481 151542 183435 151544
rect 85481 151539 85547 151542
rect 183369 151539 183435 151542
rect 71681 151466 71747 151469
rect 173157 151466 173223 151469
rect 71681 151464 173223 151466
rect 71681 151408 71686 151464
rect 71742 151408 173162 151464
rect 173218 151408 173223 151464
rect 71681 151406 173223 151408
rect 71681 151403 71747 151406
rect 173157 151403 173223 151406
rect 44081 151330 44147 151333
rect 152549 151330 152615 151333
rect 44081 151328 152615 151330
rect 44081 151272 44086 151328
rect 44142 151272 152554 151328
rect 152610 151272 152615 151328
rect 44081 151270 152615 151272
rect 44081 151267 44147 151270
rect 152549 151267 152615 151270
rect 28901 151194 28967 151197
rect 141049 151194 141115 151197
rect 28901 151192 141115 151194
rect 28901 151136 28906 151192
rect 28962 151136 141054 151192
rect 141110 151136 141115 151192
rect 28901 151134 141115 151136
rect 28901 151131 28967 151134
rect 141049 151131 141115 151134
rect 2037 151058 2103 151061
rect 118969 151058 119035 151061
rect 2037 151056 119035 151058
rect 2037 151000 2042 151056
rect 2098 151000 118974 151056
rect 119030 151000 119035 151056
rect 2037 150998 119035 151000
rect 2037 150995 2103 150998
rect 118969 150995 119035 150998
rect 519813 151058 519879 151061
rect 523200 151058 524400 151088
rect 519813 151056 524400 151058
rect 519813 151000 519818 151056
rect 519874 151000 524400 151056
rect 519813 150998 524400 151000
rect 519813 150995 519879 150998
rect 523200 150968 524400 150998
rect 36997 150650 37063 150653
rect 116945 150650 117011 150653
rect 36997 150648 117011 150650
rect 36997 150592 37002 150648
rect 37058 150592 116950 150648
rect 117006 150592 117011 150648
rect 36997 150590 117011 150592
rect 36997 150587 37063 150590
rect 116945 150587 117011 150590
rect 19793 150514 19859 150517
rect 114001 150514 114067 150517
rect 19793 150512 114067 150514
rect 19793 150456 19798 150512
rect 19854 150456 114006 150512
rect 114062 150456 114067 150512
rect 19793 150454 114067 150456
rect 19793 150451 19859 150454
rect 114001 150451 114067 150454
rect 106917 149698 106983 149701
rect 111793 149698 111859 149701
rect 106917 149696 111859 149698
rect 106917 149640 106922 149696
rect 106978 149640 111798 149696
rect 111854 149640 111859 149696
rect 106917 149638 111859 149640
rect 106917 149635 106983 149638
rect 111793 149635 111859 149638
rect 519997 149562 520063 149565
rect 523200 149562 524400 149592
rect 519997 149560 524400 149562
rect 519997 149504 520002 149560
rect 520058 149504 524400 149560
rect 519997 149502 524400 149504
rect 519997 149499 520063 149502
rect 523200 149472 524400 149502
rect 6361 149426 6427 149429
rect 16481 149426 16547 149429
rect 30281 149426 30347 149429
rect 114185 149426 114251 149429
rect 6361 149424 6930 149426
rect 6361 149368 6366 149424
rect 6422 149368 6930 149424
rect 6361 149366 6930 149368
rect 6361 149363 6427 149366
rect 6870 149154 6930 149366
rect 16481 149424 16590 149426
rect 16481 149368 16486 149424
rect 16542 149368 16590 149424
rect 16481 149363 16590 149368
rect 30281 149424 114251 149426
rect 30281 149368 30286 149424
rect 30342 149368 114190 149424
rect 114246 149368 114251 149424
rect 30281 149366 114251 149368
rect 30281 149363 30347 149366
rect 114185 149363 114251 149366
rect 16530 149290 16590 149363
rect 116577 149290 116643 149293
rect 519721 149290 519787 149293
rect 16530 149288 116643 149290
rect 16530 149232 116582 149288
rect 116638 149232 116643 149288
rect 16530 149230 116643 149232
rect 518788 149288 519787 149290
rect 518788 149232 519726 149288
rect 519782 149232 519787 149288
rect 518788 149230 519787 149232
rect 116577 149227 116643 149230
rect 519721 149227 519787 149230
rect 113909 149154 113975 149157
rect 6870 149152 113975 149154
rect 6870 149096 113914 149152
rect 113970 149096 113975 149152
rect 6870 149094 113975 149096
rect 113909 149091 113975 149094
rect 116117 149018 116183 149021
rect 116117 149016 119140 149018
rect 116117 148960 116122 149016
rect 116178 148960 119140 149016
rect 116117 148958 119140 148960
rect 116117 148955 116183 148958
rect 519721 148066 519787 148069
rect 523200 148066 524400 148096
rect 519721 148064 524400 148066
rect 519721 148008 519726 148064
rect 519782 148008 524400 148064
rect 519721 148006 524400 148008
rect 519721 148003 519787 148006
rect 523200 147976 524400 148006
rect 519537 147930 519603 147933
rect 518788 147928 519603 147930
rect 518788 147872 519542 147928
rect 519598 147872 519603 147928
rect 518788 147870 519603 147872
rect 519537 147867 519603 147870
rect 116117 147114 116183 147117
rect 116117 147112 119140 147114
rect 116117 147056 116122 147112
rect 116178 147056 119140 147112
rect 116117 147054 119140 147056
rect 116117 147051 116183 147054
rect 519629 146570 519695 146573
rect 518788 146568 519695 146570
rect 518788 146512 519634 146568
rect 519690 146512 519695 146568
rect 518788 146510 519695 146512
rect 519629 146507 519695 146510
rect 520917 146570 520983 146573
rect 523200 146570 524400 146600
rect 520917 146568 524400 146570
rect 520917 146512 520922 146568
rect 520978 146512 524400 146568
rect 520917 146510 524400 146512
rect 520917 146507 520983 146510
rect 523200 146480 524400 146510
rect 116025 145210 116091 145213
rect 519353 145210 519419 145213
rect 116025 145208 119140 145210
rect 116025 145152 116030 145208
rect 116086 145152 119140 145208
rect 116025 145150 119140 145152
rect 518788 145208 519419 145210
rect 518788 145152 519358 145208
rect 519414 145152 519419 145208
rect 518788 145150 519419 145152
rect 116025 145147 116091 145150
rect 519353 145147 519419 145150
rect 519537 144938 519603 144941
rect 523200 144938 524400 144968
rect 519537 144936 524400 144938
rect 519537 144880 519542 144936
rect 519598 144880 524400 144936
rect 519537 144878 524400 144880
rect 519537 144875 519603 144878
rect 523200 144848 524400 144878
rect 113725 144258 113791 144261
rect 110860 144256 113791 144258
rect 110860 144200 113730 144256
rect 113786 144200 113791 144256
rect 110860 144198 113791 144200
rect 113725 144195 113791 144198
rect 520089 143850 520155 143853
rect 518788 143848 520155 143850
rect 518788 143792 520094 143848
rect 520150 143792 520155 143848
rect 518788 143790 520155 143792
rect 520089 143787 520155 143790
rect 519261 143442 519327 143445
rect 523200 143442 524400 143472
rect 519261 143440 524400 143442
rect 519261 143384 519266 143440
rect 519322 143384 524400 143440
rect 519261 143382 524400 143384
rect 519261 143379 519327 143382
rect 523200 143352 524400 143382
rect 116117 143306 116183 143309
rect 116117 143304 119140 143306
rect 116117 143248 116122 143304
rect 116178 143248 119140 143304
rect 116117 143246 119140 143248
rect 116117 143243 116183 143246
rect 520181 142490 520247 142493
rect 518788 142488 520247 142490
rect 518788 142432 520186 142488
rect 520242 142432 520247 142488
rect 518788 142430 520247 142432
rect 520181 142427 520247 142430
rect 519353 141946 519419 141949
rect 523200 141946 524400 141976
rect 519353 141944 524400 141946
rect 519353 141888 519358 141944
rect 519414 141888 524400 141944
rect 519353 141886 524400 141888
rect 519353 141883 519419 141886
rect 523200 141856 524400 141886
rect 116485 141402 116551 141405
rect 116485 141400 119140 141402
rect 116485 141344 116490 141400
rect 116546 141344 119140 141400
rect 116485 141342 119140 141344
rect 116485 141339 116551 141342
rect 519905 141130 519971 141133
rect 518788 141128 519971 141130
rect 518788 141072 519910 141128
rect 519966 141072 519971 141128
rect 518788 141070 519971 141072
rect 519905 141067 519971 141070
rect 519445 140450 519511 140453
rect 523200 140450 524400 140480
rect 519445 140448 524400 140450
rect 519445 140392 519450 140448
rect 519506 140392 524400 140448
rect 519445 140390 524400 140392
rect 519445 140387 519511 140390
rect 523200 140360 524400 140390
rect 521009 139770 521075 139773
rect 518788 139768 521075 139770
rect 518788 139712 521014 139768
rect 521070 139712 521075 139768
rect 518788 139710 521075 139712
rect 521009 139707 521075 139710
rect 116485 139498 116551 139501
rect 116485 139496 119140 139498
rect 116485 139440 116490 139496
rect 116546 139440 119140 139496
rect 116485 139438 119140 139440
rect 116485 139435 116551 139438
rect 520089 138954 520155 138957
rect 523200 138954 524400 138984
rect 520089 138952 524400 138954
rect 520089 138896 520094 138952
rect 520150 138896 524400 138952
rect 520089 138894 524400 138896
rect 520089 138891 520155 138894
rect 523200 138864 524400 138894
rect 519813 138410 519879 138413
rect 518788 138408 519879 138410
rect 518788 138352 519818 138408
rect 519874 138352 519879 138408
rect 518788 138350 519879 138352
rect 519813 138347 519879 138350
rect 116393 137594 116459 137597
rect 116393 137592 119140 137594
rect 116393 137536 116398 137592
rect 116454 137536 119140 137592
rect 116393 137534 119140 137536
rect 116393 137531 116459 137534
rect 520181 137458 520247 137461
rect 523200 137458 524400 137488
rect 520181 137456 524400 137458
rect 520181 137400 520186 137456
rect 520242 137400 524400 137456
rect 520181 137398 524400 137400
rect 520181 137395 520247 137398
rect 523200 137368 524400 137398
rect 519997 137050 520063 137053
rect 518788 137048 520063 137050
rect 518788 136992 520002 137048
rect 520058 136992 520063 137048
rect 518788 136990 520063 136992
rect 519997 136987 520063 136990
rect 519905 135826 519971 135829
rect 523200 135826 524400 135856
rect 519905 135824 524400 135826
rect 519905 135768 519910 135824
rect 519966 135768 524400 135824
rect 519905 135766 524400 135768
rect 519905 135763 519971 135766
rect 523200 135736 524400 135766
rect 519721 135690 519787 135693
rect 518788 135688 519787 135690
rect 518788 135632 519726 135688
rect 519782 135632 519787 135688
rect 518788 135630 519787 135632
rect 519721 135627 519787 135630
rect 116301 135554 116367 135557
rect 116301 135552 119140 135554
rect 116301 135496 116306 135552
rect 116362 135496 119140 135552
rect 116301 135494 119140 135496
rect 116301 135491 116367 135494
rect 520917 134466 520983 134469
rect 518758 134464 520983 134466
rect 518758 134408 520922 134464
rect 520978 134408 520983 134464
rect 518758 134406 520983 134408
rect 518758 134300 518818 134406
rect 520917 134403 520983 134406
rect 519629 134330 519695 134333
rect 523200 134330 524400 134360
rect 519629 134328 524400 134330
rect 519629 134272 519634 134328
rect 519690 134272 524400 134328
rect 519629 134270 524400 134272
rect 519629 134267 519695 134270
rect 523200 134240 524400 134270
rect 117221 133650 117287 133653
rect 117221 133648 119140 133650
rect 117221 133592 117226 133648
rect 117282 133592 119140 133648
rect 117221 133590 119140 133592
rect 117221 133587 117287 133590
rect 519537 132970 519603 132973
rect 518788 132968 519603 132970
rect 518788 132912 519542 132968
rect 519598 132912 519603 132968
rect 518788 132910 519603 132912
rect 519537 132907 519603 132910
rect 114093 132834 114159 132837
rect 110860 132832 114159 132834
rect 110860 132776 114098 132832
rect 114154 132776 114159 132832
rect 110860 132774 114159 132776
rect 114093 132771 114159 132774
rect 519721 132834 519787 132837
rect 523200 132834 524400 132864
rect 519721 132832 524400 132834
rect 519721 132776 519726 132832
rect 519782 132776 524400 132832
rect 519721 132774 524400 132776
rect 519721 132771 519787 132774
rect 523200 132744 524400 132774
rect 116117 131746 116183 131749
rect 116117 131744 119140 131746
rect 116117 131688 116122 131744
rect 116178 131688 119140 131744
rect 116117 131686 119140 131688
rect 116117 131683 116183 131686
rect 519261 131474 519327 131477
rect 518788 131472 519327 131474
rect 518788 131416 519266 131472
rect 519322 131416 519327 131472
rect 518788 131414 519327 131416
rect 519261 131411 519327 131414
rect 519537 131338 519603 131341
rect 523200 131338 524400 131368
rect 519537 131336 524400 131338
rect 519537 131280 519542 131336
rect 519598 131280 524400 131336
rect 519537 131278 524400 131280
rect 519537 131275 519603 131278
rect 523200 131248 524400 131278
rect 519353 130114 519419 130117
rect 518788 130112 519419 130114
rect 518788 130056 519358 130112
rect 519414 130056 519419 130112
rect 518788 130054 519419 130056
rect 519353 130051 519419 130054
rect 115933 129842 115999 129845
rect 519813 129842 519879 129845
rect 523200 129842 524400 129872
rect 115933 129840 119140 129842
rect 115933 129784 115938 129840
rect 115994 129784 119140 129840
rect 115933 129782 119140 129784
rect 519813 129840 524400 129842
rect 519813 129784 519818 129840
rect 519874 129784 524400 129840
rect 519813 129782 524400 129784
rect 115933 129779 115999 129782
rect 519813 129779 519879 129782
rect 523200 129752 524400 129782
rect 519445 128754 519511 128757
rect 518788 128752 519511 128754
rect 518788 128696 519450 128752
rect 519506 128696 519511 128752
rect 518788 128694 519511 128696
rect 519445 128691 519511 128694
rect 519445 128346 519511 128349
rect 523200 128346 524400 128376
rect 519445 128344 524400 128346
rect 519445 128288 519450 128344
rect 519506 128288 524400 128344
rect 519445 128286 524400 128288
rect 519445 128283 519511 128286
rect 523200 128256 524400 128286
rect 116117 127938 116183 127941
rect 116117 127936 119140 127938
rect 116117 127880 116122 127936
rect 116178 127880 119140 127936
rect 116117 127878 119140 127880
rect 116117 127875 116183 127878
rect 520089 127394 520155 127397
rect 518788 127392 520155 127394
rect 518788 127336 520094 127392
rect 520150 127336 520155 127392
rect 518788 127334 520155 127336
rect 520089 127331 520155 127334
rect 519997 126714 520063 126717
rect 523200 126714 524400 126744
rect 519997 126712 524400 126714
rect 519997 126656 520002 126712
rect 520058 126656 524400 126712
rect 519997 126654 524400 126656
rect 519997 126651 520063 126654
rect 523200 126624 524400 126654
rect 116117 126034 116183 126037
rect 520181 126034 520247 126037
rect 116117 126032 119140 126034
rect 116117 125976 116122 126032
rect 116178 125976 119140 126032
rect 116117 125974 119140 125976
rect 518788 126032 520247 126034
rect 518788 125976 520186 126032
rect 520242 125976 520247 126032
rect 518788 125974 520247 125976
rect 116117 125971 116183 125974
rect 520181 125971 520247 125974
rect 520089 125218 520155 125221
rect 523200 125218 524400 125248
rect 520089 125216 524400 125218
rect 520089 125160 520094 125216
rect 520150 125160 524400 125216
rect 520089 125158 524400 125160
rect 520089 125155 520155 125158
rect 523200 125128 524400 125158
rect 519905 124674 519971 124677
rect 518788 124672 519971 124674
rect 518788 124616 519910 124672
rect 519966 124616 519971 124672
rect 518788 124614 519971 124616
rect 519905 124611 519971 124614
rect 116117 124130 116183 124133
rect 116117 124128 119140 124130
rect 116117 124072 116122 124128
rect 116178 124072 119140 124128
rect 116117 124070 119140 124072
rect 116117 124067 116183 124070
rect 519353 123722 519419 123725
rect 523200 123722 524400 123752
rect 519353 123720 524400 123722
rect 519353 123664 519358 123720
rect 519414 123664 524400 123720
rect 519353 123662 524400 123664
rect 519353 123659 519419 123662
rect 523200 123632 524400 123662
rect 519629 123314 519695 123317
rect 518788 123312 519695 123314
rect 518788 123256 519634 123312
rect 519690 123256 519695 123312
rect 518788 123254 519695 123256
rect 519629 123251 519695 123254
rect 115933 122226 115999 122229
rect 519905 122226 519971 122229
rect 523200 122226 524400 122256
rect 115933 122224 119140 122226
rect 115933 122168 115938 122224
rect 115994 122168 119140 122224
rect 115933 122166 119140 122168
rect 519905 122224 524400 122226
rect 519905 122168 519910 122224
rect 519966 122168 524400 122224
rect 519905 122166 524400 122168
rect 115933 122163 115999 122166
rect 519905 122163 519971 122166
rect 523200 122136 524400 122166
rect 519721 121954 519787 121957
rect 518788 121952 519787 121954
rect 518788 121896 519726 121952
rect 519782 121896 519787 121952
rect 518788 121894 519787 121896
rect 519721 121891 519787 121894
rect 114277 121410 114343 121413
rect 110860 121408 114343 121410
rect 110860 121352 114282 121408
rect 114338 121352 114343 121408
rect 110860 121350 114343 121352
rect 114277 121347 114343 121350
rect 520181 120730 520247 120733
rect 523200 120730 524400 120760
rect 520181 120728 524400 120730
rect 520181 120672 520186 120728
rect 520242 120672 524400 120728
rect 520181 120670 524400 120672
rect 520181 120667 520247 120670
rect 523200 120640 524400 120670
rect 519537 120594 519603 120597
rect 518788 120592 519603 120594
rect 518788 120536 519542 120592
rect 519598 120536 519603 120592
rect 518788 120534 519603 120536
rect 519537 120531 519603 120534
rect 116117 120186 116183 120189
rect 116117 120184 119140 120186
rect 116117 120128 116122 120184
rect 116178 120128 119140 120184
rect 116117 120126 119140 120128
rect 116117 120123 116183 120126
rect 519813 119234 519879 119237
rect 523200 119234 524400 119264
rect 518788 119232 519879 119234
rect 518788 119176 519818 119232
rect 519874 119176 519879 119232
rect 518788 119174 519879 119176
rect 519813 119171 519879 119174
rect 520046 119174 524400 119234
rect 519261 119098 519327 119101
rect 520046 119098 520106 119174
rect 523200 119144 524400 119174
rect 519261 119096 520106 119098
rect 519261 119040 519266 119096
rect 519322 119040 520106 119096
rect 519261 119038 520106 119040
rect 519261 119035 519327 119038
rect 116117 118282 116183 118285
rect 116117 118280 119140 118282
rect 116117 118224 116122 118280
rect 116178 118224 119140 118280
rect 116117 118222 119140 118224
rect 116117 118219 116183 118222
rect 519445 117874 519511 117877
rect 518788 117872 519511 117874
rect 518788 117816 519450 117872
rect 519506 117816 519511 117872
rect 518788 117814 519511 117816
rect 519445 117811 519511 117814
rect 519721 117602 519787 117605
rect 523200 117602 524400 117632
rect 519721 117600 524400 117602
rect 519721 117544 519726 117600
rect 519782 117544 524400 117600
rect 519721 117542 524400 117544
rect 519721 117539 519787 117542
rect 523200 117512 524400 117542
rect 519997 116514 520063 116517
rect 518788 116512 520063 116514
rect 518788 116456 520002 116512
rect 520058 116456 520063 116512
rect 518788 116454 520063 116456
rect 519997 116451 520063 116454
rect 116117 116378 116183 116381
rect 116117 116376 119140 116378
rect 116117 116320 116122 116376
rect 116178 116320 119140 116376
rect 116117 116318 119140 116320
rect 116117 116315 116183 116318
rect 519629 116106 519695 116109
rect 523200 116106 524400 116136
rect 519629 116104 524400 116106
rect 519629 116048 519634 116104
rect 519690 116048 524400 116104
rect 519629 116046 524400 116048
rect 519629 116043 519695 116046
rect 523200 116016 524400 116046
rect 520089 115154 520155 115157
rect 518788 115152 520155 115154
rect 518788 115096 520094 115152
rect 520150 115096 520155 115152
rect 518788 115094 520155 115096
rect 520089 115091 520155 115094
rect 519537 114610 519603 114613
rect 523200 114610 524400 114640
rect 519537 114608 524400 114610
rect 519537 114552 519542 114608
rect 519598 114552 524400 114608
rect 519537 114550 524400 114552
rect 519537 114547 519603 114550
rect 523200 114520 524400 114550
rect 116117 114474 116183 114477
rect 116117 114472 119140 114474
rect 116117 114416 116122 114472
rect 116178 114416 119140 114472
rect 116117 114414 119140 114416
rect 116117 114411 116183 114414
rect 519353 113794 519419 113797
rect 518788 113792 519419 113794
rect 518788 113736 519358 113792
rect 519414 113736 519419 113792
rect 518788 113734 519419 113736
rect 519353 113731 519419 113734
rect 521193 113114 521259 113117
rect 523200 113114 524400 113144
rect 521193 113112 524400 113114
rect 521193 113056 521198 113112
rect 521254 113056 524400 113112
rect 521193 113054 524400 113056
rect 521193 113051 521259 113054
rect 523200 113024 524400 113054
rect 116117 112570 116183 112573
rect 116117 112568 119140 112570
rect 116117 112512 116122 112568
rect 116178 112512 119140 112568
rect 116117 112510 119140 112512
rect 116117 112507 116183 112510
rect 519905 112298 519971 112301
rect 518788 112296 519971 112298
rect 518788 112240 519910 112296
rect 519966 112240 519971 112296
rect 518788 112238 519971 112240
rect 519905 112235 519971 112238
rect 521561 111618 521627 111621
rect 523200 111618 524400 111648
rect 521561 111616 524400 111618
rect 521561 111560 521566 111616
rect 521622 111560 524400 111616
rect 521561 111558 524400 111560
rect 521561 111555 521627 111558
rect 523200 111528 524400 111558
rect 520181 110938 520247 110941
rect 518788 110936 520247 110938
rect 518788 110880 520186 110936
rect 520242 110880 520247 110936
rect 518788 110878 520247 110880
rect 520181 110875 520247 110878
rect 117129 110666 117195 110669
rect 117129 110664 119140 110666
rect 117129 110608 117134 110664
rect 117190 110608 119140 110664
rect 117129 110606 119140 110608
rect 117129 110603 117195 110606
rect 113541 110122 113607 110125
rect 110860 110120 113607 110122
rect 110860 110064 113546 110120
rect 113602 110064 113607 110120
rect 110860 110062 113607 110064
rect 113541 110059 113607 110062
rect 521101 110122 521167 110125
rect 523200 110122 524400 110152
rect 521101 110120 524400 110122
rect 521101 110064 521106 110120
rect 521162 110064 524400 110120
rect 521101 110062 524400 110064
rect 521101 110059 521167 110062
rect 523200 110032 524400 110062
rect 519261 109578 519327 109581
rect 518788 109576 519327 109578
rect 518788 109520 519266 109576
rect 519322 109520 519327 109576
rect 518788 109518 519327 109520
rect 519261 109515 519327 109518
rect 116945 108762 117011 108765
rect 116945 108760 119140 108762
rect 116945 108704 116950 108760
rect 117006 108704 119140 108760
rect 116945 108702 119140 108704
rect 116945 108699 117011 108702
rect 521009 108490 521075 108493
rect 523200 108490 524400 108520
rect 521009 108488 524400 108490
rect 521009 108432 521014 108488
rect 521070 108432 524400 108488
rect 521009 108430 524400 108432
rect 521009 108427 521075 108430
rect 523200 108400 524400 108430
rect 519721 108218 519787 108221
rect 518788 108216 519787 108218
rect 518788 108160 519726 108216
rect 519782 108160 519787 108216
rect 518788 108158 519787 108160
rect 519721 108155 519787 108158
rect 520917 106994 520983 106997
rect 523200 106994 524400 107024
rect 520917 106992 524400 106994
rect 520917 106936 520922 106992
rect 520978 106936 524400 106992
rect 520917 106934 524400 106936
rect 520917 106931 520983 106934
rect 523200 106904 524400 106934
rect 117037 106858 117103 106861
rect 519629 106858 519695 106861
rect 117037 106856 119140 106858
rect 117037 106800 117042 106856
rect 117098 106800 119140 106856
rect 117037 106798 119140 106800
rect 518788 106856 519695 106858
rect 518788 106800 519634 106856
rect 519690 106800 519695 106856
rect 518788 106798 519695 106800
rect 117037 106795 117103 106798
rect 519629 106795 519695 106798
rect 519537 105498 519603 105501
rect 518788 105496 519603 105498
rect 518788 105440 519542 105496
rect 519598 105440 519603 105496
rect 518788 105438 519603 105440
rect 519537 105435 519603 105438
rect 520273 105498 520339 105501
rect 523200 105498 524400 105528
rect 520273 105496 524400 105498
rect 520273 105440 520278 105496
rect 520334 105440 524400 105496
rect 520273 105438 524400 105440
rect 520273 105435 520339 105438
rect 523200 105408 524400 105438
rect 115933 104818 115999 104821
rect 115933 104816 119140 104818
rect 115933 104760 115938 104816
rect 115994 104760 119140 104816
rect 115933 104758 119140 104760
rect 115933 104755 115999 104758
rect 521193 104138 521259 104141
rect 518788 104136 521259 104138
rect 518788 104080 521198 104136
rect 521254 104080 521259 104136
rect 518788 104078 521259 104080
rect 521193 104075 521259 104078
rect 521193 104002 521259 104005
rect 523200 104002 524400 104032
rect 521193 104000 524400 104002
rect 521193 103944 521198 104000
rect 521254 103944 524400 104000
rect 521193 103942 524400 103944
rect 521193 103939 521259 103942
rect 523200 103912 524400 103942
rect 116853 102914 116919 102917
rect 116853 102912 119140 102914
rect 116853 102856 116858 102912
rect 116914 102856 119140 102912
rect 116853 102854 119140 102856
rect 116853 102851 116919 102854
rect 521561 102778 521627 102781
rect 518788 102776 521627 102778
rect 518788 102720 521566 102776
rect 521622 102720 521627 102776
rect 518788 102718 521627 102720
rect 521561 102715 521627 102718
rect 520733 102506 520799 102509
rect 523200 102506 524400 102536
rect 520733 102504 524400 102506
rect 520733 102448 520738 102504
rect 520794 102448 524400 102504
rect 520733 102446 524400 102448
rect 520733 102443 520799 102446
rect 523200 102416 524400 102446
rect 521101 101418 521167 101421
rect 518788 101416 521167 101418
rect 518788 101360 521106 101416
rect 521162 101360 521167 101416
rect 518788 101358 521167 101360
rect 521101 101355 521167 101358
rect 116761 101010 116827 101013
rect 521377 101010 521443 101013
rect 523200 101010 524400 101040
rect 116761 101008 119140 101010
rect 116761 100952 116766 101008
rect 116822 100952 119140 101008
rect 116761 100950 119140 100952
rect 521377 101008 524400 101010
rect 521377 100952 521382 101008
rect 521438 100952 524400 101008
rect 521377 100950 524400 100952
rect 116761 100947 116827 100950
rect 521377 100947 521443 100950
rect 523200 100920 524400 100950
rect 521009 100058 521075 100061
rect 518788 100056 521075 100058
rect 518788 100000 521014 100056
rect 521070 100000 521075 100056
rect 518788 99998 521075 100000
rect 521009 99995 521075 99998
rect 519537 99378 519603 99381
rect 523200 99378 524400 99408
rect 519537 99376 524400 99378
rect 519537 99320 519542 99376
rect 519598 99320 524400 99376
rect 519537 99318 524400 99320
rect 519537 99315 519603 99318
rect 523200 99288 524400 99318
rect 116485 99106 116551 99109
rect 116485 99104 119140 99106
rect 116485 99048 116490 99104
rect 116546 99048 119140 99104
rect 116485 99046 119140 99048
rect 116485 99043 116551 99046
rect 114461 98698 114527 98701
rect 520917 98698 520983 98701
rect 110860 98696 114527 98698
rect 110860 98640 114466 98696
rect 114522 98640 114527 98696
rect 110860 98638 114527 98640
rect 518788 98696 520983 98698
rect 518788 98640 520922 98696
rect 520978 98640 520983 98696
rect 518788 98638 520983 98640
rect 114461 98635 114527 98638
rect 520917 98635 520983 98638
rect 520181 97882 520247 97885
rect 523200 97882 524400 97912
rect 520181 97880 524400 97882
rect 520181 97824 520186 97880
rect 520242 97824 524400 97880
rect 520181 97822 524400 97824
rect 520181 97819 520247 97822
rect 523200 97792 524400 97822
rect 520273 97338 520339 97341
rect 518788 97336 520339 97338
rect 518788 97280 520278 97336
rect 520334 97280 520339 97336
rect 518788 97278 520339 97280
rect 520273 97275 520339 97278
rect 116577 97202 116643 97205
rect 116577 97200 119140 97202
rect 116577 97144 116582 97200
rect 116638 97144 119140 97200
rect 116577 97142 119140 97144
rect 116577 97139 116643 97142
rect 519997 96386 520063 96389
rect 523200 96386 524400 96416
rect 519997 96384 524400 96386
rect 519997 96328 520002 96384
rect 520058 96328 524400 96384
rect 519997 96326 524400 96328
rect 519997 96323 520063 96326
rect 523200 96296 524400 96326
rect 521193 95978 521259 95981
rect 518788 95976 521259 95978
rect 518788 95920 521198 95976
rect 521254 95920 521259 95976
rect 518788 95918 521259 95920
rect 521193 95915 521259 95918
rect 116669 95298 116735 95301
rect 116669 95296 119140 95298
rect 116669 95240 116674 95296
rect 116730 95240 119140 95296
rect 116669 95238 119140 95240
rect 116669 95235 116735 95238
rect 519261 94890 519327 94893
rect 523200 94890 524400 94920
rect 519261 94888 524400 94890
rect 519261 94832 519266 94888
rect 519322 94832 524400 94888
rect 519261 94830 524400 94832
rect 519261 94827 519327 94830
rect 523200 94800 524400 94830
rect 520733 94482 520799 94485
rect 518788 94480 520799 94482
rect 518788 94424 520738 94480
rect 520794 94424 520799 94480
rect 518788 94422 520799 94424
rect 520733 94419 520799 94422
rect 116485 93394 116551 93397
rect 520089 93394 520155 93397
rect 523200 93394 524400 93424
rect 116485 93392 119140 93394
rect 116485 93336 116490 93392
rect 116546 93336 119140 93392
rect 116485 93334 119140 93336
rect 520089 93392 524400 93394
rect 520089 93336 520094 93392
rect 520150 93336 524400 93392
rect 520089 93334 524400 93336
rect 116485 93331 116551 93334
rect 520089 93331 520155 93334
rect 523200 93304 524400 93334
rect 521377 93122 521443 93125
rect 518788 93120 521443 93122
rect 518788 93064 521382 93120
rect 521438 93064 521443 93120
rect 518788 93062 521443 93064
rect 521377 93059 521443 93062
rect 519445 91898 519511 91901
rect 523200 91898 524400 91928
rect 519445 91896 524400 91898
rect 519445 91840 519450 91896
rect 519506 91840 524400 91896
rect 519445 91838 524400 91840
rect 519445 91835 519511 91838
rect 523200 91808 524400 91838
rect 519537 91762 519603 91765
rect 518788 91760 519603 91762
rect 518788 91704 519542 91760
rect 519598 91704 519603 91760
rect 518788 91702 519603 91704
rect 519537 91699 519603 91702
rect 116117 91354 116183 91357
rect 116117 91352 119140 91354
rect 116117 91296 116122 91352
rect 116178 91296 119140 91352
rect 116117 91294 119140 91296
rect 116117 91291 116183 91294
rect 520181 90402 520247 90405
rect 518788 90400 520247 90402
rect 518788 90344 520186 90400
rect 520242 90344 520247 90400
rect 518788 90342 520247 90344
rect 520181 90339 520247 90342
rect 519813 90266 519879 90269
rect 523200 90266 524400 90296
rect 519813 90264 524400 90266
rect 519813 90208 519818 90264
rect 519874 90208 524400 90264
rect 519813 90206 524400 90208
rect 519813 90203 519879 90206
rect 523200 90176 524400 90206
rect 116526 89388 116532 89452
rect 116596 89450 116602 89452
rect 116596 89390 119140 89450
rect 116596 89388 116602 89390
rect 519997 89042 520063 89045
rect 518788 89040 520063 89042
rect 518788 88984 520002 89040
rect 520058 88984 520063 89040
rect 518788 88982 520063 88984
rect 519997 88979 520063 88982
rect 519721 88770 519787 88773
rect 523200 88770 524400 88800
rect 519721 88768 524400 88770
rect 519721 88712 519726 88768
rect 519782 88712 524400 88768
rect 519721 88710 524400 88712
rect 519721 88707 519787 88710
rect 523200 88680 524400 88710
rect 519261 87682 519327 87685
rect 518788 87680 519327 87682
rect 518788 87624 519266 87680
rect 519322 87624 519327 87680
rect 518788 87622 519327 87624
rect 519261 87619 519327 87622
rect 116853 87546 116919 87549
rect 116853 87544 119140 87546
rect 116853 87488 116858 87544
rect 116914 87488 119140 87544
rect 116853 87486 119140 87488
rect 116853 87483 116919 87486
rect 114461 87274 114527 87277
rect 110860 87272 114527 87274
rect 110860 87216 114466 87272
rect 114522 87216 114527 87272
rect 110860 87214 114527 87216
rect 114461 87211 114527 87214
rect 519997 87274 520063 87277
rect 523200 87274 524400 87304
rect 519997 87272 524400 87274
rect 519997 87216 520002 87272
rect 520058 87216 524400 87272
rect 519997 87214 524400 87216
rect 519997 87211 520063 87214
rect 523200 87184 524400 87214
rect 520089 86322 520155 86325
rect 518788 86320 520155 86322
rect 518788 86264 520094 86320
rect 520150 86264 520155 86320
rect 518788 86262 520155 86264
rect 520089 86259 520155 86262
rect 519077 85778 519143 85781
rect 523200 85778 524400 85808
rect 519077 85776 524400 85778
rect 519077 85720 519082 85776
rect 519138 85720 524400 85776
rect 519077 85718 524400 85720
rect 519077 85715 519143 85718
rect 523200 85688 524400 85718
rect 116209 85642 116275 85645
rect 116209 85640 119140 85642
rect 116209 85584 116214 85640
rect 116270 85584 119140 85640
rect 116209 85582 119140 85584
rect 116209 85579 116275 85582
rect 519445 84962 519511 84965
rect 518788 84960 519511 84962
rect 518788 84904 519450 84960
rect 519506 84904 519511 84960
rect 518788 84902 519511 84904
rect 519445 84899 519511 84902
rect 519261 84282 519327 84285
rect 523200 84282 524400 84312
rect 519261 84280 524400 84282
rect 519261 84224 519266 84280
rect 519322 84224 524400 84280
rect 519261 84222 524400 84224
rect 519261 84219 519327 84222
rect 523200 84192 524400 84222
rect 115289 83738 115355 83741
rect 115289 83736 119140 83738
rect 115289 83680 115294 83736
rect 115350 83680 119140 83736
rect 115289 83678 119140 83680
rect 115289 83675 115355 83678
rect 519813 83602 519879 83605
rect 518788 83600 519879 83602
rect 518788 83544 519818 83600
rect 519874 83544 519879 83600
rect 518788 83542 519879 83544
rect 519813 83539 519879 83542
rect 519445 82786 519511 82789
rect 523200 82786 524400 82816
rect 519445 82784 524400 82786
rect 519445 82728 519450 82784
rect 519506 82728 524400 82784
rect 519445 82726 524400 82728
rect 519445 82723 519511 82726
rect 523200 82696 524400 82726
rect 519721 82242 519787 82245
rect 518788 82240 519787 82242
rect 518788 82184 519726 82240
rect 519782 82184 519787 82240
rect 518788 82182 519787 82184
rect 519721 82179 519787 82182
rect 115381 81834 115447 81837
rect 115381 81832 119140 81834
rect 115381 81776 115386 81832
rect 115442 81776 119140 81832
rect 115381 81774 119140 81776
rect 115381 81771 115447 81774
rect 519629 81154 519695 81157
rect 523200 81154 524400 81184
rect 519629 81152 524400 81154
rect 519629 81096 519634 81152
rect 519690 81096 524400 81152
rect 519629 81094 524400 81096
rect 519629 81091 519695 81094
rect 523200 81064 524400 81094
rect 519997 80882 520063 80885
rect 518788 80880 520063 80882
rect 518788 80824 520002 80880
rect 520058 80824 520063 80880
rect 518788 80822 520063 80824
rect 519997 80819 520063 80822
rect 116761 79930 116827 79933
rect 116761 79928 119140 79930
rect 116761 79872 116766 79928
rect 116822 79872 119140 79928
rect 116761 79870 119140 79872
rect 116761 79867 116827 79870
rect 519997 79658 520063 79661
rect 523200 79658 524400 79688
rect 519997 79656 524400 79658
rect 519997 79600 520002 79656
rect 520058 79600 524400 79656
rect 519997 79598 524400 79600
rect 519997 79595 520063 79598
rect 523200 79568 524400 79598
rect 519077 79522 519143 79525
rect 518788 79520 519143 79522
rect 518788 79464 519082 79520
rect 519138 79464 519143 79520
rect 518788 79462 519143 79464
rect 519077 79459 519143 79462
rect 519261 78162 519327 78165
rect 518788 78160 519327 78162
rect 518788 78104 519266 78160
rect 519322 78104 519327 78160
rect 518788 78102 519327 78104
rect 519261 78099 519327 78102
rect 519721 78162 519787 78165
rect 523200 78162 524400 78192
rect 519721 78160 524400 78162
rect 519721 78104 519726 78160
rect 519782 78104 524400 78160
rect 519721 78102 524400 78104
rect 519721 78099 519787 78102
rect 523200 78072 524400 78102
rect 116669 78026 116735 78029
rect 116669 78024 119140 78026
rect 116669 77968 116674 78024
rect 116730 77968 119140 78024
rect 116669 77966 119140 77968
rect 116669 77963 116735 77966
rect 519445 76802 519511 76805
rect 518788 76800 519511 76802
rect 518788 76744 519450 76800
rect 519506 76744 519511 76800
rect 518788 76742 519511 76744
rect 519445 76739 519511 76742
rect 519077 76666 519143 76669
rect 523200 76666 524400 76696
rect 519077 76664 524400 76666
rect 519077 76608 519082 76664
rect 519138 76608 524400 76664
rect 519077 76606 524400 76608
rect 519077 76603 519143 76606
rect 523200 76576 524400 76606
rect 110860 75926 119140 75986
rect 519629 75306 519695 75309
rect 518788 75304 519695 75306
rect 518788 75248 519634 75304
rect 519690 75248 519695 75304
rect 518788 75246 519695 75248
rect 519629 75243 519695 75246
rect 519905 75170 519971 75173
rect 523200 75170 524400 75200
rect 519905 75168 524400 75170
rect 519905 75112 519910 75168
rect 519966 75112 524400 75168
rect 519905 75110 524400 75112
rect 519905 75107 519971 75110
rect 523200 75080 524400 75110
rect 116577 74082 116643 74085
rect 116577 74080 119140 74082
rect 116577 74024 116582 74080
rect 116638 74024 119140 74080
rect 116577 74022 119140 74024
rect 116577 74019 116643 74022
rect 519997 73946 520063 73949
rect 518788 73944 520063 73946
rect 518788 73888 520002 73944
rect 520058 73888 520063 73944
rect 518788 73886 520063 73888
rect 519997 73883 520063 73886
rect 519261 73674 519327 73677
rect 523200 73674 524400 73704
rect 519261 73672 524400 73674
rect 519261 73616 519266 73672
rect 519322 73616 524400 73672
rect 519261 73614 524400 73616
rect 519261 73611 519327 73614
rect 523200 73584 524400 73614
rect 519721 72586 519787 72589
rect 518788 72584 519787 72586
rect 518788 72528 519726 72584
rect 519782 72528 519787 72584
rect 518788 72526 519787 72528
rect 519721 72523 519787 72526
rect 116485 72178 116551 72181
rect 116485 72176 119140 72178
rect 116485 72120 116490 72176
rect 116546 72120 119140 72176
rect 116485 72118 119140 72120
rect 116485 72115 116551 72118
rect 520089 72042 520155 72045
rect 523200 72042 524400 72072
rect 520089 72040 524400 72042
rect 520089 71984 520094 72040
rect 520150 71984 524400 72040
rect 520089 71982 524400 71984
rect 520089 71979 520155 71982
rect 523200 71952 524400 71982
rect 519077 71226 519143 71229
rect 518788 71224 519143 71226
rect 518788 71168 519082 71224
rect 519138 71168 519143 71224
rect 518788 71166 519143 71168
rect 519077 71163 519143 71166
rect 520181 70546 520247 70549
rect 523200 70546 524400 70576
rect 520181 70544 524400 70546
rect 520181 70488 520186 70544
rect 520242 70488 524400 70544
rect 520181 70486 524400 70488
rect 520181 70483 520247 70486
rect 523200 70456 524400 70486
rect 116301 70274 116367 70277
rect 116301 70272 119140 70274
rect 116301 70216 116306 70272
rect 116362 70216 119140 70272
rect 116301 70214 119140 70216
rect 116301 70211 116367 70214
rect 519905 69866 519971 69869
rect 518788 69864 519971 69866
rect 518788 69808 519910 69864
rect 519966 69808 519971 69864
rect 518788 69806 519971 69808
rect 519905 69803 519971 69806
rect 519629 69050 519695 69053
rect 523200 69050 524400 69080
rect 519629 69048 524400 69050
rect 519629 68992 519634 69048
rect 519690 68992 524400 69048
rect 519629 68990 524400 68992
rect 519629 68987 519695 68990
rect 523200 68960 524400 68990
rect 519261 68506 519327 68509
rect 518788 68504 519327 68506
rect 518788 68448 519266 68504
rect 519322 68448 519327 68504
rect 518788 68446 519327 68448
rect 519261 68443 519327 68446
rect 116209 68370 116275 68373
rect 116209 68368 119140 68370
rect 116209 68312 116214 68368
rect 116270 68312 119140 68368
rect 116209 68310 119140 68312
rect 116209 68307 116275 68310
rect 520457 67554 520523 67557
rect 523200 67554 524400 67584
rect 520457 67552 524400 67554
rect 520457 67496 520462 67552
rect 520518 67496 524400 67552
rect 520457 67494 524400 67496
rect 520457 67491 520523 67494
rect 523200 67464 524400 67494
rect 520089 67146 520155 67149
rect 518788 67144 520155 67146
rect 518788 67088 520094 67144
rect 520150 67088 520155 67144
rect 518788 67086 520155 67088
rect 520089 67083 520155 67086
rect 117129 66466 117195 66469
rect 117129 66464 119140 66466
rect 117129 66408 117134 66464
rect 117190 66408 119140 66464
rect 117129 66406 119140 66408
rect 117129 66403 117195 66406
rect 520365 66058 520431 66061
rect 523200 66058 524400 66088
rect 520365 66056 524400 66058
rect 520365 66000 520370 66056
rect 520426 66000 524400 66056
rect 520365 65998 524400 66000
rect 520365 65995 520431 65998
rect 523200 65968 524400 65998
rect 520181 65786 520247 65789
rect 518788 65784 520247 65786
rect 518788 65728 520186 65784
rect 520242 65728 520247 65784
rect 518788 65726 520247 65728
rect 520181 65723 520247 65726
rect 113541 64562 113607 64565
rect 110860 64560 113607 64562
rect 110860 64504 113546 64560
rect 113602 64504 113607 64560
rect 110860 64502 113607 64504
rect 113541 64499 113607 64502
rect 115197 64562 115263 64565
rect 520733 64562 520799 64565
rect 523200 64562 524400 64592
rect 115197 64560 119140 64562
rect 115197 64504 115202 64560
rect 115258 64504 119140 64560
rect 115197 64502 119140 64504
rect 520733 64560 524400 64562
rect 520733 64504 520738 64560
rect 520794 64504 524400 64560
rect 520733 64502 524400 64504
rect 115197 64499 115263 64502
rect 520733 64499 520799 64502
rect 523200 64472 524400 64502
rect 519629 64426 519695 64429
rect 518788 64424 519695 64426
rect 518788 64368 519634 64424
rect 519690 64368 519695 64424
rect 518788 64366 519695 64368
rect 519629 64363 519695 64366
rect 520457 63066 520523 63069
rect 518788 63064 520523 63066
rect 518788 63008 520462 63064
rect 520518 63008 520523 63064
rect 518788 63006 520523 63008
rect 520457 63003 520523 63006
rect 521009 62930 521075 62933
rect 523200 62930 524400 62960
rect 521009 62928 524400 62930
rect 521009 62872 521014 62928
rect 521070 62872 524400 62928
rect 521009 62870 524400 62872
rect 521009 62867 521075 62870
rect 523200 62840 524400 62870
rect 116117 62658 116183 62661
rect 116117 62656 119140 62658
rect 116117 62600 116122 62656
rect 116178 62600 119140 62656
rect 116117 62598 119140 62600
rect 116117 62595 116183 62598
rect 520365 61706 520431 61709
rect 518788 61704 520431 61706
rect 518788 61648 520370 61704
rect 520426 61648 520431 61704
rect 518788 61646 520431 61648
rect 520365 61643 520431 61646
rect 521101 61434 521167 61437
rect 523200 61434 524400 61464
rect 521101 61432 524400 61434
rect 521101 61376 521106 61432
rect 521162 61376 524400 61432
rect 521101 61374 524400 61376
rect 521101 61371 521167 61374
rect 523200 61344 524400 61374
rect 116577 60618 116643 60621
rect 116577 60616 119140 60618
rect 116577 60560 116582 60616
rect 116638 60560 119140 60616
rect 116577 60558 119140 60560
rect 116577 60555 116643 60558
rect 520733 60346 520799 60349
rect 518788 60344 520799 60346
rect 518788 60288 520738 60344
rect 520794 60288 520799 60344
rect 518788 60286 520799 60288
rect 520733 60283 520799 60286
rect 520733 59938 520799 59941
rect 523200 59938 524400 59968
rect 520733 59936 524400 59938
rect 520733 59880 520738 59936
rect 520794 59880 524400 59936
rect 520733 59878 524400 59880
rect 520733 59875 520799 59878
rect 523200 59848 524400 59878
rect 521009 58986 521075 58989
rect 518788 58984 521075 58986
rect 518788 58928 521014 58984
rect 521070 58928 521075 58984
rect 518788 58926 521075 58928
rect 521009 58923 521075 58926
rect 116669 58714 116735 58717
rect 116669 58712 119140 58714
rect 116669 58656 116674 58712
rect 116730 58656 119140 58712
rect 116669 58654 119140 58656
rect 116669 58651 116735 58654
rect 521285 58442 521351 58445
rect 523200 58442 524400 58472
rect 521285 58440 524400 58442
rect 521285 58384 521290 58440
rect 521346 58384 524400 58440
rect 521285 58382 524400 58384
rect 521285 58379 521351 58382
rect 523200 58352 524400 58382
rect 521101 57490 521167 57493
rect 518788 57488 521167 57490
rect 518788 57432 521106 57488
rect 521162 57432 521167 57488
rect 518788 57430 521167 57432
rect 521101 57427 521167 57430
rect 520365 56946 520431 56949
rect 523200 56946 524400 56976
rect 520365 56944 524400 56946
rect 520365 56888 520370 56944
rect 520426 56888 524400 56944
rect 520365 56886 524400 56888
rect 520365 56883 520431 56886
rect 523200 56856 524400 56886
rect 116761 56810 116827 56813
rect 116761 56808 119140 56810
rect 116761 56752 116766 56808
rect 116822 56752 119140 56808
rect 116761 56750 119140 56752
rect 116761 56747 116827 56750
rect 520733 56130 520799 56133
rect 518788 56128 520799 56130
rect 518788 56072 520738 56128
rect 520794 56072 520799 56128
rect 518788 56070 520799 56072
rect 520733 56067 520799 56070
rect 520273 55450 520339 55453
rect 523200 55450 524400 55480
rect 520273 55448 524400 55450
rect 520273 55392 520278 55448
rect 520334 55392 524400 55448
rect 520273 55390 524400 55392
rect 520273 55387 520339 55390
rect 523200 55360 524400 55390
rect 116853 54906 116919 54909
rect 116853 54904 119140 54906
rect 116853 54848 116858 54904
rect 116914 54848 119140 54904
rect 116853 54846 119140 54848
rect 116853 54843 116919 54846
rect 521285 54770 521351 54773
rect 518788 54768 521351 54770
rect 518788 54712 521290 54768
rect 521346 54712 521351 54768
rect 518788 54710 521351 54712
rect 521285 54707 521351 54710
rect 519077 53818 519143 53821
rect 523200 53818 524400 53848
rect 519077 53816 524400 53818
rect 519077 53760 519082 53816
rect 519138 53760 524400 53816
rect 519077 53758 524400 53760
rect 519077 53755 519143 53758
rect 523200 53728 524400 53758
rect 520365 53410 520431 53413
rect 518788 53408 520431 53410
rect 518788 53352 520370 53408
rect 520426 53352 520431 53408
rect 518788 53350 520431 53352
rect 520365 53347 520431 53350
rect 113909 53138 113975 53141
rect 110860 53136 113975 53138
rect 110860 53080 113914 53136
rect 113970 53080 113975 53136
rect 110860 53078 113975 53080
rect 113909 53075 113975 53078
rect 116393 53002 116459 53005
rect 116393 53000 119140 53002
rect 116393 52944 116398 53000
rect 116454 52944 119140 53000
rect 116393 52942 119140 52944
rect 116393 52939 116459 52942
rect 519905 52322 519971 52325
rect 523200 52322 524400 52352
rect 519905 52320 524400 52322
rect 519905 52264 519910 52320
rect 519966 52264 524400 52320
rect 519905 52262 524400 52264
rect 519905 52259 519971 52262
rect 523200 52232 524400 52262
rect 520273 52050 520339 52053
rect 518788 52048 520339 52050
rect 518788 51992 520278 52048
rect 520334 51992 520339 52048
rect 518788 51990 520339 51992
rect 520273 51987 520339 51990
rect 116945 51098 117011 51101
rect 116945 51096 119140 51098
rect 116945 51040 116950 51096
rect 117006 51040 119140 51096
rect 116945 51038 119140 51040
rect 116945 51035 117011 51038
rect 519997 50826 520063 50829
rect 523200 50826 524400 50856
rect 519997 50824 524400 50826
rect 519997 50768 520002 50824
rect 520058 50768 524400 50824
rect 519997 50766 524400 50768
rect 519997 50763 520063 50766
rect 523200 50736 524400 50766
rect 519077 50690 519143 50693
rect 518788 50688 519143 50690
rect 518788 50632 519082 50688
rect 519138 50632 519143 50688
rect 518788 50630 519143 50632
rect 519077 50627 519143 50630
rect 519905 49330 519971 49333
rect 518788 49328 519971 49330
rect 518788 49272 519910 49328
rect 519966 49272 519971 49328
rect 518788 49270 519971 49272
rect 519905 49267 519971 49270
rect 520181 49330 520247 49333
rect 523200 49330 524400 49360
rect 520181 49328 524400 49330
rect 520181 49272 520186 49328
rect 520242 49272 524400 49328
rect 520181 49270 524400 49272
rect 520181 49267 520247 49270
rect 523200 49240 524400 49270
rect 115933 49194 115999 49197
rect 115933 49192 119140 49194
rect 115933 49136 115938 49192
rect 115994 49136 119140 49192
rect 115933 49134 119140 49136
rect 115933 49131 115999 49134
rect 519997 47970 520063 47973
rect 518788 47968 520063 47970
rect 518788 47912 520002 47968
rect 520058 47912 520063 47968
rect 518788 47910 520063 47912
rect 519997 47907 520063 47910
rect 519261 47834 519327 47837
rect 523200 47834 524400 47864
rect 519261 47832 524400 47834
rect 519261 47776 519266 47832
rect 519322 47776 524400 47832
rect 519261 47774 524400 47776
rect 519261 47771 519327 47774
rect 523200 47744 524400 47774
rect 116025 47154 116091 47157
rect 116025 47152 119140 47154
rect 116025 47096 116030 47152
rect 116086 47096 119140 47152
rect 116025 47094 119140 47096
rect 116025 47091 116091 47094
rect 520181 46610 520247 46613
rect 518788 46608 520247 46610
rect 518788 46552 520186 46608
rect 520242 46552 520247 46608
rect 518788 46550 520247 46552
rect 520181 46547 520247 46550
rect 519905 46338 519971 46341
rect 523200 46338 524400 46368
rect 519905 46336 524400 46338
rect 519905 46280 519910 46336
rect 519966 46280 524400 46336
rect 519905 46278 524400 46280
rect 519905 46275 519971 46278
rect 523200 46248 524400 46278
rect 117037 45250 117103 45253
rect 519261 45250 519327 45253
rect 117037 45248 119140 45250
rect 117037 45192 117042 45248
rect 117098 45192 119140 45248
rect 117037 45190 119140 45192
rect 518788 45248 519327 45250
rect 518788 45192 519266 45248
rect 519322 45192 519327 45248
rect 518788 45190 519327 45192
rect 117037 45187 117103 45190
rect 519261 45187 519327 45190
rect 519813 44706 519879 44709
rect 523200 44706 524400 44736
rect 519813 44704 524400 44706
rect 519813 44648 519818 44704
rect 519874 44648 524400 44704
rect 519813 44646 524400 44648
rect 519813 44643 519879 44646
rect 523200 44616 524400 44646
rect 519905 43890 519971 43893
rect 518788 43888 519971 43890
rect 518788 43832 519910 43888
rect 519966 43832 519971 43888
rect 518788 43830 519971 43832
rect 519905 43827 519971 43830
rect 117129 43346 117195 43349
rect 117129 43344 119140 43346
rect 117129 43288 117134 43344
rect 117190 43288 119140 43344
rect 117129 43286 119140 43288
rect 117129 43283 117195 43286
rect 520089 43210 520155 43213
rect 523200 43210 524400 43240
rect 520089 43208 524400 43210
rect 520089 43152 520094 43208
rect 520150 43152 524400 43208
rect 520089 43150 524400 43152
rect 520089 43147 520155 43150
rect 523200 43120 524400 43150
rect 519813 42530 519879 42533
rect 518788 42528 519879 42530
rect 518788 42472 519818 42528
rect 519874 42472 519879 42528
rect 518788 42470 519879 42472
rect 519813 42467 519879 42470
rect 114093 41850 114159 41853
rect 110860 41848 114159 41850
rect 110860 41792 114098 41848
rect 114154 41792 114159 41848
rect 110860 41790 114159 41792
rect 114093 41787 114159 41790
rect 520181 41714 520247 41717
rect 523200 41714 524400 41744
rect 520181 41712 524400 41714
rect 520181 41656 520186 41712
rect 520242 41656 524400 41712
rect 520181 41654 524400 41656
rect 520181 41651 520247 41654
rect 523200 41624 524400 41654
rect 115933 41442 115999 41445
rect 115933 41440 119140 41442
rect 115933 41384 115938 41440
rect 115994 41384 119140 41440
rect 115933 41382 119140 41384
rect 115933 41379 115999 41382
rect 520089 41170 520155 41173
rect 518788 41168 520155 41170
rect 518788 41112 520094 41168
rect 520150 41112 520155 41168
rect 518788 41110 520155 41112
rect 520089 41107 520155 41110
rect 519813 40218 519879 40221
rect 523200 40218 524400 40248
rect 519813 40216 524400 40218
rect 519813 40160 519818 40216
rect 519874 40160 524400 40216
rect 519813 40158 524400 40160
rect 519813 40155 519879 40158
rect 523200 40128 524400 40158
rect 520181 39810 520247 39813
rect 518788 39808 520247 39810
rect 518788 39752 520186 39808
rect 520242 39752 520247 39808
rect 518788 39750 520247 39752
rect 520181 39747 520247 39750
rect 115933 39538 115999 39541
rect 115933 39536 119140 39538
rect 115933 39480 115938 39536
rect 115994 39480 119140 39536
rect 115933 39478 119140 39480
rect 115933 39475 115999 39478
rect 520181 38722 520247 38725
rect 523200 38722 524400 38752
rect 520181 38720 524400 38722
rect 520181 38664 520186 38720
rect 520242 38664 524400 38720
rect 520181 38662 524400 38664
rect 520181 38659 520247 38662
rect 523200 38632 524400 38662
rect 519813 38314 519879 38317
rect 518788 38312 519879 38314
rect 518788 38256 519818 38312
rect 519874 38256 519879 38312
rect 518788 38254 519879 38256
rect 519813 38251 519879 38254
rect 116393 37634 116459 37637
rect 116393 37632 119140 37634
rect 116393 37576 116398 37632
rect 116454 37576 119140 37632
rect 116393 37574 119140 37576
rect 116393 37571 116459 37574
rect 521101 37226 521167 37229
rect 523200 37226 524400 37256
rect 521101 37224 524400 37226
rect 521101 37168 521106 37224
rect 521162 37168 524400 37224
rect 521101 37166 524400 37168
rect 521101 37163 521167 37166
rect 523200 37136 524400 37166
rect 520181 36954 520247 36957
rect 518788 36952 520247 36954
rect 518788 36896 520186 36952
rect 520242 36896 520247 36952
rect 518788 36894 520247 36896
rect 520181 36891 520247 36894
rect 521101 36002 521167 36005
rect 518758 36000 521167 36002
rect 518758 35944 521106 36000
rect 521162 35944 521167 36000
rect 518758 35942 521167 35944
rect 115933 35730 115999 35733
rect 115933 35728 119140 35730
rect 115933 35672 115938 35728
rect 115994 35672 119140 35728
rect 115933 35670 119140 35672
rect 115933 35667 115999 35670
rect 518758 35564 518818 35942
rect 521101 35939 521167 35942
rect 520917 35594 520983 35597
rect 523200 35594 524400 35624
rect 520917 35592 524400 35594
rect 520917 35536 520922 35592
rect 520978 35536 524400 35592
rect 520917 35534 524400 35536
rect 520917 35531 520983 35534
rect 523200 35504 524400 35534
rect 520917 34642 520983 34645
rect 518758 34640 520983 34642
rect 518758 34584 520922 34640
rect 520978 34584 520983 34640
rect 518758 34582 520983 34584
rect 518758 34204 518818 34582
rect 520917 34579 520983 34582
rect 520825 34098 520891 34101
rect 523200 34098 524400 34128
rect 520825 34096 524400 34098
rect 520825 34040 520830 34096
rect 520886 34040 524400 34096
rect 520825 34038 524400 34040
rect 520825 34035 520891 34038
rect 523200 34008 524400 34038
rect 116393 33826 116459 33829
rect 116393 33824 119140 33826
rect 116393 33768 116398 33824
rect 116454 33768 119140 33824
rect 116393 33766 119140 33768
rect 116393 33763 116459 33766
rect 520825 33282 520891 33285
rect 518758 33280 520891 33282
rect 518758 33224 520830 33280
rect 520886 33224 520891 33280
rect 518758 33222 520891 33224
rect 518758 32844 518818 33222
rect 520825 33219 520891 33222
rect 521101 32602 521167 32605
rect 523200 32602 524400 32632
rect 521101 32600 524400 32602
rect 521101 32544 521106 32600
rect 521162 32544 524400 32600
rect 521101 32542 524400 32544
rect 521101 32539 521167 32542
rect 523200 32512 524400 32542
rect 115933 31786 115999 31789
rect 521101 31786 521167 31789
rect 115933 31784 119140 31786
rect 115933 31728 115938 31784
rect 115994 31728 119140 31784
rect 115933 31726 119140 31728
rect 518758 31784 521167 31786
rect 518758 31728 521106 31784
rect 521162 31728 521167 31784
rect 518758 31726 521167 31728
rect 115933 31723 115999 31726
rect 518758 31484 518818 31726
rect 521101 31723 521167 31726
rect 521101 31106 521167 31109
rect 523200 31106 524400 31136
rect 521101 31104 524400 31106
rect 521101 31048 521106 31104
rect 521162 31048 524400 31104
rect 521101 31046 524400 31048
rect 521101 31043 521167 31046
rect 523200 31016 524400 31046
rect 114185 30426 114251 30429
rect 521101 30426 521167 30429
rect 110860 30424 114251 30426
rect 110860 30368 114190 30424
rect 114246 30368 114251 30424
rect 110860 30366 114251 30368
rect 114185 30363 114251 30366
rect 518758 30424 521167 30426
rect 518758 30368 521106 30424
rect 521162 30368 521167 30424
rect 518758 30366 521167 30368
rect 518758 30124 518818 30366
rect 521101 30363 521167 30366
rect 116117 29882 116183 29885
rect 116117 29880 119140 29882
rect 116117 29824 116122 29880
rect 116178 29824 119140 29880
rect 116117 29822 119140 29824
rect 116117 29819 116183 29822
rect 521101 29610 521167 29613
rect 523200 29610 524400 29640
rect 521101 29608 524400 29610
rect 521101 29552 521106 29608
rect 521162 29552 524400 29608
rect 521101 29550 524400 29552
rect 521101 29547 521167 29550
rect 523200 29520 524400 29550
rect 521101 28794 521167 28797
rect 518788 28792 521167 28794
rect 518788 28736 521106 28792
rect 521162 28736 521167 28792
rect 518788 28734 521167 28736
rect 521101 28731 521167 28734
rect 523200 28114 524400 28144
rect 518850 28054 524400 28114
rect 116117 27978 116183 27981
rect 518850 27978 518910 28054
rect 523200 28024 524400 28054
rect 116117 27976 119140 27978
rect 116117 27920 116122 27976
rect 116178 27920 119140 27976
rect 116117 27918 119140 27920
rect 518758 27918 518910 27978
rect 116117 27915 116183 27918
rect 518758 27404 518818 27918
rect 523200 26482 524400 26512
rect 518850 26422 524400 26482
rect 518850 26346 518910 26422
rect 523200 26392 524400 26422
rect 518758 26286 518910 26346
rect 116117 26074 116183 26077
rect 116117 26072 119140 26074
rect 116117 26016 116122 26072
rect 116178 26016 119140 26072
rect 518758 26044 518818 26286
rect 116117 26014 119140 26016
rect 116117 26011 116183 26014
rect 523200 24986 524400 25016
rect 518758 24926 524400 24986
rect 518758 24684 518818 24926
rect 523200 24896 524400 24926
rect 117221 24170 117287 24173
rect 117221 24168 119140 24170
rect 117221 24112 117226 24168
rect 117282 24112 119140 24168
rect 117221 24110 119140 24112
rect 117221 24107 117287 24110
rect 523200 23490 524400 23520
rect 518758 23430 524400 23490
rect 518758 23324 518818 23430
rect 523200 23400 524400 23430
rect 115933 22266 115999 22269
rect 115933 22264 119140 22266
rect 115933 22208 115938 22264
rect 115994 22208 119140 22264
rect 115933 22206 119140 22208
rect 115933 22203 115999 22206
rect 523200 21994 524400 22024
rect 518788 21934 524400 21994
rect 523200 21904 524400 21934
rect 521101 20498 521167 20501
rect 523200 20498 524400 20528
rect 521101 20496 524400 20498
rect 116117 20362 116183 20365
rect 116117 20360 119140 20362
rect 116117 20304 116122 20360
rect 116178 20304 119140 20360
rect 116117 20302 119140 20304
rect 116117 20299 116183 20302
rect 518758 19818 518818 20468
rect 521101 20440 521106 20496
rect 521162 20440 524400 20496
rect 521101 20438 524400 20440
rect 521101 20435 521167 20438
rect 523200 20408 524400 20438
rect 521101 19818 521167 19821
rect 518758 19816 521167 19818
rect 518758 19760 521106 19816
rect 521162 19760 521167 19816
rect 518758 19758 521167 19760
rect 521101 19755 521167 19758
rect 113633 19002 113699 19005
rect 110860 19000 113699 19002
rect 110860 18944 113638 19000
rect 113694 18944 113699 19000
rect 110860 18942 113699 18944
rect 113633 18939 113699 18942
rect 116301 18458 116367 18461
rect 518758 18458 518818 19108
rect 523200 19002 524400 19032
rect 521150 18942 524400 19002
rect 521150 18458 521210 18942
rect 523200 18912 524400 18942
rect 116301 18456 119140 18458
rect 116301 18400 116306 18456
rect 116362 18400 119140 18456
rect 116301 18398 119140 18400
rect 518758 18398 521210 18458
rect 116301 18395 116367 18398
rect 518758 17098 518818 17748
rect 523200 17370 524400 17400
rect 521150 17310 524400 17370
rect 521150 17098 521210 17310
rect 523200 17280 524400 17310
rect 518758 17038 521210 17098
rect 116393 16418 116459 16421
rect 116393 16416 119140 16418
rect 116393 16360 116398 16416
rect 116454 16360 119140 16416
rect 116393 16358 119140 16360
rect 116393 16355 116459 16358
rect 518758 15738 518818 16388
rect 523200 15874 524400 15904
rect 521104 15814 524400 15874
rect 521104 15738 521164 15814
rect 523200 15784 524400 15814
rect 518758 15678 521164 15738
rect 521101 15058 521167 15061
rect 518788 15056 521167 15058
rect 518788 15000 521106 15056
rect 521162 15000 521167 15056
rect 518788 14998 521167 15000
rect 521101 14995 521167 14998
rect 116209 14514 116275 14517
rect 116209 14512 119140 14514
rect 116209 14456 116214 14512
rect 116270 14456 119140 14512
rect 116209 14454 119140 14456
rect 116209 14451 116275 14454
rect 521101 14378 521167 14381
rect 523200 14378 524400 14408
rect 521101 14376 524400 14378
rect 521101 14320 521106 14376
rect 521162 14320 524400 14376
rect 521101 14318 524400 14320
rect 521101 14315 521167 14318
rect 523200 14288 524400 14318
rect 521101 13698 521167 13701
rect 518788 13696 521167 13698
rect 518788 13640 521106 13696
rect 521162 13640 521167 13696
rect 518788 13638 521167 13640
rect 521101 13635 521167 13638
rect 521101 12882 521167 12885
rect 523200 12882 524400 12912
rect 521101 12880 524400 12882
rect 521101 12824 521106 12880
rect 521162 12824 524400 12880
rect 521101 12822 524400 12824
rect 521101 12819 521167 12822
rect 523200 12792 524400 12822
rect 116526 12548 116532 12612
rect 116596 12610 116602 12612
rect 116596 12550 119140 12610
rect 116596 12548 116602 12550
rect 519629 12338 519695 12341
rect 518788 12336 519695 12338
rect 518788 12280 519634 12336
rect 519690 12280 519695 12336
rect 518788 12278 519695 12280
rect 519629 12275 519695 12278
rect 519629 11386 519695 11389
rect 523200 11386 524400 11416
rect 519629 11384 524400 11386
rect 519629 11328 519634 11384
rect 519690 11328 524400 11384
rect 519629 11326 524400 11328
rect 519629 11323 519695 11326
rect 523200 11296 524400 11326
rect 521101 10978 521167 10981
rect 518788 10976 521167 10978
rect 518788 10920 521106 10976
rect 521162 10920 521167 10976
rect 518788 10918 521167 10920
rect 521101 10915 521167 10918
rect 113766 10644 113772 10708
rect 113836 10706 113842 10708
rect 113836 10646 119140 10706
rect 113836 10644 113842 10646
rect 521101 9890 521167 9893
rect 523200 9890 524400 9920
rect 521101 9888 524400 9890
rect 521101 9832 521106 9888
rect 521162 9832 524400 9888
rect 521101 9830 524400 9832
rect 521101 9827 521167 9830
rect 523200 9800 524400 9830
rect 521101 9618 521167 9621
rect 518788 9616 521167 9618
rect 518788 9560 521106 9616
rect 521162 9560 521167 9616
rect 518788 9558 521167 9560
rect 521101 9555 521167 9558
rect 117078 8740 117084 8804
rect 117148 8802 117154 8804
rect 117148 8742 119140 8802
rect 117148 8740 117154 8742
rect 520365 8258 520431 8261
rect 518788 8256 520431 8258
rect 518788 8200 520370 8256
rect 520426 8200 520431 8256
rect 518788 8198 520431 8200
rect 520365 8195 520431 8198
rect 521101 8258 521167 8261
rect 523200 8258 524400 8288
rect 521101 8256 524400 8258
rect 521101 8200 521106 8256
rect 521162 8200 524400 8256
rect 521101 8198 524400 8200
rect 521101 8195 521167 8198
rect 523200 8168 524400 8198
rect 113633 7714 113699 7717
rect 110860 7712 113699 7714
rect 110860 7656 113638 7712
rect 113694 7656 113699 7712
rect 110860 7654 113699 7656
rect 113633 7651 113699 7654
rect 116158 6836 116164 6900
rect 116228 6898 116234 6900
rect 521101 6898 521167 6901
rect 116228 6838 119140 6898
rect 518788 6896 521167 6898
rect 518788 6840 521106 6896
rect 521162 6840 521167 6896
rect 518788 6838 521167 6840
rect 116228 6836 116234 6838
rect 521101 6835 521167 6838
rect 520365 6762 520431 6765
rect 523200 6762 524400 6792
rect 520365 6760 524400 6762
rect 520365 6704 520370 6760
rect 520426 6704 524400 6760
rect 520365 6702 524400 6704
rect 520365 6699 520431 6702
rect 523200 6672 524400 6702
rect 521009 5538 521075 5541
rect 518788 5536 521075 5538
rect 518788 5480 521014 5536
rect 521070 5480 521075 5536
rect 518788 5478 521075 5480
rect 521009 5475 521075 5478
rect 521101 5266 521167 5269
rect 523200 5266 524400 5296
rect 521101 5264 524400 5266
rect 521101 5208 521106 5264
rect 521162 5208 524400 5264
rect 521101 5206 524400 5208
rect 521101 5203 521167 5206
rect 523200 5176 524400 5206
rect 116117 4994 116183 4997
rect 116117 4992 119140 4994
rect 116117 4936 116122 4992
rect 116178 4936 119140 4992
rect 116117 4934 119140 4936
rect 116117 4931 116183 4934
rect 521101 4178 521167 4181
rect 518788 4176 521167 4178
rect 518788 4120 521106 4176
rect 521162 4120 521167 4176
rect 518788 4118 521167 4120
rect 521101 4115 521167 4118
rect 521009 3770 521075 3773
rect 523200 3770 524400 3800
rect 521009 3768 524400 3770
rect 521009 3712 521014 3768
rect 521070 3712 524400 3768
rect 521009 3710 524400 3712
rect 521009 3707 521075 3710
rect 523200 3680 524400 3710
rect 116117 3090 116183 3093
rect 116117 3088 119140 3090
rect 116117 3032 116122 3088
rect 116178 3032 119140 3088
rect 116117 3030 119140 3032
rect 116117 3027 116183 3030
rect 519997 2818 520063 2821
rect 518788 2816 520063 2818
rect 518788 2760 520002 2816
rect 520058 2760 520063 2816
rect 518788 2758 520063 2760
rect 519997 2755 520063 2758
rect 33041 2274 33107 2277
rect 111333 2274 111399 2277
rect 33041 2272 111399 2274
rect 33041 2216 33046 2272
rect 33102 2216 111338 2272
rect 111394 2216 111399 2272
rect 33041 2214 111399 2216
rect 33041 2211 33107 2214
rect 111333 2211 111399 2214
rect 521101 2274 521167 2277
rect 523200 2274 524400 2304
rect 521101 2272 524400 2274
rect 521101 2216 521106 2272
rect 521162 2216 524400 2272
rect 521101 2214 524400 2216
rect 521101 2211 521167 2214
rect 523200 2184 524400 2214
rect 29545 2138 29611 2141
rect 109677 2138 109743 2141
rect 29545 2136 109743 2138
rect 29545 2080 29550 2136
rect 29606 2080 109682 2136
rect 109738 2080 109743 2136
rect 29545 2078 109743 2080
rect 29545 2075 29611 2078
rect 109677 2075 109743 2078
rect 26049 2002 26115 2005
rect 109861 2002 109927 2005
rect 26049 2000 109927 2002
rect 26049 1944 26054 2000
rect 26110 1944 109866 2000
rect 109922 1944 109927 2000
rect 26049 1942 109927 1944
rect 26049 1939 26115 1942
rect 109861 1939 109927 1942
rect 19333 1866 19399 1869
rect 116526 1866 116532 1868
rect 19333 1864 116532 1866
rect 19333 1808 19338 1864
rect 19394 1808 116532 1864
rect 19333 1806 116532 1808
rect 19333 1803 19399 1806
rect 116526 1804 116532 1806
rect 116596 1804 116602 1868
rect 5993 1730 6059 1733
rect 109953 1730 110019 1733
rect 5993 1728 110019 1730
rect 5993 1672 5998 1728
rect 6054 1672 109958 1728
rect 110014 1672 110019 1728
rect 5993 1670 110019 1672
rect 5993 1667 6059 1670
rect 109953 1667 110019 1670
rect 229277 1730 229343 1733
rect 293585 1730 293651 1733
rect 229277 1728 293651 1730
rect 229277 1672 229282 1728
rect 229338 1672 293590 1728
rect 293646 1672 293651 1728
rect 229277 1670 293651 1672
rect 229277 1667 229343 1670
rect 293585 1667 293651 1670
rect 9305 1594 9371 1597
rect 116158 1594 116164 1596
rect 9305 1592 116164 1594
rect 9305 1536 9310 1592
rect 9366 1536 116164 1592
rect 9305 1534 116164 1536
rect 9305 1531 9371 1534
rect 116158 1532 116164 1534
rect 116228 1532 116234 1596
rect 163773 1594 163839 1597
rect 243629 1594 243695 1597
rect 163773 1592 243695 1594
rect 163773 1536 163778 1592
rect 163834 1536 243634 1592
rect 243690 1536 243695 1592
rect 163773 1534 243695 1536
rect 163773 1531 163839 1534
rect 243629 1531 243695 1534
rect 55949 1458 56015 1461
rect 294781 1458 294847 1461
rect 343633 1458 343699 1461
rect 55949 1456 343699 1458
rect 55949 1400 55954 1456
rect 56010 1400 294786 1456
rect 294842 1400 343638 1456
rect 343694 1400 343699 1456
rect 55949 1398 343699 1400
rect 55949 1395 56015 1398
rect 294781 1395 294847 1398
rect 343633 1395 343699 1398
rect 360285 1458 360351 1461
rect 393589 1458 393655 1461
rect 360285 1456 393655 1458
rect 360285 1400 360290 1456
rect 360346 1400 393594 1456
rect 393650 1400 393655 1456
rect 360285 1398 393655 1400
rect 360285 1395 360351 1398
rect 393589 1395 393655 1398
rect 425789 1458 425855 1461
rect 443637 1458 443703 1461
rect 425789 1456 443703 1458
rect 425789 1400 425794 1456
rect 425850 1400 443642 1456
rect 443698 1400 443703 1456
rect 425789 1398 443703 1400
rect 425789 1395 425855 1398
rect 443637 1395 443703 1398
rect 100753 1322 100819 1325
rect 117078 1322 117084 1324
rect 100753 1320 117084 1322
rect 100753 1264 100758 1320
rect 100814 1264 117084 1320
rect 100753 1262 117084 1264
rect 100753 1259 100819 1262
rect 117078 1260 117084 1262
rect 117148 1260 117154 1324
rect 98637 1186 98703 1189
rect 113766 1186 113772 1188
rect 98637 1184 113772 1186
rect 98637 1128 98642 1184
rect 98698 1128 113772 1184
rect 98637 1126 113772 1128
rect 98637 1123 98703 1126
rect 113766 1124 113772 1126
rect 113836 1124 113842 1188
rect 519997 778 520063 781
rect 523200 778 524400 808
rect 519997 776 524400 778
rect 519997 720 520002 776
rect 520058 720 524400 776
rect 519997 718 524400 720
rect 519997 715 520063 718
rect 523200 688 524400 718
<< via3 >>
rect 116532 151812 116596 151876
rect 116532 89388 116596 89452
rect 116532 12548 116596 12612
rect 113772 10644 113836 10708
rect 117084 8740 117148 8804
rect 116164 6836 116228 6900
rect 116532 1804 116596 1868
rect 116164 1532 116228 1596
rect 117084 1260 117148 1324
rect 113772 1124 113836 1188
<< metal4 >>
rect 116531 151876 116597 151877
rect 116531 151812 116532 151876
rect 116596 151812 116597 151876
rect 116531 151811 116597 151812
rect 1664 144454 1984 144496
rect 1664 144218 1706 144454
rect 1942 144218 1984 144454
rect 1664 144134 1984 144218
rect 1664 143898 1706 144134
rect 1942 143898 1984 144134
rect 1664 143856 1984 143898
rect 109956 144454 110276 144496
rect 109956 144218 109998 144454
rect 110234 144218 110276 144454
rect 109956 144134 110276 144218
rect 109956 143898 109998 144134
rect 110234 143898 110276 144134
rect 109956 143856 110276 143898
rect 1096 131454 1332 131496
rect 1096 131134 1332 131218
rect 1096 130856 1332 130898
rect 110616 131454 110936 131496
rect 110616 131218 110658 131454
rect 110894 131218 110936 131454
rect 110616 131134 110936 131218
rect 110616 130898 110658 131134
rect 110894 130898 110936 131134
rect 110616 130856 110936 130898
rect 1664 118454 1984 118496
rect 1664 118218 1706 118454
rect 1942 118218 1984 118454
rect 1664 118134 1984 118218
rect 1664 117898 1706 118134
rect 1942 117898 1984 118134
rect 1664 117856 1984 117898
rect 109956 118454 110276 118496
rect 109956 118218 109998 118454
rect 110234 118218 110276 118454
rect 109956 118134 110276 118218
rect 109956 117898 109998 118134
rect 110234 117898 110276 118134
rect 109956 117856 110276 117898
rect 1096 105454 1332 105496
rect 1096 105134 1332 105218
rect 1096 104856 1332 104898
rect 110616 105454 110936 105496
rect 110616 105218 110658 105454
rect 110894 105218 110936 105454
rect 110616 105134 110936 105218
rect 110616 104898 110658 105134
rect 110894 104898 110936 105134
rect 110616 104856 110936 104898
rect 1664 92454 1984 92496
rect 1664 92218 1706 92454
rect 1942 92218 1984 92454
rect 1664 92134 1984 92218
rect 1664 91898 1706 92134
rect 1942 91898 1984 92134
rect 1664 91856 1984 91898
rect 109956 92454 110276 92496
rect 109956 92218 109998 92454
rect 110234 92218 110276 92454
rect 109956 92134 110276 92218
rect 109956 91898 109998 92134
rect 110234 91898 110276 92134
rect 109956 91856 110276 91898
rect 116534 89453 116594 151811
rect 119664 144454 119984 144496
rect 119664 144218 119706 144454
rect 119942 144218 119984 144454
rect 119664 144134 119984 144218
rect 119664 143898 119706 144134
rect 119942 143898 119984 144134
rect 119664 143856 119984 143898
rect 517940 144454 518260 144496
rect 517940 144218 517982 144454
rect 518218 144218 518260 144454
rect 517940 144134 518260 144218
rect 517940 143898 517982 144134
rect 518218 143898 518260 144134
rect 517940 143856 518260 143898
rect 119004 131454 119324 131496
rect 119004 131218 119046 131454
rect 119282 131218 119324 131454
rect 119004 131134 119324 131218
rect 119004 130898 119046 131134
rect 119282 130898 119324 131134
rect 119004 130856 119324 130898
rect 518600 131454 518920 131496
rect 518600 131218 518642 131454
rect 518878 131218 518920 131454
rect 518600 131134 518920 131218
rect 518600 130898 518642 131134
rect 518878 130898 518920 131134
rect 518600 130856 518920 130898
rect 119664 118454 119984 118496
rect 119664 118218 119706 118454
rect 119942 118218 119984 118454
rect 119664 118134 119984 118218
rect 119664 117898 119706 118134
rect 119942 117898 119984 118134
rect 119664 117856 119984 117898
rect 517940 118454 518260 118496
rect 517940 118218 517982 118454
rect 518218 118218 518260 118454
rect 517940 118134 518260 118218
rect 517940 117898 517982 118134
rect 518218 117898 518260 118134
rect 517940 117856 518260 117898
rect 119004 105454 119324 105496
rect 119004 105218 119046 105454
rect 119282 105218 119324 105454
rect 119004 105134 119324 105218
rect 119004 104898 119046 105134
rect 119282 104898 119324 105134
rect 119004 104856 119324 104898
rect 518600 105454 518920 105496
rect 518600 105218 518642 105454
rect 518878 105218 518920 105454
rect 518600 105134 518920 105218
rect 518600 104898 518642 105134
rect 518878 104898 518920 105134
rect 518600 104856 518920 104898
rect 119664 92454 119984 92496
rect 119664 92218 119706 92454
rect 119942 92218 119984 92454
rect 119664 92134 119984 92218
rect 119664 91898 119706 92134
rect 119942 91898 119984 92134
rect 119664 91856 119984 91898
rect 517940 92454 518260 92496
rect 517940 92218 517982 92454
rect 518218 92218 518260 92454
rect 517940 92134 518260 92218
rect 517940 91898 517982 92134
rect 518218 91898 518260 92134
rect 517940 91856 518260 91898
rect 116531 89452 116597 89453
rect 116531 89388 116532 89452
rect 116596 89388 116597 89452
rect 116531 89387 116597 89388
rect 1096 79454 1332 79496
rect 1096 79134 1332 79218
rect 1096 78856 1332 78898
rect 110616 79454 110936 79496
rect 110616 79218 110658 79454
rect 110894 79218 110936 79454
rect 110616 79134 110936 79218
rect 110616 78898 110658 79134
rect 110894 78898 110936 79134
rect 110616 78856 110936 78898
rect 119004 79454 119324 79496
rect 119004 79218 119046 79454
rect 119282 79218 119324 79454
rect 119004 79134 119324 79218
rect 119004 78898 119046 79134
rect 119282 78898 119324 79134
rect 119004 78856 119324 78898
rect 518600 79454 518920 79496
rect 518600 79218 518642 79454
rect 518878 79218 518920 79454
rect 518600 79134 518920 79218
rect 518600 78898 518642 79134
rect 518878 78898 518920 79134
rect 518600 78856 518920 78898
rect 1664 66454 1984 66496
rect 1664 66218 1706 66454
rect 1942 66218 1984 66454
rect 1664 66134 1984 66218
rect 1664 65898 1706 66134
rect 1942 65898 1984 66134
rect 1664 65856 1984 65898
rect 109956 66454 110276 66496
rect 109956 66218 109998 66454
rect 110234 66218 110276 66454
rect 109956 66134 110276 66218
rect 109956 65898 109998 66134
rect 110234 65898 110276 66134
rect 109956 65856 110276 65898
rect 119664 66454 119984 66496
rect 119664 66218 119706 66454
rect 119942 66218 119984 66454
rect 119664 66134 119984 66218
rect 119664 65898 119706 66134
rect 119942 65898 119984 66134
rect 119664 65856 119984 65898
rect 517940 66454 518260 66496
rect 517940 66218 517982 66454
rect 518218 66218 518260 66454
rect 517940 66134 518260 66218
rect 517940 65898 517982 66134
rect 518218 65898 518260 66134
rect 517940 65856 518260 65898
rect 1096 53454 1332 53496
rect 1096 53134 1332 53218
rect 1096 52856 1332 52898
rect 110616 53454 110936 53496
rect 110616 53218 110658 53454
rect 110894 53218 110936 53454
rect 110616 53134 110936 53218
rect 110616 52898 110658 53134
rect 110894 52898 110936 53134
rect 110616 52856 110936 52898
rect 119004 53454 119324 53496
rect 119004 53218 119046 53454
rect 119282 53218 119324 53454
rect 119004 53134 119324 53218
rect 119004 52898 119046 53134
rect 119282 52898 119324 53134
rect 119004 52856 119324 52898
rect 518600 53454 518920 53496
rect 518600 53218 518642 53454
rect 518878 53218 518920 53454
rect 518600 53134 518920 53218
rect 518600 52898 518642 53134
rect 518878 52898 518920 53134
rect 518600 52856 518920 52898
rect 1664 40454 1984 40496
rect 1664 40218 1706 40454
rect 1942 40218 1984 40454
rect 1664 40134 1984 40218
rect 1664 39898 1706 40134
rect 1942 39898 1984 40134
rect 1664 39856 1984 39898
rect 109956 40454 110276 40496
rect 109956 40218 109998 40454
rect 110234 40218 110276 40454
rect 109956 40134 110276 40218
rect 109956 39898 109998 40134
rect 110234 39898 110276 40134
rect 109956 39856 110276 39898
rect 119664 40454 119984 40496
rect 119664 40218 119706 40454
rect 119942 40218 119984 40454
rect 119664 40134 119984 40218
rect 119664 39898 119706 40134
rect 119942 39898 119984 40134
rect 119664 39856 119984 39898
rect 517940 40454 518260 40496
rect 517940 40218 517982 40454
rect 518218 40218 518260 40454
rect 517940 40134 518260 40218
rect 517940 39898 517982 40134
rect 518218 39898 518260 40134
rect 517940 39856 518260 39898
rect 1096 27454 1332 27496
rect 1096 27134 1332 27218
rect 1096 26856 1332 26898
rect 110616 27454 110936 27496
rect 110616 27218 110658 27454
rect 110894 27218 110936 27454
rect 110616 27134 110936 27218
rect 110616 26898 110658 27134
rect 110894 26898 110936 27134
rect 110616 26856 110936 26898
rect 119004 27454 119324 27496
rect 119004 27218 119046 27454
rect 119282 27218 119324 27454
rect 119004 27134 119324 27218
rect 119004 26898 119046 27134
rect 119282 26898 119324 27134
rect 119004 26856 119324 26898
rect 518600 27454 518920 27496
rect 518600 27218 518642 27454
rect 518878 27218 518920 27454
rect 518600 27134 518920 27218
rect 518600 26898 518642 27134
rect 518878 26898 518920 27134
rect 518600 26856 518920 26898
rect 1664 14454 1984 14496
rect 1664 14218 1706 14454
rect 1942 14218 1984 14454
rect 1664 14134 1984 14218
rect 1664 13898 1706 14134
rect 1942 13898 1984 14134
rect 1664 13856 1984 13898
rect 109956 14454 110276 14496
rect 109956 14218 109998 14454
rect 110234 14218 110276 14454
rect 109956 14134 110276 14218
rect 109956 13898 109998 14134
rect 110234 13898 110276 14134
rect 109956 13856 110276 13898
rect 119664 14454 119984 14496
rect 119664 14218 119706 14454
rect 119942 14218 119984 14454
rect 119664 14134 119984 14218
rect 119664 13898 119706 14134
rect 119942 13898 119984 14134
rect 119664 13856 119984 13898
rect 517940 14454 518260 14496
rect 517940 14218 517982 14454
rect 518218 14218 518260 14454
rect 517940 14134 518260 14218
rect 517940 13898 517982 14134
rect 518218 13898 518260 14134
rect 517940 13856 518260 13898
rect 116531 12612 116597 12613
rect 116531 12548 116532 12612
rect 116596 12548 116597 12612
rect 116531 12547 116597 12548
rect 113771 10708 113837 10709
rect 113771 10644 113772 10708
rect 113836 10644 113837 10708
rect 113771 10643 113837 10644
rect 113774 1189 113834 10643
rect 116163 6900 116229 6901
rect 116163 6836 116164 6900
rect 116228 6836 116229 6900
rect 116163 6835 116229 6836
rect 116166 1597 116226 6835
rect 116534 1869 116594 12547
rect 117083 8804 117149 8805
rect 117083 8740 117084 8804
rect 117148 8740 117149 8804
rect 117083 8739 117149 8740
rect 116531 1868 116597 1869
rect 116531 1804 116532 1868
rect 116596 1804 116597 1868
rect 116531 1803 116597 1804
rect 116163 1596 116229 1597
rect 116163 1532 116164 1596
rect 116228 1532 116229 1596
rect 116163 1531 116229 1532
rect 117086 1325 117146 8739
rect 117083 1324 117149 1325
rect 117083 1260 117084 1324
rect 117148 1260 117149 1324
rect 117083 1259 117149 1260
rect 113771 1188 113837 1189
rect 113771 1124 113772 1188
rect 113836 1124 113837 1188
rect 113771 1123 113837 1124
<< via4 >>
rect 1706 144218 1942 144454
rect 1706 143898 1942 144134
rect 109998 144218 110234 144454
rect 109998 143898 110234 144134
rect 1096 131218 1332 131454
rect 1096 130898 1332 131134
rect 110658 131218 110894 131454
rect 110658 130898 110894 131134
rect 1706 118218 1942 118454
rect 1706 117898 1942 118134
rect 109998 118218 110234 118454
rect 109998 117898 110234 118134
rect 1096 105218 1332 105454
rect 1096 104898 1332 105134
rect 110658 105218 110894 105454
rect 110658 104898 110894 105134
rect 1706 92218 1942 92454
rect 1706 91898 1942 92134
rect 109998 92218 110234 92454
rect 109998 91898 110234 92134
rect 119706 144218 119942 144454
rect 119706 143898 119942 144134
rect 517982 144218 518218 144454
rect 517982 143898 518218 144134
rect 119046 131218 119282 131454
rect 119046 130898 119282 131134
rect 518642 131218 518878 131454
rect 518642 130898 518878 131134
rect 119706 118218 119942 118454
rect 119706 117898 119942 118134
rect 517982 118218 518218 118454
rect 517982 117898 518218 118134
rect 119046 105218 119282 105454
rect 119046 104898 119282 105134
rect 518642 105218 518878 105454
rect 518642 104898 518878 105134
rect 119706 92218 119942 92454
rect 119706 91898 119942 92134
rect 517982 92218 518218 92454
rect 517982 91898 518218 92134
rect 1096 79218 1332 79454
rect 1096 78898 1332 79134
rect 110658 79218 110894 79454
rect 110658 78898 110894 79134
rect 119046 79218 119282 79454
rect 119046 78898 119282 79134
rect 518642 79218 518878 79454
rect 518642 78898 518878 79134
rect 1706 66218 1942 66454
rect 1706 65898 1942 66134
rect 109998 66218 110234 66454
rect 109998 65898 110234 66134
rect 119706 66218 119942 66454
rect 119706 65898 119942 66134
rect 517982 66218 518218 66454
rect 517982 65898 518218 66134
rect 1096 53218 1332 53454
rect 1096 52898 1332 53134
rect 110658 53218 110894 53454
rect 110658 52898 110894 53134
rect 119046 53218 119282 53454
rect 119046 52898 119282 53134
rect 518642 53218 518878 53454
rect 518642 52898 518878 53134
rect 1706 40218 1942 40454
rect 1706 39898 1942 40134
rect 109998 40218 110234 40454
rect 109998 39898 110234 40134
rect 119706 40218 119942 40454
rect 119706 39898 119942 40134
rect 517982 40218 518218 40454
rect 517982 39898 518218 40134
rect 1096 27218 1332 27454
rect 1096 26898 1332 27134
rect 110658 27218 110894 27454
rect 110658 26898 110894 27134
rect 119046 27218 119282 27454
rect 119046 26898 119282 27134
rect 518642 27218 518878 27454
rect 518642 26898 518878 27134
rect 1706 14218 1942 14454
rect 1706 13898 1942 14134
rect 109998 14218 110234 14454
rect 109998 13898 110234 14134
rect 119706 14218 119942 14454
rect 119706 13898 119942 14134
rect 517982 14218 518218 14454
rect 517982 13898 518218 14134
<< metal5 >>
rect 1104 156856 522836 157496
rect 1104 144454 2200 144496
rect 1104 144218 1706 144454
rect 1942 144218 2200 144454
rect 1104 144134 2200 144218
rect 1104 143898 1706 144134
rect 1942 143898 2200 144134
rect 1104 143856 2200 143898
rect 109800 144454 120200 144496
rect 109800 144218 109998 144454
rect 110234 144218 119706 144454
rect 119942 144218 120200 144454
rect 109800 144134 120200 144218
rect 109800 143898 109998 144134
rect 110234 143898 119706 144134
rect 119942 143898 120200 144134
rect 109800 143856 120200 143898
rect 517800 144454 522836 144496
rect 517800 144218 517982 144454
rect 518218 144218 522836 144454
rect 517800 144134 522836 144218
rect 517800 143898 517982 144134
rect 518218 143898 522836 144134
rect 517800 143856 522836 143898
rect 1072 131454 2200 131496
rect 1072 131218 1096 131454
rect 1332 131218 2200 131454
rect 1072 131134 2200 131218
rect 1072 130898 1096 131134
rect 1332 130898 2200 131134
rect 1072 130856 2200 130898
rect 109800 131454 120200 131496
rect 109800 131218 110658 131454
rect 110894 131218 119046 131454
rect 119282 131218 120200 131454
rect 109800 131134 120200 131218
rect 109800 130898 110658 131134
rect 110894 130898 119046 131134
rect 119282 130898 120200 131134
rect 109800 130856 120200 130898
rect 517800 131454 522836 131496
rect 517800 131218 518642 131454
rect 518878 131218 522836 131454
rect 517800 131134 522836 131218
rect 517800 130898 518642 131134
rect 518878 130898 522836 131134
rect 517800 130856 522836 130898
rect 1104 118454 2200 118496
rect 1104 118218 1706 118454
rect 1942 118218 2200 118454
rect 1104 118134 2200 118218
rect 1104 117898 1706 118134
rect 1942 117898 2200 118134
rect 1104 117856 2200 117898
rect 109800 118454 120200 118496
rect 109800 118218 109998 118454
rect 110234 118218 119706 118454
rect 119942 118218 120200 118454
rect 109800 118134 120200 118218
rect 109800 117898 109998 118134
rect 110234 117898 119706 118134
rect 119942 117898 120200 118134
rect 109800 117856 120200 117898
rect 517800 118454 522836 118496
rect 517800 118218 517982 118454
rect 518218 118218 522836 118454
rect 517800 118134 522836 118218
rect 517800 117898 517982 118134
rect 518218 117898 522836 118134
rect 517800 117856 522836 117898
rect 1072 105454 2200 105496
rect 1072 105218 1096 105454
rect 1332 105218 2200 105454
rect 1072 105134 2200 105218
rect 1072 104898 1096 105134
rect 1332 104898 2200 105134
rect 1072 104856 2200 104898
rect 109800 105454 120200 105496
rect 109800 105218 110658 105454
rect 110894 105218 119046 105454
rect 119282 105218 120200 105454
rect 109800 105134 120200 105218
rect 109800 104898 110658 105134
rect 110894 104898 119046 105134
rect 119282 104898 120200 105134
rect 109800 104856 120200 104898
rect 517800 105454 522836 105496
rect 517800 105218 518642 105454
rect 518878 105218 522836 105454
rect 517800 105134 522836 105218
rect 517800 104898 518642 105134
rect 518878 104898 522836 105134
rect 517800 104856 522836 104898
rect 1104 92454 2200 92496
rect 1104 92218 1706 92454
rect 1942 92218 2200 92454
rect 1104 92134 2200 92218
rect 1104 91898 1706 92134
rect 1942 91898 2200 92134
rect 1104 91856 2200 91898
rect 109800 92454 120200 92496
rect 109800 92218 109998 92454
rect 110234 92218 119706 92454
rect 119942 92218 120200 92454
rect 109800 92134 120200 92218
rect 109800 91898 109998 92134
rect 110234 91898 119706 92134
rect 119942 91898 120200 92134
rect 109800 91856 120200 91898
rect 517800 92454 522836 92496
rect 517800 92218 517982 92454
rect 518218 92218 522836 92454
rect 517800 92134 522836 92218
rect 517800 91898 517982 92134
rect 518218 91898 522836 92134
rect 517800 91856 522836 91898
rect 1072 79454 2200 79496
rect 1072 79218 1096 79454
rect 1332 79218 2200 79454
rect 1072 79134 2200 79218
rect 1072 78898 1096 79134
rect 1332 78898 2200 79134
rect 1072 78856 2200 78898
rect 109800 79454 120200 79496
rect 109800 79218 110658 79454
rect 110894 79218 119046 79454
rect 119282 79218 120200 79454
rect 109800 79134 120200 79218
rect 109800 78898 110658 79134
rect 110894 78898 119046 79134
rect 119282 78898 120200 79134
rect 109800 78856 120200 78898
rect 517800 79454 522836 79496
rect 517800 79218 518642 79454
rect 518878 79218 522836 79454
rect 517800 79134 522836 79218
rect 517800 78898 518642 79134
rect 518878 78898 522836 79134
rect 517800 78856 522836 78898
rect 1104 66454 2200 66496
rect 1104 66218 1706 66454
rect 1942 66218 2200 66454
rect 1104 66134 2200 66218
rect 1104 65898 1706 66134
rect 1942 65898 2200 66134
rect 1104 65856 2200 65898
rect 109800 66454 120200 66496
rect 109800 66218 109998 66454
rect 110234 66218 119706 66454
rect 119942 66218 120200 66454
rect 109800 66134 120200 66218
rect 109800 65898 109998 66134
rect 110234 65898 119706 66134
rect 119942 65898 120200 66134
rect 109800 65856 120200 65898
rect 517800 66454 522836 66496
rect 517800 66218 517982 66454
rect 518218 66218 522836 66454
rect 517800 66134 522836 66218
rect 517800 65898 517982 66134
rect 518218 65898 522836 66134
rect 517800 65856 522836 65898
rect 1072 53454 2200 53496
rect 1072 53218 1096 53454
rect 1332 53218 2200 53454
rect 1072 53134 2200 53218
rect 1072 52898 1096 53134
rect 1332 52898 2200 53134
rect 1072 52856 2200 52898
rect 109800 53454 120200 53496
rect 109800 53218 110658 53454
rect 110894 53218 119046 53454
rect 119282 53218 120200 53454
rect 109800 53134 120200 53218
rect 109800 52898 110658 53134
rect 110894 52898 119046 53134
rect 119282 52898 120200 53134
rect 109800 52856 120200 52898
rect 517800 53454 522836 53496
rect 517800 53218 518642 53454
rect 518878 53218 522836 53454
rect 517800 53134 522836 53218
rect 517800 52898 518642 53134
rect 518878 52898 522836 53134
rect 517800 52856 522836 52898
rect 1104 40454 2200 40496
rect 1104 40218 1706 40454
rect 1942 40218 2200 40454
rect 1104 40134 2200 40218
rect 1104 39898 1706 40134
rect 1942 39898 2200 40134
rect 1104 39856 2200 39898
rect 109800 40454 120200 40496
rect 109800 40218 109998 40454
rect 110234 40218 119706 40454
rect 119942 40218 120200 40454
rect 109800 40134 120200 40218
rect 109800 39898 109998 40134
rect 110234 39898 119706 40134
rect 119942 39898 120200 40134
rect 109800 39856 120200 39898
rect 517800 40454 522836 40496
rect 517800 40218 517982 40454
rect 518218 40218 522836 40454
rect 517800 40134 522836 40218
rect 517800 39898 517982 40134
rect 518218 39898 522836 40134
rect 517800 39856 522836 39898
rect 1072 27454 2200 27496
rect 1072 27218 1096 27454
rect 1332 27218 2200 27454
rect 1072 27134 2200 27218
rect 1072 26898 1096 27134
rect 1332 26898 2200 27134
rect 1072 26856 2200 26898
rect 109800 27454 120200 27496
rect 109800 27218 110658 27454
rect 110894 27218 119046 27454
rect 119282 27218 120200 27454
rect 109800 27134 120200 27218
rect 109800 26898 110658 27134
rect 110894 26898 119046 27134
rect 119282 26898 120200 27134
rect 109800 26856 120200 26898
rect 517800 27454 522836 27496
rect 517800 27218 518642 27454
rect 518878 27218 522836 27454
rect 517800 27134 522836 27218
rect 517800 26898 518642 27134
rect 518878 26898 522836 27134
rect 517800 26856 522836 26898
rect 1104 14454 2200 14496
rect 1104 14218 1706 14454
rect 1942 14218 2200 14454
rect 1104 14134 2200 14218
rect 1104 13898 1706 14134
rect 1942 13898 2200 14134
rect 1104 13856 2200 13898
rect 109800 14454 120200 14496
rect 109800 14218 109998 14454
rect 110234 14218 119706 14454
rect 119942 14218 120200 14454
rect 109800 14134 120200 14218
rect 109800 13898 109998 14134
rect 110234 13898 119706 14134
rect 119942 13898 120200 14134
rect 109800 13856 120200 13898
rect 517800 14454 522836 14496
rect 517800 14218 517982 14454
rect 518218 14218 522836 14454
rect 517800 14134 522836 14218
rect 517800 13898 517982 14134
rect 518218 13898 522836 14134
rect 517800 13856 522836 13898
use mgmt_core  core
timestamp 1637331822
transform 1 0 119000 0 1 2000
box 0 0 400000 148000
use DFFRAM  DFFRAM
timestamp 1637331822
transform 1 0 1000 0 1 2000
box 4 0 110000 148000
<< labels >>
rlabel metal5 s 1104 26856 2200 27496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 26856 120200 27496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 26856 522836 27496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 52856 2200 53496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 52856 120200 53496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 52856 522836 53496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 78856 2200 79496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 78856 120200 79496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 78856 522836 79496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 104856 2200 105496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 104856 120200 105496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 104856 522836 105496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 130856 2200 131496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 130856 120200 131496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 130856 522836 131496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 156856 522836 157496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 13856 2200 14496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 13856 120200 14496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 13856 522836 14496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 39856 2200 40496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 39856 120200 40496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 39856 522836 40496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 65856 2200 66496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 65856 120200 66496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 65856 522836 66496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 91856 2200 92496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 91856 120200 92496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 91856 522836 92496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 117856 2200 118496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 117856 120200 118496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 117856 522836 118496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 143856 2200 144496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 143856 120200 144496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 143856 522836 144496 6 VPWR
port 1 nsew power input
rlabel metal2 s 294786 -400 294842 800 6 core_clk
port 2 nsew signal input
rlabel metal2 s 98274 -400 98330 800 6 core_rstn
port 3 nsew signal input
rlabel metal3 s 523200 64472 524400 64592 6 debug_in
port 4 nsew signal input
rlabel metal3 s 523200 65968 524400 66088 6 debug_mode
port 5 nsew signal tristate
rlabel metal3 s 523200 67464 524400 67584 6 debug_oeb
port 6 nsew signal tristate
rlabel metal3 s 523200 68960 524400 69080 6 debug_out
port 7 nsew signal tristate
rlabel metal3 s 523200 144848 524400 144968 6 flash_clk
port 8 nsew signal tristate
rlabel metal3 s 523200 143352 524400 143472 6 flash_csb
port 9 nsew signal tristate
rlabel metal3 s 523200 146480 524400 146600 6 flash_io0_di
port 10 nsew signal input
rlabel metal3 s 523200 147976 524400 148096 6 flash_io0_do
port 11 nsew signal tristate
rlabel metal3 s 523200 149472 524400 149592 6 flash_io0_oeb
port 12 nsew signal tristate
rlabel metal3 s 523200 150968 524400 151088 6 flash_io1_di
port 13 nsew signal input
rlabel metal3 s 523200 152464 524400 152584 6 flash_io1_do
port 14 nsew signal tristate
rlabel metal3 s 523200 153960 524400 154080 6 flash_io1_oeb
port 15 nsew signal tristate
rlabel metal3 s 523200 155592 524400 155712 6 flash_io2_di
port 16 nsew signal input
rlabel metal3 s 523200 157088 524400 157208 6 flash_io2_do
port 17 nsew signal tristate
rlabel metal3 s 523200 158584 524400 158704 6 flash_io2_oeb
port 18 nsew signal tristate
rlabel metal3 s 523200 160080 524400 160200 6 flash_io3_di
port 19 nsew signal input
rlabel metal3 s 523200 161576 524400 161696 6 flash_io3_do
port 20 nsew signal tristate
rlabel metal3 s 523200 163072 524400 163192 6 flash_io3_oeb
port 21 nsew signal tristate
rlabel metal2 s 32770 -400 32826 800 6 gpio_in_pad
port 22 nsew signal input
rlabel metal2 s 163778 -400 163834 800 6 gpio_inenb_pad
port 23 nsew signal tristate
rlabel metal2 s 229282 -400 229338 800 6 gpio_mode0_pad
port 24 nsew signal tristate
rlabel metal2 s 360290 -400 360346 800 6 gpio_mode1_pad
port 25 nsew signal tristate
rlabel metal2 s 425794 -400 425850 800 6 gpio_out_pad
port 26 nsew signal tristate
rlabel metal2 s 491298 -400 491354 800 6 gpio_outenb_pad
port 27 nsew signal tristate
rlabel metal3 s 523200 91808 524400 91928 6 hk_ack_i
port 28 nsew signal input
rlabel metal3 s 523200 94800 524400 94920 6 hk_dat_i[0]
port 29 nsew signal input
rlabel metal3 s 523200 110032 524400 110152 6 hk_dat_i[10]
port 30 nsew signal input
rlabel metal3 s 523200 111528 524400 111648 6 hk_dat_i[11]
port 31 nsew signal input
rlabel metal3 s 523200 113024 524400 113144 6 hk_dat_i[12]
port 32 nsew signal input
rlabel metal3 s 523200 114520 524400 114640 6 hk_dat_i[13]
port 33 nsew signal input
rlabel metal3 s 523200 116016 524400 116136 6 hk_dat_i[14]
port 34 nsew signal input
rlabel metal3 s 523200 117512 524400 117632 6 hk_dat_i[15]
port 35 nsew signal input
rlabel metal3 s 523200 119144 524400 119264 6 hk_dat_i[16]
port 36 nsew signal input
rlabel metal3 s 523200 120640 524400 120760 6 hk_dat_i[17]
port 37 nsew signal input
rlabel metal3 s 523200 122136 524400 122256 6 hk_dat_i[18]
port 38 nsew signal input
rlabel metal3 s 523200 123632 524400 123752 6 hk_dat_i[19]
port 39 nsew signal input
rlabel metal3 s 523200 96296 524400 96416 6 hk_dat_i[1]
port 40 nsew signal input
rlabel metal3 s 523200 125128 524400 125248 6 hk_dat_i[20]
port 41 nsew signal input
rlabel metal3 s 523200 126624 524400 126744 6 hk_dat_i[21]
port 42 nsew signal input
rlabel metal3 s 523200 128256 524400 128376 6 hk_dat_i[22]
port 43 nsew signal input
rlabel metal3 s 523200 129752 524400 129872 6 hk_dat_i[23]
port 44 nsew signal input
rlabel metal3 s 523200 131248 524400 131368 6 hk_dat_i[24]
port 45 nsew signal input
rlabel metal3 s 523200 132744 524400 132864 6 hk_dat_i[25]
port 46 nsew signal input
rlabel metal3 s 523200 134240 524400 134360 6 hk_dat_i[26]
port 47 nsew signal input
rlabel metal3 s 523200 135736 524400 135856 6 hk_dat_i[27]
port 48 nsew signal input
rlabel metal3 s 523200 137368 524400 137488 6 hk_dat_i[28]
port 49 nsew signal input
rlabel metal3 s 523200 138864 524400 138984 6 hk_dat_i[29]
port 50 nsew signal input
rlabel metal3 s 523200 97792 524400 97912 6 hk_dat_i[2]
port 51 nsew signal input
rlabel metal3 s 523200 140360 524400 140480 6 hk_dat_i[30]
port 52 nsew signal input
rlabel metal3 s 523200 141856 524400 141976 6 hk_dat_i[31]
port 53 nsew signal input
rlabel metal3 s 523200 99288 524400 99408 6 hk_dat_i[3]
port 54 nsew signal input
rlabel metal3 s 523200 100920 524400 101040 6 hk_dat_i[4]
port 55 nsew signal input
rlabel metal3 s 523200 102416 524400 102536 6 hk_dat_i[5]
port 56 nsew signal input
rlabel metal3 s 523200 103912 524400 104032 6 hk_dat_i[6]
port 57 nsew signal input
rlabel metal3 s 523200 105408 524400 105528 6 hk_dat_i[7]
port 58 nsew signal input
rlabel metal3 s 523200 106904 524400 107024 6 hk_dat_i[8]
port 59 nsew signal input
rlabel metal3 s 523200 108400 524400 108520 6 hk_dat_i[9]
port 60 nsew signal input
rlabel metal3 s 523200 93304 524400 93424 6 hk_stb_o
port 61 nsew signal tristate
rlabel metal2 s 521842 163200 521898 164400 6 irq[0]
port 62 nsew signal input
rlabel metal2 s 522670 163200 522726 164400 6 irq[1]
port 63 nsew signal input
rlabel metal2 s 523498 163200 523554 164400 6 irq[2]
port 64 nsew signal input
rlabel metal3 s 523200 75080 524400 75200 6 irq[3]
port 65 nsew signal input
rlabel metal3 s 523200 73584 524400 73704 6 irq[4]
port 66 nsew signal input
rlabel metal3 s 523200 71952 524400 72072 6 irq[5]
port 67 nsew signal input
rlabel metal2 s 386 163200 442 164400 6 la_iena[0]
port 68 nsew signal tristate
rlabel metal2 s 336830 163200 336886 164400 6 la_iena[100]
port 69 nsew signal tristate
rlabel metal2 s 340142 163200 340198 164400 6 la_iena[101]
port 70 nsew signal tristate
rlabel metal2 s 343546 163200 343602 164400 6 la_iena[102]
port 71 nsew signal tristate
rlabel metal2 s 346858 163200 346914 164400 6 la_iena[103]
port 72 nsew signal tristate
rlabel metal2 s 350262 163200 350318 164400 6 la_iena[104]
port 73 nsew signal tristate
rlabel metal2 s 353666 163200 353722 164400 6 la_iena[105]
port 74 nsew signal tristate
rlabel metal2 s 356978 163200 357034 164400 6 la_iena[106]
port 75 nsew signal tristate
rlabel metal2 s 360382 163200 360438 164400 6 la_iena[107]
port 76 nsew signal tristate
rlabel metal2 s 363694 163200 363750 164400 6 la_iena[108]
port 77 nsew signal tristate
rlabel metal2 s 367098 163200 367154 164400 6 la_iena[109]
port 78 nsew signal tristate
rlabel metal2 s 33966 163200 34022 164400 6 la_iena[10]
port 79 nsew signal tristate
rlabel metal2 s 370410 163200 370466 164400 6 la_iena[110]
port 80 nsew signal tristate
rlabel metal2 s 373814 163200 373870 164400 6 la_iena[111]
port 81 nsew signal tristate
rlabel metal2 s 377218 163200 377274 164400 6 la_iena[112]
port 82 nsew signal tristate
rlabel metal2 s 380530 163200 380586 164400 6 la_iena[113]
port 83 nsew signal tristate
rlabel metal2 s 383934 163200 383990 164400 6 la_iena[114]
port 84 nsew signal tristate
rlabel metal2 s 387246 163200 387302 164400 6 la_iena[115]
port 85 nsew signal tristate
rlabel metal2 s 390650 163200 390706 164400 6 la_iena[116]
port 86 nsew signal tristate
rlabel metal2 s 393962 163200 394018 164400 6 la_iena[117]
port 87 nsew signal tristate
rlabel metal2 s 397366 163200 397422 164400 6 la_iena[118]
port 88 nsew signal tristate
rlabel metal2 s 400770 163200 400826 164400 6 la_iena[119]
port 89 nsew signal tristate
rlabel metal2 s 37370 163200 37426 164400 6 la_iena[11]
port 90 nsew signal tristate
rlabel metal2 s 404082 163200 404138 164400 6 la_iena[120]
port 91 nsew signal tristate
rlabel metal2 s 407486 163200 407542 164400 6 la_iena[121]
port 92 nsew signal tristate
rlabel metal2 s 410798 163200 410854 164400 6 la_iena[122]
port 93 nsew signal tristate
rlabel metal2 s 414202 163200 414258 164400 6 la_iena[123]
port 94 nsew signal tristate
rlabel metal2 s 417514 163200 417570 164400 6 la_iena[124]
port 95 nsew signal tristate
rlabel metal2 s 420918 163200 420974 164400 6 la_iena[125]
port 96 nsew signal tristate
rlabel metal2 s 424322 163200 424378 164400 6 la_iena[126]
port 97 nsew signal tristate
rlabel metal2 s 427634 163200 427690 164400 6 la_iena[127]
port 98 nsew signal tristate
rlabel metal2 s 40682 163200 40738 164400 6 la_iena[12]
port 99 nsew signal tristate
rlabel metal2 s 44086 163200 44142 164400 6 la_iena[13]
port 100 nsew signal tristate
rlabel metal2 s 47490 163200 47546 164400 6 la_iena[14]
port 101 nsew signal tristate
rlabel metal2 s 50802 163200 50858 164400 6 la_iena[15]
port 102 nsew signal tristate
rlabel metal2 s 54206 163200 54262 164400 6 la_iena[16]
port 103 nsew signal tristate
rlabel metal2 s 57518 163200 57574 164400 6 la_iena[17]
port 104 nsew signal tristate
rlabel metal2 s 60922 163200 60978 164400 6 la_iena[18]
port 105 nsew signal tristate
rlabel metal2 s 64234 163200 64290 164400 6 la_iena[19]
port 106 nsew signal tristate
rlabel metal2 s 3698 163200 3754 164400 6 la_iena[1]
port 107 nsew signal tristate
rlabel metal2 s 67638 163200 67694 164400 6 la_iena[20]
port 108 nsew signal tristate
rlabel metal2 s 71042 163200 71098 164400 6 la_iena[21]
port 109 nsew signal tristate
rlabel metal2 s 74354 163200 74410 164400 6 la_iena[22]
port 110 nsew signal tristate
rlabel metal2 s 77758 163200 77814 164400 6 la_iena[23]
port 111 nsew signal tristate
rlabel metal2 s 81070 163200 81126 164400 6 la_iena[24]
port 112 nsew signal tristate
rlabel metal2 s 84474 163200 84530 164400 6 la_iena[25]
port 113 nsew signal tristate
rlabel metal2 s 87786 163200 87842 164400 6 la_iena[26]
port 114 nsew signal tristate
rlabel metal2 s 91190 163200 91246 164400 6 la_iena[27]
port 115 nsew signal tristate
rlabel metal2 s 94594 163200 94650 164400 6 la_iena[28]
port 116 nsew signal tristate
rlabel metal2 s 97906 163200 97962 164400 6 la_iena[29]
port 117 nsew signal tristate
rlabel metal2 s 7102 163200 7158 164400 6 la_iena[2]
port 118 nsew signal tristate
rlabel metal2 s 101310 163200 101366 164400 6 la_iena[30]
port 119 nsew signal tristate
rlabel metal2 s 104622 163200 104678 164400 6 la_iena[31]
port 120 nsew signal tristate
rlabel metal2 s 108026 163200 108082 164400 6 la_iena[32]
port 121 nsew signal tristate
rlabel metal2 s 111338 163200 111394 164400 6 la_iena[33]
port 122 nsew signal tristate
rlabel metal2 s 114742 163200 114798 164400 6 la_iena[34]
port 123 nsew signal tristate
rlabel metal2 s 118146 163200 118202 164400 6 la_iena[35]
port 124 nsew signal tristate
rlabel metal2 s 121458 163200 121514 164400 6 la_iena[36]
port 125 nsew signal tristate
rlabel metal2 s 124862 163200 124918 164400 6 la_iena[37]
port 126 nsew signal tristate
rlabel metal2 s 128174 163200 128230 164400 6 la_iena[38]
port 127 nsew signal tristate
rlabel metal2 s 131578 163200 131634 164400 6 la_iena[39]
port 128 nsew signal tristate
rlabel metal2 s 10414 163200 10470 164400 6 la_iena[3]
port 129 nsew signal tristate
rlabel metal2 s 134890 163200 134946 164400 6 la_iena[40]
port 130 nsew signal tristate
rlabel metal2 s 138294 163200 138350 164400 6 la_iena[41]
port 131 nsew signal tristate
rlabel metal2 s 141698 163200 141754 164400 6 la_iena[42]
port 132 nsew signal tristate
rlabel metal2 s 145010 163200 145066 164400 6 la_iena[43]
port 133 nsew signal tristate
rlabel metal2 s 148414 163200 148470 164400 6 la_iena[44]
port 134 nsew signal tristate
rlabel metal2 s 151726 163200 151782 164400 6 la_iena[45]
port 135 nsew signal tristate
rlabel metal2 s 155130 163200 155186 164400 6 la_iena[46]
port 136 nsew signal tristate
rlabel metal2 s 158442 163200 158498 164400 6 la_iena[47]
port 137 nsew signal tristate
rlabel metal2 s 161846 163200 161902 164400 6 la_iena[48]
port 138 nsew signal tristate
rlabel metal2 s 165250 163200 165306 164400 6 la_iena[49]
port 139 nsew signal tristate
rlabel metal2 s 13818 163200 13874 164400 6 la_iena[4]
port 140 nsew signal tristate
rlabel metal2 s 168562 163200 168618 164400 6 la_iena[50]
port 141 nsew signal tristate
rlabel metal2 s 171966 163200 172022 164400 6 la_iena[51]
port 142 nsew signal tristate
rlabel metal2 s 175278 163200 175334 164400 6 la_iena[52]
port 143 nsew signal tristate
rlabel metal2 s 178682 163200 178738 164400 6 la_iena[53]
port 144 nsew signal tristate
rlabel metal2 s 181994 163200 182050 164400 6 la_iena[54]
port 145 nsew signal tristate
rlabel metal2 s 185398 163200 185454 164400 6 la_iena[55]
port 146 nsew signal tristate
rlabel metal2 s 188802 163200 188858 164400 6 la_iena[56]
port 147 nsew signal tristate
rlabel metal2 s 192114 163200 192170 164400 6 la_iena[57]
port 148 nsew signal tristate
rlabel metal2 s 195518 163200 195574 164400 6 la_iena[58]
port 149 nsew signal tristate
rlabel metal2 s 198830 163200 198886 164400 6 la_iena[59]
port 150 nsew signal tristate
rlabel metal2 s 17130 163200 17186 164400 6 la_iena[5]
port 151 nsew signal tristate
rlabel metal2 s 202234 163200 202290 164400 6 la_iena[60]
port 152 nsew signal tristate
rlabel metal2 s 205546 163200 205602 164400 6 la_iena[61]
port 153 nsew signal tristate
rlabel metal2 s 208950 163200 209006 164400 6 la_iena[62]
port 154 nsew signal tristate
rlabel metal2 s 212354 163200 212410 164400 6 la_iena[63]
port 155 nsew signal tristate
rlabel metal2 s 215666 163200 215722 164400 6 la_iena[64]
port 156 nsew signal tristate
rlabel metal2 s 219070 163200 219126 164400 6 la_iena[65]
port 157 nsew signal tristate
rlabel metal2 s 222382 163200 222438 164400 6 la_iena[66]
port 158 nsew signal tristate
rlabel metal2 s 225786 163200 225842 164400 6 la_iena[67]
port 159 nsew signal tristate
rlabel metal2 s 229098 163200 229154 164400 6 la_iena[68]
port 160 nsew signal tristate
rlabel metal2 s 232502 163200 232558 164400 6 la_iena[69]
port 161 nsew signal tristate
rlabel metal2 s 20534 163200 20590 164400 6 la_iena[6]
port 162 nsew signal tristate
rlabel metal2 s 235906 163200 235962 164400 6 la_iena[70]
port 163 nsew signal tristate
rlabel metal2 s 239218 163200 239274 164400 6 la_iena[71]
port 164 nsew signal tristate
rlabel metal2 s 242622 163200 242678 164400 6 la_iena[72]
port 165 nsew signal tristate
rlabel metal2 s 245934 163200 245990 164400 6 la_iena[73]
port 166 nsew signal tristate
rlabel metal2 s 249338 163200 249394 164400 6 la_iena[74]
port 167 nsew signal tristate
rlabel metal2 s 252650 163200 252706 164400 6 la_iena[75]
port 168 nsew signal tristate
rlabel metal2 s 256054 163200 256110 164400 6 la_iena[76]
port 169 nsew signal tristate
rlabel metal2 s 259458 163200 259514 164400 6 la_iena[77]
port 170 nsew signal tristate
rlabel metal2 s 262770 163200 262826 164400 6 la_iena[78]
port 171 nsew signal tristate
rlabel metal2 s 266174 163200 266230 164400 6 la_iena[79]
port 172 nsew signal tristate
rlabel metal2 s 23938 163200 23994 164400 6 la_iena[7]
port 173 nsew signal tristate
rlabel metal2 s 269486 163200 269542 164400 6 la_iena[80]
port 174 nsew signal tristate
rlabel metal2 s 272890 163200 272946 164400 6 la_iena[81]
port 175 nsew signal tristate
rlabel metal2 s 276202 163200 276258 164400 6 la_iena[82]
port 176 nsew signal tristate
rlabel metal2 s 279606 163200 279662 164400 6 la_iena[83]
port 177 nsew signal tristate
rlabel metal2 s 283010 163200 283066 164400 6 la_iena[84]
port 178 nsew signal tristate
rlabel metal2 s 286322 163200 286378 164400 6 la_iena[85]
port 179 nsew signal tristate
rlabel metal2 s 289726 163200 289782 164400 6 la_iena[86]
port 180 nsew signal tristate
rlabel metal2 s 293038 163200 293094 164400 6 la_iena[87]
port 181 nsew signal tristate
rlabel metal2 s 296442 163200 296498 164400 6 la_iena[88]
port 182 nsew signal tristate
rlabel metal2 s 299754 163200 299810 164400 6 la_iena[89]
port 183 nsew signal tristate
rlabel metal2 s 27250 163200 27306 164400 6 la_iena[8]
port 184 nsew signal tristate
rlabel metal2 s 303158 163200 303214 164400 6 la_iena[90]
port 185 nsew signal tristate
rlabel metal2 s 306562 163200 306618 164400 6 la_iena[91]
port 186 nsew signal tristate
rlabel metal2 s 309874 163200 309930 164400 6 la_iena[92]
port 187 nsew signal tristate
rlabel metal2 s 313278 163200 313334 164400 6 la_iena[93]
port 188 nsew signal tristate
rlabel metal2 s 316590 163200 316646 164400 6 la_iena[94]
port 189 nsew signal tristate
rlabel metal2 s 319994 163200 320050 164400 6 la_iena[95]
port 190 nsew signal tristate
rlabel metal2 s 323306 163200 323362 164400 6 la_iena[96]
port 191 nsew signal tristate
rlabel metal2 s 326710 163200 326766 164400 6 la_iena[97]
port 192 nsew signal tristate
rlabel metal2 s 330114 163200 330170 164400 6 la_iena[98]
port 193 nsew signal tristate
rlabel metal2 s 333426 163200 333482 164400 6 la_iena[99]
port 194 nsew signal tristate
rlabel metal2 s 30654 163200 30710 164400 6 la_iena[9]
port 195 nsew signal tristate
rlabel metal2 s 1214 163200 1270 164400 6 la_input[0]
port 196 nsew signal input
rlabel metal2 s 337658 163200 337714 164400 6 la_input[100]
port 197 nsew signal input
rlabel metal2 s 340970 163200 341026 164400 6 la_input[101]
port 198 nsew signal input
rlabel metal2 s 344374 163200 344430 164400 6 la_input[102]
port 199 nsew signal input
rlabel metal2 s 347778 163200 347834 164400 6 la_input[103]
port 200 nsew signal input
rlabel metal2 s 351090 163200 351146 164400 6 la_input[104]
port 201 nsew signal input
rlabel metal2 s 354494 163200 354550 164400 6 la_input[105]
port 202 nsew signal input
rlabel metal2 s 357806 163200 357862 164400 6 la_input[106]
port 203 nsew signal input
rlabel metal2 s 361210 163200 361266 164400 6 la_input[107]
port 204 nsew signal input
rlabel metal2 s 364522 163200 364578 164400 6 la_input[108]
port 205 nsew signal input
rlabel metal2 s 367926 163200 367982 164400 6 la_input[109]
port 206 nsew signal input
rlabel metal2 s 34794 163200 34850 164400 6 la_input[10]
port 207 nsew signal input
rlabel metal2 s 371330 163200 371386 164400 6 la_input[110]
port 208 nsew signal input
rlabel metal2 s 374642 163200 374698 164400 6 la_input[111]
port 209 nsew signal input
rlabel metal2 s 378046 163200 378102 164400 6 la_input[112]
port 210 nsew signal input
rlabel metal2 s 381358 163200 381414 164400 6 la_input[113]
port 211 nsew signal input
rlabel metal2 s 384762 163200 384818 164400 6 la_input[114]
port 212 nsew signal input
rlabel metal2 s 388074 163200 388130 164400 6 la_input[115]
port 213 nsew signal input
rlabel metal2 s 391478 163200 391534 164400 6 la_input[116]
port 214 nsew signal input
rlabel metal2 s 394882 163200 394938 164400 6 la_input[117]
port 215 nsew signal input
rlabel metal2 s 398194 163200 398250 164400 6 la_input[118]
port 216 nsew signal input
rlabel metal2 s 401598 163200 401654 164400 6 la_input[119]
port 217 nsew signal input
rlabel metal2 s 38198 163200 38254 164400 6 la_input[11]
port 218 nsew signal input
rlabel metal2 s 404910 163200 404966 164400 6 la_input[120]
port 219 nsew signal input
rlabel metal2 s 408314 163200 408370 164400 6 la_input[121]
port 220 nsew signal input
rlabel metal2 s 411626 163200 411682 164400 6 la_input[122]
port 221 nsew signal input
rlabel metal2 s 415030 163200 415086 164400 6 la_input[123]
port 222 nsew signal input
rlabel metal2 s 418434 163200 418490 164400 6 la_input[124]
port 223 nsew signal input
rlabel metal2 s 421746 163200 421802 164400 6 la_input[125]
port 224 nsew signal input
rlabel metal2 s 425150 163200 425206 164400 6 la_input[126]
port 225 nsew signal input
rlabel metal2 s 428462 163200 428518 164400 6 la_input[127]
port 226 nsew signal input
rlabel metal2 s 41602 163200 41658 164400 6 la_input[12]
port 227 nsew signal input
rlabel metal2 s 44914 163200 44970 164400 6 la_input[13]
port 228 nsew signal input
rlabel metal2 s 48318 163200 48374 164400 6 la_input[14]
port 229 nsew signal input
rlabel metal2 s 51630 163200 51686 164400 6 la_input[15]
port 230 nsew signal input
rlabel metal2 s 55034 163200 55090 164400 6 la_input[16]
port 231 nsew signal input
rlabel metal2 s 58346 163200 58402 164400 6 la_input[17]
port 232 nsew signal input
rlabel metal2 s 61750 163200 61806 164400 6 la_input[18]
port 233 nsew signal input
rlabel metal2 s 65154 163200 65210 164400 6 la_input[19]
port 234 nsew signal input
rlabel metal2 s 4526 163200 4582 164400 6 la_input[1]
port 235 nsew signal input
rlabel metal2 s 68466 163200 68522 164400 6 la_input[20]
port 236 nsew signal input
rlabel metal2 s 71870 163200 71926 164400 6 la_input[21]
port 237 nsew signal input
rlabel metal2 s 75182 163200 75238 164400 6 la_input[22]
port 238 nsew signal input
rlabel metal2 s 78586 163200 78642 164400 6 la_input[23]
port 239 nsew signal input
rlabel metal2 s 81898 163200 81954 164400 6 la_input[24]
port 240 nsew signal input
rlabel metal2 s 85302 163200 85358 164400 6 la_input[25]
port 241 nsew signal input
rlabel metal2 s 88706 163200 88762 164400 6 la_input[26]
port 242 nsew signal input
rlabel metal2 s 92018 163200 92074 164400 6 la_input[27]
port 243 nsew signal input
rlabel metal2 s 95422 163200 95478 164400 6 la_input[28]
port 244 nsew signal input
rlabel metal2 s 98734 163200 98790 164400 6 la_input[29]
port 245 nsew signal input
rlabel metal2 s 7930 163200 7986 164400 6 la_input[2]
port 246 nsew signal input
rlabel metal2 s 102138 163200 102194 164400 6 la_input[30]
port 247 nsew signal input
rlabel metal2 s 105450 163200 105506 164400 6 la_input[31]
port 248 nsew signal input
rlabel metal2 s 108854 163200 108910 164400 6 la_input[32]
port 249 nsew signal input
rlabel metal2 s 112258 163200 112314 164400 6 la_input[33]
port 250 nsew signal input
rlabel metal2 s 115570 163200 115626 164400 6 la_input[34]
port 251 nsew signal input
rlabel metal2 s 118974 163200 119030 164400 6 la_input[35]
port 252 nsew signal input
rlabel metal2 s 122286 163200 122342 164400 6 la_input[36]
port 253 nsew signal input
rlabel metal2 s 125690 163200 125746 164400 6 la_input[37]
port 254 nsew signal input
rlabel metal2 s 129002 163200 129058 164400 6 la_input[38]
port 255 nsew signal input
rlabel metal2 s 132406 163200 132462 164400 6 la_input[39]
port 256 nsew signal input
rlabel metal2 s 11242 163200 11298 164400 6 la_input[3]
port 257 nsew signal input
rlabel metal2 s 135810 163200 135866 164400 6 la_input[40]
port 258 nsew signal input
rlabel metal2 s 139122 163200 139178 164400 6 la_input[41]
port 259 nsew signal input
rlabel metal2 s 142526 163200 142582 164400 6 la_input[42]
port 260 nsew signal input
rlabel metal2 s 145838 163200 145894 164400 6 la_input[43]
port 261 nsew signal input
rlabel metal2 s 149242 163200 149298 164400 6 la_input[44]
port 262 nsew signal input
rlabel metal2 s 152554 163200 152610 164400 6 la_input[45]
port 263 nsew signal input
rlabel metal2 s 155958 163200 156014 164400 6 la_input[46]
port 264 nsew signal input
rlabel metal2 s 159362 163200 159418 164400 6 la_input[47]
port 265 nsew signal input
rlabel metal2 s 162674 163200 162730 164400 6 la_input[48]
port 266 nsew signal input
rlabel metal2 s 166078 163200 166134 164400 6 la_input[49]
port 267 nsew signal input
rlabel metal2 s 14646 163200 14702 164400 6 la_input[4]
port 268 nsew signal input
rlabel metal2 s 169390 163200 169446 164400 6 la_input[50]
port 269 nsew signal input
rlabel metal2 s 172794 163200 172850 164400 6 la_input[51]
port 270 nsew signal input
rlabel metal2 s 176106 163200 176162 164400 6 la_input[52]
port 271 nsew signal input
rlabel metal2 s 179510 163200 179566 164400 6 la_input[53]
port 272 nsew signal input
rlabel metal2 s 182914 163200 182970 164400 6 la_input[54]
port 273 nsew signal input
rlabel metal2 s 186226 163200 186282 164400 6 la_input[55]
port 274 nsew signal input
rlabel metal2 s 189630 163200 189686 164400 6 la_input[56]
port 275 nsew signal input
rlabel metal2 s 192942 163200 192998 164400 6 la_input[57]
port 276 nsew signal input
rlabel metal2 s 196346 163200 196402 164400 6 la_input[58]
port 277 nsew signal input
rlabel metal2 s 199658 163200 199714 164400 6 la_input[59]
port 278 nsew signal input
rlabel metal2 s 18050 163200 18106 164400 6 la_input[5]
port 279 nsew signal input
rlabel metal2 s 203062 163200 203118 164400 6 la_input[60]
port 280 nsew signal input
rlabel metal2 s 206466 163200 206522 164400 6 la_input[61]
port 281 nsew signal input
rlabel metal2 s 209778 163200 209834 164400 6 la_input[62]
port 282 nsew signal input
rlabel metal2 s 213182 163200 213238 164400 6 la_input[63]
port 283 nsew signal input
rlabel metal2 s 216494 163200 216550 164400 6 la_input[64]
port 284 nsew signal input
rlabel metal2 s 219898 163200 219954 164400 6 la_input[65]
port 285 nsew signal input
rlabel metal2 s 223210 163200 223266 164400 6 la_input[66]
port 286 nsew signal input
rlabel metal2 s 226614 163200 226670 164400 6 la_input[67]
port 287 nsew signal input
rlabel metal2 s 230018 163200 230074 164400 6 la_input[68]
port 288 nsew signal input
rlabel metal2 s 233330 163200 233386 164400 6 la_input[69]
port 289 nsew signal input
rlabel metal2 s 21362 163200 21418 164400 6 la_input[6]
port 290 nsew signal input
rlabel metal2 s 236734 163200 236790 164400 6 la_input[70]
port 291 nsew signal input
rlabel metal2 s 240046 163200 240102 164400 6 la_input[71]
port 292 nsew signal input
rlabel metal2 s 243450 163200 243506 164400 6 la_input[72]
port 293 nsew signal input
rlabel metal2 s 246762 163200 246818 164400 6 la_input[73]
port 294 nsew signal input
rlabel metal2 s 250166 163200 250222 164400 6 la_input[74]
port 295 nsew signal input
rlabel metal2 s 253570 163200 253626 164400 6 la_input[75]
port 296 nsew signal input
rlabel metal2 s 256882 163200 256938 164400 6 la_input[76]
port 297 nsew signal input
rlabel metal2 s 260286 163200 260342 164400 6 la_input[77]
port 298 nsew signal input
rlabel metal2 s 263598 163200 263654 164400 6 la_input[78]
port 299 nsew signal input
rlabel metal2 s 267002 163200 267058 164400 6 la_input[79]
port 300 nsew signal input
rlabel metal2 s 24766 163200 24822 164400 6 la_input[7]
port 301 nsew signal input
rlabel metal2 s 270314 163200 270370 164400 6 la_input[80]
port 302 nsew signal input
rlabel metal2 s 273718 163200 273774 164400 6 la_input[81]
port 303 nsew signal input
rlabel metal2 s 277122 163200 277178 164400 6 la_input[82]
port 304 nsew signal input
rlabel metal2 s 280434 163200 280490 164400 6 la_input[83]
port 305 nsew signal input
rlabel metal2 s 283838 163200 283894 164400 6 la_input[84]
port 306 nsew signal input
rlabel metal2 s 287150 163200 287206 164400 6 la_input[85]
port 307 nsew signal input
rlabel metal2 s 290554 163200 290610 164400 6 la_input[86]
port 308 nsew signal input
rlabel metal2 s 293866 163200 293922 164400 6 la_input[87]
port 309 nsew signal input
rlabel metal2 s 297270 163200 297326 164400 6 la_input[88]
port 310 nsew signal input
rlabel metal2 s 300674 163200 300730 164400 6 la_input[89]
port 311 nsew signal input
rlabel metal2 s 28078 163200 28134 164400 6 la_input[8]
port 312 nsew signal input
rlabel metal2 s 303986 163200 304042 164400 6 la_input[90]
port 313 nsew signal input
rlabel metal2 s 307390 163200 307446 164400 6 la_input[91]
port 314 nsew signal input
rlabel metal2 s 310702 163200 310758 164400 6 la_input[92]
port 315 nsew signal input
rlabel metal2 s 314106 163200 314162 164400 6 la_input[93]
port 316 nsew signal input
rlabel metal2 s 317418 163200 317474 164400 6 la_input[94]
port 317 nsew signal input
rlabel metal2 s 320822 163200 320878 164400 6 la_input[95]
port 318 nsew signal input
rlabel metal2 s 324226 163200 324282 164400 6 la_input[96]
port 319 nsew signal input
rlabel metal2 s 327538 163200 327594 164400 6 la_input[97]
port 320 nsew signal input
rlabel metal2 s 330942 163200 330998 164400 6 la_input[98]
port 321 nsew signal input
rlabel metal2 s 334254 163200 334310 164400 6 la_input[99]
port 322 nsew signal input
rlabel metal2 s 31482 163200 31538 164400 6 la_input[9]
port 323 nsew signal input
rlabel metal2 s 2042 163200 2098 164400 6 la_oenb[0]
port 324 nsew signal tristate
rlabel metal2 s 338486 163200 338542 164400 6 la_oenb[100]
port 325 nsew signal tristate
rlabel metal2 s 341890 163200 341946 164400 6 la_oenb[101]
port 326 nsew signal tristate
rlabel metal2 s 345202 163200 345258 164400 6 la_oenb[102]
port 327 nsew signal tristate
rlabel metal2 s 348606 163200 348662 164400 6 la_oenb[103]
port 328 nsew signal tristate
rlabel metal2 s 351918 163200 351974 164400 6 la_oenb[104]
port 329 nsew signal tristate
rlabel metal2 s 355322 163200 355378 164400 6 la_oenb[105]
port 330 nsew signal tristate
rlabel metal2 s 358634 163200 358690 164400 6 la_oenb[106]
port 331 nsew signal tristate
rlabel metal2 s 362038 163200 362094 164400 6 la_oenb[107]
port 332 nsew signal tristate
rlabel metal2 s 365442 163200 365498 164400 6 la_oenb[108]
port 333 nsew signal tristate
rlabel metal2 s 368754 163200 368810 164400 6 la_oenb[109]
port 334 nsew signal tristate
rlabel metal2 s 35714 163200 35770 164400 6 la_oenb[10]
port 335 nsew signal tristate
rlabel metal2 s 372158 163200 372214 164400 6 la_oenb[110]
port 336 nsew signal tristate
rlabel metal2 s 375470 163200 375526 164400 6 la_oenb[111]
port 337 nsew signal tristate
rlabel metal2 s 378874 163200 378930 164400 6 la_oenb[112]
port 338 nsew signal tristate
rlabel metal2 s 382186 163200 382242 164400 6 la_oenb[113]
port 339 nsew signal tristate
rlabel metal2 s 385590 163200 385646 164400 6 la_oenb[114]
port 340 nsew signal tristate
rlabel metal2 s 388994 163200 389050 164400 6 la_oenb[115]
port 341 nsew signal tristate
rlabel metal2 s 392306 163200 392362 164400 6 la_oenb[116]
port 342 nsew signal tristate
rlabel metal2 s 395710 163200 395766 164400 6 la_oenb[117]
port 343 nsew signal tristate
rlabel metal2 s 399022 163200 399078 164400 6 la_oenb[118]
port 344 nsew signal tristate
rlabel metal2 s 402426 163200 402482 164400 6 la_oenb[119]
port 345 nsew signal tristate
rlabel metal2 s 39026 163200 39082 164400 6 la_oenb[11]
port 346 nsew signal tristate
rlabel metal2 s 405738 163200 405794 164400 6 la_oenb[120]
port 347 nsew signal tristate
rlabel metal2 s 409142 163200 409198 164400 6 la_oenb[121]
port 348 nsew signal tristate
rlabel metal2 s 412546 163200 412602 164400 6 la_oenb[122]
port 349 nsew signal tristate
rlabel metal2 s 415858 163200 415914 164400 6 la_oenb[123]
port 350 nsew signal tristate
rlabel metal2 s 419262 163200 419318 164400 6 la_oenb[124]
port 351 nsew signal tristate
rlabel metal2 s 422574 163200 422630 164400 6 la_oenb[125]
port 352 nsew signal tristate
rlabel metal2 s 425978 163200 426034 164400 6 la_oenb[126]
port 353 nsew signal tristate
rlabel metal2 s 429290 163200 429346 164400 6 la_oenb[127]
port 354 nsew signal tristate
rlabel metal2 s 42430 163200 42486 164400 6 la_oenb[12]
port 355 nsew signal tristate
rlabel metal2 s 45742 163200 45798 164400 6 la_oenb[13]
port 356 nsew signal tristate
rlabel metal2 s 49146 163200 49202 164400 6 la_oenb[14]
port 357 nsew signal tristate
rlabel metal2 s 52458 163200 52514 164400 6 la_oenb[15]
port 358 nsew signal tristate
rlabel metal2 s 55862 163200 55918 164400 6 la_oenb[16]
port 359 nsew signal tristate
rlabel metal2 s 59266 163200 59322 164400 6 la_oenb[17]
port 360 nsew signal tristate
rlabel metal2 s 62578 163200 62634 164400 6 la_oenb[18]
port 361 nsew signal tristate
rlabel metal2 s 65982 163200 66038 164400 6 la_oenb[19]
port 362 nsew signal tristate
rlabel metal2 s 5354 163200 5410 164400 6 la_oenb[1]
port 363 nsew signal tristate
rlabel metal2 s 69294 163200 69350 164400 6 la_oenb[20]
port 364 nsew signal tristate
rlabel metal2 s 72698 163200 72754 164400 6 la_oenb[21]
port 365 nsew signal tristate
rlabel metal2 s 76010 163200 76066 164400 6 la_oenb[22]
port 366 nsew signal tristate
rlabel metal2 s 79414 163200 79470 164400 6 la_oenb[23]
port 367 nsew signal tristate
rlabel metal2 s 82818 163200 82874 164400 6 la_oenb[24]
port 368 nsew signal tristate
rlabel metal2 s 86130 163200 86186 164400 6 la_oenb[25]
port 369 nsew signal tristate
rlabel metal2 s 89534 163200 89590 164400 6 la_oenb[26]
port 370 nsew signal tristate
rlabel metal2 s 92846 163200 92902 164400 6 la_oenb[27]
port 371 nsew signal tristate
rlabel metal2 s 96250 163200 96306 164400 6 la_oenb[28]
port 372 nsew signal tristate
rlabel metal2 s 99562 163200 99618 164400 6 la_oenb[29]
port 373 nsew signal tristate
rlabel metal2 s 8758 163200 8814 164400 6 la_oenb[2]
port 374 nsew signal tristate
rlabel metal2 s 102966 163200 103022 164400 6 la_oenb[30]
port 375 nsew signal tristate
rlabel metal2 s 106370 163200 106426 164400 6 la_oenb[31]
port 376 nsew signal tristate
rlabel metal2 s 109682 163200 109738 164400 6 la_oenb[32]
port 377 nsew signal tristate
rlabel metal2 s 113086 163200 113142 164400 6 la_oenb[33]
port 378 nsew signal tristate
rlabel metal2 s 116398 163200 116454 164400 6 la_oenb[34]
port 379 nsew signal tristate
rlabel metal2 s 119802 163200 119858 164400 6 la_oenb[35]
port 380 nsew signal tristate
rlabel metal2 s 123114 163200 123170 164400 6 la_oenb[36]
port 381 nsew signal tristate
rlabel metal2 s 126518 163200 126574 164400 6 la_oenb[37]
port 382 nsew signal tristate
rlabel metal2 s 129922 163200 129978 164400 6 la_oenb[38]
port 383 nsew signal tristate
rlabel metal2 s 133234 163200 133290 164400 6 la_oenb[39]
port 384 nsew signal tristate
rlabel metal2 s 12162 163200 12218 164400 6 la_oenb[3]
port 385 nsew signal tristate
rlabel metal2 s 136638 163200 136694 164400 6 la_oenb[40]
port 386 nsew signal tristate
rlabel metal2 s 139950 163200 140006 164400 6 la_oenb[41]
port 387 nsew signal tristate
rlabel metal2 s 143354 163200 143410 164400 6 la_oenb[42]
port 388 nsew signal tristate
rlabel metal2 s 146666 163200 146722 164400 6 la_oenb[43]
port 389 nsew signal tristate
rlabel metal2 s 150070 163200 150126 164400 6 la_oenb[44]
port 390 nsew signal tristate
rlabel metal2 s 153474 163200 153530 164400 6 la_oenb[45]
port 391 nsew signal tristate
rlabel metal2 s 156786 163200 156842 164400 6 la_oenb[46]
port 392 nsew signal tristate
rlabel metal2 s 160190 163200 160246 164400 6 la_oenb[47]
port 393 nsew signal tristate
rlabel metal2 s 163502 163200 163558 164400 6 la_oenb[48]
port 394 nsew signal tristate
rlabel metal2 s 166906 163200 166962 164400 6 la_oenb[49]
port 395 nsew signal tristate
rlabel metal2 s 15474 163200 15530 164400 6 la_oenb[4]
port 396 nsew signal tristate
rlabel metal2 s 170218 163200 170274 164400 6 la_oenb[50]
port 397 nsew signal tristate
rlabel metal2 s 173622 163200 173678 164400 6 la_oenb[51]
port 398 nsew signal tristate
rlabel metal2 s 177026 163200 177082 164400 6 la_oenb[52]
port 399 nsew signal tristate
rlabel metal2 s 180338 163200 180394 164400 6 la_oenb[53]
port 400 nsew signal tristate
rlabel metal2 s 183742 163200 183798 164400 6 la_oenb[54]
port 401 nsew signal tristate
rlabel metal2 s 187054 163200 187110 164400 6 la_oenb[55]
port 402 nsew signal tristate
rlabel metal2 s 190458 163200 190514 164400 6 la_oenb[56]
port 403 nsew signal tristate
rlabel metal2 s 193770 163200 193826 164400 6 la_oenb[57]
port 404 nsew signal tristate
rlabel metal2 s 197174 163200 197230 164400 6 la_oenb[58]
port 405 nsew signal tristate
rlabel metal2 s 200578 163200 200634 164400 6 la_oenb[59]
port 406 nsew signal tristate
rlabel metal2 s 18878 163200 18934 164400 6 la_oenb[5]
port 407 nsew signal tristate
rlabel metal2 s 203890 163200 203946 164400 6 la_oenb[60]
port 408 nsew signal tristate
rlabel metal2 s 207294 163200 207350 164400 6 la_oenb[61]
port 409 nsew signal tristate
rlabel metal2 s 210606 163200 210662 164400 6 la_oenb[62]
port 410 nsew signal tristate
rlabel metal2 s 214010 163200 214066 164400 6 la_oenb[63]
port 411 nsew signal tristate
rlabel metal2 s 217322 163200 217378 164400 6 la_oenb[64]
port 412 nsew signal tristate
rlabel metal2 s 220726 163200 220782 164400 6 la_oenb[65]
port 413 nsew signal tristate
rlabel metal2 s 224130 163200 224186 164400 6 la_oenb[66]
port 414 nsew signal tristate
rlabel metal2 s 227442 163200 227498 164400 6 la_oenb[67]
port 415 nsew signal tristate
rlabel metal2 s 230846 163200 230902 164400 6 la_oenb[68]
port 416 nsew signal tristate
rlabel metal2 s 234158 163200 234214 164400 6 la_oenb[69]
port 417 nsew signal tristate
rlabel metal2 s 22190 163200 22246 164400 6 la_oenb[6]
port 418 nsew signal tristate
rlabel metal2 s 237562 163200 237618 164400 6 la_oenb[70]
port 419 nsew signal tristate
rlabel metal2 s 240874 163200 240930 164400 6 la_oenb[71]
port 420 nsew signal tristate
rlabel metal2 s 244278 163200 244334 164400 6 la_oenb[72]
port 421 nsew signal tristate
rlabel metal2 s 247682 163200 247738 164400 6 la_oenb[73]
port 422 nsew signal tristate
rlabel metal2 s 250994 163200 251050 164400 6 la_oenb[74]
port 423 nsew signal tristate
rlabel metal2 s 254398 163200 254454 164400 6 la_oenb[75]
port 424 nsew signal tristate
rlabel metal2 s 257710 163200 257766 164400 6 la_oenb[76]
port 425 nsew signal tristate
rlabel metal2 s 261114 163200 261170 164400 6 la_oenb[77]
port 426 nsew signal tristate
rlabel metal2 s 264426 163200 264482 164400 6 la_oenb[78]
port 427 nsew signal tristate
rlabel metal2 s 267830 163200 267886 164400 6 la_oenb[79]
port 428 nsew signal tristate
rlabel metal2 s 25594 163200 25650 164400 6 la_oenb[7]
port 429 nsew signal tristate
rlabel metal2 s 271234 163200 271290 164400 6 la_oenb[80]
port 430 nsew signal tristate
rlabel metal2 s 274546 163200 274602 164400 6 la_oenb[81]
port 431 nsew signal tristate
rlabel metal2 s 277950 163200 278006 164400 6 la_oenb[82]
port 432 nsew signal tristate
rlabel metal2 s 281262 163200 281318 164400 6 la_oenb[83]
port 433 nsew signal tristate
rlabel metal2 s 284666 163200 284722 164400 6 la_oenb[84]
port 434 nsew signal tristate
rlabel metal2 s 287978 163200 288034 164400 6 la_oenb[85]
port 435 nsew signal tristate
rlabel metal2 s 291382 163200 291438 164400 6 la_oenb[86]
port 436 nsew signal tristate
rlabel metal2 s 294786 163200 294842 164400 6 la_oenb[87]
port 437 nsew signal tristate
rlabel metal2 s 298098 163200 298154 164400 6 la_oenb[88]
port 438 nsew signal tristate
rlabel metal2 s 301502 163200 301558 164400 6 la_oenb[89]
port 439 nsew signal tristate
rlabel metal2 s 28906 163200 28962 164400 6 la_oenb[8]
port 440 nsew signal tristate
rlabel metal2 s 304814 163200 304870 164400 6 la_oenb[90]
port 441 nsew signal tristate
rlabel metal2 s 308218 163200 308274 164400 6 la_oenb[91]
port 442 nsew signal tristate
rlabel metal2 s 311530 163200 311586 164400 6 la_oenb[92]
port 443 nsew signal tristate
rlabel metal2 s 314934 163200 314990 164400 6 la_oenb[93]
port 444 nsew signal tristate
rlabel metal2 s 318338 163200 318394 164400 6 la_oenb[94]
port 445 nsew signal tristate
rlabel metal2 s 321650 163200 321706 164400 6 la_oenb[95]
port 446 nsew signal tristate
rlabel metal2 s 325054 163200 325110 164400 6 la_oenb[96]
port 447 nsew signal tristate
rlabel metal2 s 328366 163200 328422 164400 6 la_oenb[97]
port 448 nsew signal tristate
rlabel metal2 s 331770 163200 331826 164400 6 la_oenb[98]
port 449 nsew signal tristate
rlabel metal2 s 335082 163200 335138 164400 6 la_oenb[99]
port 450 nsew signal tristate
rlabel metal2 s 32310 163200 32366 164400 6 la_oenb[9]
port 451 nsew signal tristate
rlabel metal2 s 2870 163200 2926 164400 6 la_output[0]
port 452 nsew signal tristate
rlabel metal2 s 339314 163200 339370 164400 6 la_output[100]
port 453 nsew signal tristate
rlabel metal2 s 342718 163200 342774 164400 6 la_output[101]
port 454 nsew signal tristate
rlabel metal2 s 346030 163200 346086 164400 6 la_output[102]
port 455 nsew signal tristate
rlabel metal2 s 349434 163200 349490 164400 6 la_output[103]
port 456 nsew signal tristate
rlabel metal2 s 352746 163200 352802 164400 6 la_output[104]
port 457 nsew signal tristate
rlabel metal2 s 356150 163200 356206 164400 6 la_output[105]
port 458 nsew signal tristate
rlabel metal2 s 359554 163200 359610 164400 6 la_output[106]
port 459 nsew signal tristate
rlabel metal2 s 362866 163200 362922 164400 6 la_output[107]
port 460 nsew signal tristate
rlabel metal2 s 366270 163200 366326 164400 6 la_output[108]
port 461 nsew signal tristate
rlabel metal2 s 369582 163200 369638 164400 6 la_output[109]
port 462 nsew signal tristate
rlabel metal2 s 36542 163200 36598 164400 6 la_output[10]
port 463 nsew signal tristate
rlabel metal2 s 372986 163200 373042 164400 6 la_output[110]
port 464 nsew signal tristate
rlabel metal2 s 376298 163200 376354 164400 6 la_output[111]
port 465 nsew signal tristate
rlabel metal2 s 379702 163200 379758 164400 6 la_output[112]
port 466 nsew signal tristate
rlabel metal2 s 383106 163200 383162 164400 6 la_output[113]
port 467 nsew signal tristate
rlabel metal2 s 386418 163200 386474 164400 6 la_output[114]
port 468 nsew signal tristate
rlabel metal2 s 389822 163200 389878 164400 6 la_output[115]
port 469 nsew signal tristate
rlabel metal2 s 393134 163200 393190 164400 6 la_output[116]
port 470 nsew signal tristate
rlabel metal2 s 396538 163200 396594 164400 6 la_output[117]
port 471 nsew signal tristate
rlabel metal2 s 399850 163200 399906 164400 6 la_output[118]
port 472 nsew signal tristate
rlabel metal2 s 403254 163200 403310 164400 6 la_output[119]
port 473 nsew signal tristate
rlabel metal2 s 39854 163200 39910 164400 6 la_output[11]
port 474 nsew signal tristate
rlabel metal2 s 406658 163200 406714 164400 6 la_output[120]
port 475 nsew signal tristate
rlabel metal2 s 409970 163200 410026 164400 6 la_output[121]
port 476 nsew signal tristate
rlabel metal2 s 413374 163200 413430 164400 6 la_output[122]
port 477 nsew signal tristate
rlabel metal2 s 416686 163200 416742 164400 6 la_output[123]
port 478 nsew signal tristate
rlabel metal2 s 420090 163200 420146 164400 6 la_output[124]
port 479 nsew signal tristate
rlabel metal2 s 423402 163200 423458 164400 6 la_output[125]
port 480 nsew signal tristate
rlabel metal2 s 426806 163200 426862 164400 6 la_output[126]
port 481 nsew signal tristate
rlabel metal2 s 430210 163200 430266 164400 6 la_output[127]
port 482 nsew signal tristate
rlabel metal2 s 43258 163200 43314 164400 6 la_output[12]
port 483 nsew signal tristate
rlabel metal2 s 46570 163200 46626 164400 6 la_output[13]
port 484 nsew signal tristate
rlabel metal2 s 49974 163200 50030 164400 6 la_output[14]
port 485 nsew signal tristate
rlabel metal2 s 53378 163200 53434 164400 6 la_output[15]
port 486 nsew signal tristate
rlabel metal2 s 56690 163200 56746 164400 6 la_output[16]
port 487 nsew signal tristate
rlabel metal2 s 60094 163200 60150 164400 6 la_output[17]
port 488 nsew signal tristate
rlabel metal2 s 63406 163200 63462 164400 6 la_output[18]
port 489 nsew signal tristate
rlabel metal2 s 66810 163200 66866 164400 6 la_output[19]
port 490 nsew signal tristate
rlabel metal2 s 6274 163200 6330 164400 6 la_output[1]
port 491 nsew signal tristate
rlabel metal2 s 70122 163200 70178 164400 6 la_output[20]
port 492 nsew signal tristate
rlabel metal2 s 73526 163200 73582 164400 6 la_output[21]
port 493 nsew signal tristate
rlabel metal2 s 76930 163200 76986 164400 6 la_output[22]
port 494 nsew signal tristate
rlabel metal2 s 80242 163200 80298 164400 6 la_output[23]
port 495 nsew signal tristate
rlabel metal2 s 83646 163200 83702 164400 6 la_output[24]
port 496 nsew signal tristate
rlabel metal2 s 86958 163200 87014 164400 6 la_output[25]
port 497 nsew signal tristate
rlabel metal2 s 90362 163200 90418 164400 6 la_output[26]
port 498 nsew signal tristate
rlabel metal2 s 93674 163200 93730 164400 6 la_output[27]
port 499 nsew signal tristate
rlabel metal2 s 97078 163200 97134 164400 6 la_output[28]
port 500 nsew signal tristate
rlabel metal2 s 100482 163200 100538 164400 6 la_output[29]
port 501 nsew signal tristate
rlabel metal2 s 9586 163200 9642 164400 6 la_output[2]
port 502 nsew signal tristate
rlabel metal2 s 103794 163200 103850 164400 6 la_output[30]
port 503 nsew signal tristate
rlabel metal2 s 107198 163200 107254 164400 6 la_output[31]
port 504 nsew signal tristate
rlabel metal2 s 110510 163200 110566 164400 6 la_output[32]
port 505 nsew signal tristate
rlabel metal2 s 113914 163200 113970 164400 6 la_output[33]
port 506 nsew signal tristate
rlabel metal2 s 117226 163200 117282 164400 6 la_output[34]
port 507 nsew signal tristate
rlabel metal2 s 120630 163200 120686 164400 6 la_output[35]
port 508 nsew signal tristate
rlabel metal2 s 124034 163200 124090 164400 6 la_output[36]
port 509 nsew signal tristate
rlabel metal2 s 127346 163200 127402 164400 6 la_output[37]
port 510 nsew signal tristate
rlabel metal2 s 130750 163200 130806 164400 6 la_output[38]
port 511 nsew signal tristate
rlabel metal2 s 134062 163200 134118 164400 6 la_output[39]
port 512 nsew signal tristate
rlabel metal2 s 12990 163200 13046 164400 6 la_output[3]
port 513 nsew signal tristate
rlabel metal2 s 137466 163200 137522 164400 6 la_output[40]
port 514 nsew signal tristate
rlabel metal2 s 140778 163200 140834 164400 6 la_output[41]
port 515 nsew signal tristate
rlabel metal2 s 144182 163200 144238 164400 6 la_output[42]
port 516 nsew signal tristate
rlabel metal2 s 147586 163200 147642 164400 6 la_output[43]
port 517 nsew signal tristate
rlabel metal2 s 150898 163200 150954 164400 6 la_output[44]
port 518 nsew signal tristate
rlabel metal2 s 154302 163200 154358 164400 6 la_output[45]
port 519 nsew signal tristate
rlabel metal2 s 157614 163200 157670 164400 6 la_output[46]
port 520 nsew signal tristate
rlabel metal2 s 161018 163200 161074 164400 6 la_output[47]
port 521 nsew signal tristate
rlabel metal2 s 164330 163200 164386 164400 6 la_output[48]
port 522 nsew signal tristate
rlabel metal2 s 167734 163200 167790 164400 6 la_output[49]
port 523 nsew signal tristate
rlabel metal2 s 16302 163200 16358 164400 6 la_output[4]
port 524 nsew signal tristate
rlabel metal2 s 171138 163200 171194 164400 6 la_output[50]
port 525 nsew signal tristate
rlabel metal2 s 174450 163200 174506 164400 6 la_output[51]
port 526 nsew signal tristate
rlabel metal2 s 177854 163200 177910 164400 6 la_output[52]
port 527 nsew signal tristate
rlabel metal2 s 181166 163200 181222 164400 6 la_output[53]
port 528 nsew signal tristate
rlabel metal2 s 184570 163200 184626 164400 6 la_output[54]
port 529 nsew signal tristate
rlabel metal2 s 187882 163200 187938 164400 6 la_output[55]
port 530 nsew signal tristate
rlabel metal2 s 191286 163200 191342 164400 6 la_output[56]
port 531 nsew signal tristate
rlabel metal2 s 194690 163200 194746 164400 6 la_output[57]
port 532 nsew signal tristate
rlabel metal2 s 198002 163200 198058 164400 6 la_output[58]
port 533 nsew signal tristate
rlabel metal2 s 201406 163200 201462 164400 6 la_output[59]
port 534 nsew signal tristate
rlabel metal2 s 19706 163200 19762 164400 6 la_output[5]
port 535 nsew signal tristate
rlabel metal2 s 204718 163200 204774 164400 6 la_output[60]
port 536 nsew signal tristate
rlabel metal2 s 208122 163200 208178 164400 6 la_output[61]
port 537 nsew signal tristate
rlabel metal2 s 211434 163200 211490 164400 6 la_output[62]
port 538 nsew signal tristate
rlabel metal2 s 214838 163200 214894 164400 6 la_output[63]
port 539 nsew signal tristate
rlabel metal2 s 218242 163200 218298 164400 6 la_output[64]
port 540 nsew signal tristate
rlabel metal2 s 221554 163200 221610 164400 6 la_output[65]
port 541 nsew signal tristate
rlabel metal2 s 224958 163200 225014 164400 6 la_output[66]
port 542 nsew signal tristate
rlabel metal2 s 228270 163200 228326 164400 6 la_output[67]
port 543 nsew signal tristate
rlabel metal2 s 231674 163200 231730 164400 6 la_output[68]
port 544 nsew signal tristate
rlabel metal2 s 234986 163200 235042 164400 6 la_output[69]
port 545 nsew signal tristate
rlabel metal2 s 23018 163200 23074 164400 6 la_output[6]
port 546 nsew signal tristate
rlabel metal2 s 238390 163200 238446 164400 6 la_output[70]
port 547 nsew signal tristate
rlabel metal2 s 241794 163200 241850 164400 6 la_output[71]
port 548 nsew signal tristate
rlabel metal2 s 245106 163200 245162 164400 6 la_output[72]
port 549 nsew signal tristate
rlabel metal2 s 248510 163200 248566 164400 6 la_output[73]
port 550 nsew signal tristate
rlabel metal2 s 251822 163200 251878 164400 6 la_output[74]
port 551 nsew signal tristate
rlabel metal2 s 255226 163200 255282 164400 6 la_output[75]
port 552 nsew signal tristate
rlabel metal2 s 258538 163200 258594 164400 6 la_output[76]
port 553 nsew signal tristate
rlabel metal2 s 261942 163200 261998 164400 6 la_output[77]
port 554 nsew signal tristate
rlabel metal2 s 265346 163200 265402 164400 6 la_output[78]
port 555 nsew signal tristate
rlabel metal2 s 268658 163200 268714 164400 6 la_output[79]
port 556 nsew signal tristate
rlabel metal2 s 26422 163200 26478 164400 6 la_output[7]
port 557 nsew signal tristate
rlabel metal2 s 272062 163200 272118 164400 6 la_output[80]
port 558 nsew signal tristate
rlabel metal2 s 275374 163200 275430 164400 6 la_output[81]
port 559 nsew signal tristate
rlabel metal2 s 278778 163200 278834 164400 6 la_output[82]
port 560 nsew signal tristate
rlabel metal2 s 282090 163200 282146 164400 6 la_output[83]
port 561 nsew signal tristate
rlabel metal2 s 285494 163200 285550 164400 6 la_output[84]
port 562 nsew signal tristate
rlabel metal2 s 288898 163200 288954 164400 6 la_output[85]
port 563 nsew signal tristate
rlabel metal2 s 292210 163200 292266 164400 6 la_output[86]
port 564 nsew signal tristate
rlabel metal2 s 295614 163200 295670 164400 6 la_output[87]
port 565 nsew signal tristate
rlabel metal2 s 298926 163200 298982 164400 6 la_output[88]
port 566 nsew signal tristate
rlabel metal2 s 302330 163200 302386 164400 6 la_output[89]
port 567 nsew signal tristate
rlabel metal2 s 29826 163200 29882 164400 6 la_output[8]
port 568 nsew signal tristate
rlabel metal2 s 305642 163200 305698 164400 6 la_output[90]
port 569 nsew signal tristate
rlabel metal2 s 309046 163200 309102 164400 6 la_output[91]
port 570 nsew signal tristate
rlabel metal2 s 312450 163200 312506 164400 6 la_output[92]
port 571 nsew signal tristate
rlabel metal2 s 315762 163200 315818 164400 6 la_output[93]
port 572 nsew signal tristate
rlabel metal2 s 319166 163200 319222 164400 6 la_output[94]
port 573 nsew signal tristate
rlabel metal2 s 322478 163200 322534 164400 6 la_output[95]
port 574 nsew signal tristate
rlabel metal2 s 325882 163200 325938 164400 6 la_output[96]
port 575 nsew signal tristate
rlabel metal2 s 329194 163200 329250 164400 6 la_output[97]
port 576 nsew signal tristate
rlabel metal2 s 332598 163200 332654 164400 6 la_output[98]
port 577 nsew signal tristate
rlabel metal2 s 336002 163200 336058 164400 6 la_output[99]
port 578 nsew signal tristate
rlabel metal2 s 33138 163200 33194 164400 6 la_output[9]
port 579 nsew signal tristate
rlabel metal2 s 431038 163200 431094 164400 6 mprj_ack_i
port 580 nsew signal input
rlabel metal2 s 435178 163200 435234 164400 6 mprj_adr_o[0]
port 581 nsew signal tristate
rlabel metal2 s 463790 163200 463846 164400 6 mprj_adr_o[10]
port 582 nsew signal tristate
rlabel metal2 s 466366 163200 466422 164400 6 mprj_adr_o[11]
port 583 nsew signal tristate
rlabel metal2 s 468850 163200 468906 164400 6 mprj_adr_o[12]
port 584 nsew signal tristate
rlabel metal2 s 471426 163200 471482 164400 6 mprj_adr_o[13]
port 585 nsew signal tristate
rlabel metal2 s 473910 163200 473966 164400 6 mprj_adr_o[14]
port 586 nsew signal tristate
rlabel metal2 s 476394 163200 476450 164400 6 mprj_adr_o[15]
port 587 nsew signal tristate
rlabel metal2 s 478970 163200 479026 164400 6 mprj_adr_o[16]
port 588 nsew signal tristate
rlabel metal2 s 481454 163200 481510 164400 6 mprj_adr_o[17]
port 589 nsew signal tristate
rlabel metal2 s 484030 163200 484086 164400 6 mprj_adr_o[18]
port 590 nsew signal tristate
rlabel metal2 s 486514 163200 486570 164400 6 mprj_adr_o[19]
port 591 nsew signal tristate
rlabel metal2 s 438582 163200 438638 164400 6 mprj_adr_o[1]
port 592 nsew signal tristate
rlabel metal2 s 489090 163200 489146 164400 6 mprj_adr_o[20]
port 593 nsew signal tristate
rlabel metal2 s 491574 163200 491630 164400 6 mprj_adr_o[21]
port 594 nsew signal tristate
rlabel metal2 s 494058 163200 494114 164400 6 mprj_adr_o[22]
port 595 nsew signal tristate
rlabel metal2 s 496634 163200 496690 164400 6 mprj_adr_o[23]
port 596 nsew signal tristate
rlabel metal2 s 499118 163200 499174 164400 6 mprj_adr_o[24]
port 597 nsew signal tristate
rlabel metal2 s 501694 163200 501750 164400 6 mprj_adr_o[25]
port 598 nsew signal tristate
rlabel metal2 s 504178 163200 504234 164400 6 mprj_adr_o[26]
port 599 nsew signal tristate
rlabel metal2 s 506754 163200 506810 164400 6 mprj_adr_o[27]
port 600 nsew signal tristate
rlabel metal2 s 509238 163200 509294 164400 6 mprj_adr_o[28]
port 601 nsew signal tristate
rlabel metal2 s 511722 163200 511778 164400 6 mprj_adr_o[29]
port 602 nsew signal tristate
rlabel metal2 s 441986 163200 442042 164400 6 mprj_adr_o[2]
port 603 nsew signal tristate
rlabel metal2 s 514298 163200 514354 164400 6 mprj_adr_o[30]
port 604 nsew signal tristate
rlabel metal2 s 516782 163200 516838 164400 6 mprj_adr_o[31]
port 605 nsew signal tristate
rlabel metal2 s 445298 163200 445354 164400 6 mprj_adr_o[3]
port 606 nsew signal tristate
rlabel metal2 s 448702 163200 448758 164400 6 mprj_adr_o[4]
port 607 nsew signal tristate
rlabel metal2 s 451186 163200 451242 164400 6 mprj_adr_o[5]
port 608 nsew signal tristate
rlabel metal2 s 453762 163200 453818 164400 6 mprj_adr_o[6]
port 609 nsew signal tristate
rlabel metal2 s 456246 163200 456302 164400 6 mprj_adr_o[7]
port 610 nsew signal tristate
rlabel metal2 s 458730 163200 458786 164400 6 mprj_adr_o[8]
port 611 nsew signal tristate
rlabel metal2 s 461306 163200 461362 164400 6 mprj_adr_o[9]
port 612 nsew signal tristate
rlabel metal2 s 431866 163200 431922 164400 6 mprj_cyc_o
port 613 nsew signal tristate
rlabel metal2 s 436098 163200 436154 164400 6 mprj_dat_i[0]
port 614 nsew signal input
rlabel metal2 s 464618 163200 464674 164400 6 mprj_dat_i[10]
port 615 nsew signal input
rlabel metal2 s 467194 163200 467250 164400 6 mprj_dat_i[11]
port 616 nsew signal input
rlabel metal2 s 469678 163200 469734 164400 6 mprj_dat_i[12]
port 617 nsew signal input
rlabel metal2 s 472254 163200 472310 164400 6 mprj_dat_i[13]
port 618 nsew signal input
rlabel metal2 s 474738 163200 474794 164400 6 mprj_dat_i[14]
port 619 nsew signal input
rlabel metal2 s 477314 163200 477370 164400 6 mprj_dat_i[15]
port 620 nsew signal input
rlabel metal2 s 479798 163200 479854 164400 6 mprj_dat_i[16]
port 621 nsew signal input
rlabel metal2 s 482282 163200 482338 164400 6 mprj_dat_i[17]
port 622 nsew signal input
rlabel metal2 s 484858 163200 484914 164400 6 mprj_dat_i[18]
port 623 nsew signal input
rlabel metal2 s 487342 163200 487398 164400 6 mprj_dat_i[19]
port 624 nsew signal input
rlabel metal2 s 439410 163200 439466 164400 6 mprj_dat_i[1]
port 625 nsew signal input
rlabel metal2 s 489918 163200 489974 164400 6 mprj_dat_i[20]
port 626 nsew signal input
rlabel metal2 s 492402 163200 492458 164400 6 mprj_dat_i[21]
port 627 nsew signal input
rlabel metal2 s 494978 163200 495034 164400 6 mprj_dat_i[22]
port 628 nsew signal input
rlabel metal2 s 497462 163200 497518 164400 6 mprj_dat_i[23]
port 629 nsew signal input
rlabel metal2 s 499946 163200 500002 164400 6 mprj_dat_i[24]
port 630 nsew signal input
rlabel metal2 s 502522 163200 502578 164400 6 mprj_dat_i[25]
port 631 nsew signal input
rlabel metal2 s 505006 163200 505062 164400 6 mprj_dat_i[26]
port 632 nsew signal input
rlabel metal2 s 507582 163200 507638 164400 6 mprj_dat_i[27]
port 633 nsew signal input
rlabel metal2 s 510066 163200 510122 164400 6 mprj_dat_i[28]
port 634 nsew signal input
rlabel metal2 s 512642 163200 512698 164400 6 mprj_dat_i[29]
port 635 nsew signal input
rlabel metal2 s 442814 163200 442870 164400 6 mprj_dat_i[2]
port 636 nsew signal input
rlabel metal2 s 515126 163200 515182 164400 6 mprj_dat_i[30]
port 637 nsew signal input
rlabel metal2 s 517610 163200 517666 164400 6 mprj_dat_i[31]
port 638 nsew signal input
rlabel metal2 s 446126 163200 446182 164400 6 mprj_dat_i[3]
port 639 nsew signal input
rlabel metal2 s 449530 163200 449586 164400 6 mprj_dat_i[4]
port 640 nsew signal input
rlabel metal2 s 452014 163200 452070 164400 6 mprj_dat_i[5]
port 641 nsew signal input
rlabel metal2 s 454590 163200 454646 164400 6 mprj_dat_i[6]
port 642 nsew signal input
rlabel metal2 s 457074 163200 457130 164400 6 mprj_dat_i[7]
port 643 nsew signal input
rlabel metal2 s 459650 163200 459706 164400 6 mprj_dat_i[8]
port 644 nsew signal input
rlabel metal2 s 462134 163200 462190 164400 6 mprj_dat_i[9]
port 645 nsew signal input
rlabel metal2 s 436926 163200 436982 164400 6 mprj_dat_o[0]
port 646 nsew signal tristate
rlabel metal2 s 465538 163200 465594 164400 6 mprj_dat_o[10]
port 647 nsew signal tristate
rlabel metal2 s 468022 163200 468078 164400 6 mprj_dat_o[11]
port 648 nsew signal tristate
rlabel metal2 s 470506 163200 470562 164400 6 mprj_dat_o[12]
port 649 nsew signal tristate
rlabel metal2 s 473082 163200 473138 164400 6 mprj_dat_o[13]
port 650 nsew signal tristate
rlabel metal2 s 475566 163200 475622 164400 6 mprj_dat_o[14]
port 651 nsew signal tristate
rlabel metal2 s 478142 163200 478198 164400 6 mprj_dat_o[15]
port 652 nsew signal tristate
rlabel metal2 s 480626 163200 480682 164400 6 mprj_dat_o[16]
port 653 nsew signal tristate
rlabel metal2 s 483202 163200 483258 164400 6 mprj_dat_o[17]
port 654 nsew signal tristate
rlabel metal2 s 485686 163200 485742 164400 6 mprj_dat_o[18]
port 655 nsew signal tristate
rlabel metal2 s 488170 163200 488226 164400 6 mprj_dat_o[19]
port 656 nsew signal tristate
rlabel metal2 s 440238 163200 440294 164400 6 mprj_dat_o[1]
port 657 nsew signal tristate
rlabel metal2 s 490746 163200 490802 164400 6 mprj_dat_o[20]
port 658 nsew signal tristate
rlabel metal2 s 493230 163200 493286 164400 6 mprj_dat_o[21]
port 659 nsew signal tristate
rlabel metal2 s 495806 163200 495862 164400 6 mprj_dat_o[22]
port 660 nsew signal tristate
rlabel metal2 s 498290 163200 498346 164400 6 mprj_dat_o[23]
port 661 nsew signal tristate
rlabel metal2 s 500866 163200 500922 164400 6 mprj_dat_o[24]
port 662 nsew signal tristate
rlabel metal2 s 503350 163200 503406 164400 6 mprj_dat_o[25]
port 663 nsew signal tristate
rlabel metal2 s 505834 163200 505890 164400 6 mprj_dat_o[26]
port 664 nsew signal tristate
rlabel metal2 s 508410 163200 508466 164400 6 mprj_dat_o[27]
port 665 nsew signal tristate
rlabel metal2 s 510894 163200 510950 164400 6 mprj_dat_o[28]
port 666 nsew signal tristate
rlabel metal2 s 513470 163200 513526 164400 6 mprj_dat_o[29]
port 667 nsew signal tristate
rlabel metal2 s 443642 163200 443698 164400 6 mprj_dat_o[2]
port 668 nsew signal tristate
rlabel metal2 s 515954 163200 516010 164400 6 mprj_dat_o[30]
port 669 nsew signal tristate
rlabel metal2 s 518530 163200 518586 164400 6 mprj_dat_o[31]
port 670 nsew signal tristate
rlabel metal2 s 446954 163200 447010 164400 6 mprj_dat_o[3]
port 671 nsew signal tristate
rlabel metal2 s 450358 163200 450414 164400 6 mprj_dat_o[4]
port 672 nsew signal tristate
rlabel metal2 s 452842 163200 452898 164400 6 mprj_dat_o[5]
port 673 nsew signal tristate
rlabel metal2 s 455418 163200 455474 164400 6 mprj_dat_o[6]
port 674 nsew signal tristate
rlabel metal2 s 457902 163200 457958 164400 6 mprj_dat_o[7]
port 675 nsew signal tristate
rlabel metal2 s 460478 163200 460534 164400 6 mprj_dat_o[8]
port 676 nsew signal tristate
rlabel metal2 s 462962 163200 463018 164400 6 mprj_dat_o[9]
port 677 nsew signal tristate
rlabel metal2 s 437754 163200 437810 164400 6 mprj_sel_o[0]
port 678 nsew signal tristate
rlabel metal2 s 441066 163200 441122 164400 6 mprj_sel_o[1]
port 679 nsew signal tristate
rlabel metal2 s 444470 163200 444526 164400 6 mprj_sel_o[2]
port 680 nsew signal tristate
rlabel metal2 s 447874 163200 447930 164400 6 mprj_sel_o[3]
port 681 nsew signal tristate
rlabel metal2 s 432694 163200 432750 164400 6 mprj_stb_o
port 682 nsew signal tristate
rlabel metal2 s 433522 163200 433578 164400 6 mprj_wb_iena
port 683 nsew signal tristate
rlabel metal2 s 434350 163200 434406 164400 6 mprj_we_o
port 684 nsew signal tristate
rlabel metal3 s 523200 90176 524400 90296 6 qspi_enabled
port 685 nsew signal tristate
rlabel metal3 s 523200 84192 524400 84312 6 ser_rx
port 686 nsew signal input
rlabel metal3 s 523200 85688 524400 85808 6 ser_tx
port 687 nsew signal tristate
rlabel metal3 s 523200 81064 524400 81184 6 spi_csb
port 688 nsew signal tristate
rlabel metal3 s 523200 87184 524400 87304 6 spi_enabled
port 689 nsew signal tristate
rlabel metal3 s 523200 79568 524400 79688 6 spi_sck
port 690 nsew signal tristate
rlabel metal3 s 523200 82696 524400 82816 6 spi_sdi
port 691 nsew signal input
rlabel metal3 s 523200 78072 524400 78192 6 spi_sdo
port 692 nsew signal tristate
rlabel metal3 s 523200 76576 524400 76696 6 spi_sdoenb
port 693 nsew signal tristate
rlabel metal3 s 523200 2184 524400 2304 6 sram_ro_addr[0]
port 694 nsew signal input
rlabel metal3 s 523200 3680 524400 3800 6 sram_ro_addr[1]
port 695 nsew signal input
rlabel metal3 s 523200 5176 524400 5296 6 sram_ro_addr[2]
port 696 nsew signal input
rlabel metal3 s 523200 6672 524400 6792 6 sram_ro_addr[3]
port 697 nsew signal input
rlabel metal3 s 523200 8168 524400 8288 6 sram_ro_addr[4]
port 698 nsew signal input
rlabel metal3 s 523200 9800 524400 9920 6 sram_ro_addr[5]
port 699 nsew signal input
rlabel metal3 s 523200 11296 524400 11416 6 sram_ro_addr[6]
port 700 nsew signal input
rlabel metal3 s 523200 12792 524400 12912 6 sram_ro_addr[7]
port 701 nsew signal input
rlabel metal3 s 523200 14288 524400 14408 6 sram_ro_clk
port 702 nsew signal input
rlabel metal3 s 523200 688 524400 808 6 sram_ro_csb
port 703 nsew signal input
rlabel metal3 s 523200 15784 524400 15904 6 sram_ro_data[0]
port 704 nsew signal tristate
rlabel metal3 s 523200 31016 524400 31136 6 sram_ro_data[10]
port 705 nsew signal tristate
rlabel metal3 s 523200 32512 524400 32632 6 sram_ro_data[11]
port 706 nsew signal tristate
rlabel metal3 s 523200 34008 524400 34128 6 sram_ro_data[12]
port 707 nsew signal tristate
rlabel metal3 s 523200 35504 524400 35624 6 sram_ro_data[13]
port 708 nsew signal tristate
rlabel metal3 s 523200 37136 524400 37256 6 sram_ro_data[14]
port 709 nsew signal tristate
rlabel metal3 s 523200 38632 524400 38752 6 sram_ro_data[15]
port 710 nsew signal tristate
rlabel metal3 s 523200 40128 524400 40248 6 sram_ro_data[16]
port 711 nsew signal tristate
rlabel metal3 s 523200 41624 524400 41744 6 sram_ro_data[17]
port 712 nsew signal tristate
rlabel metal3 s 523200 43120 524400 43240 6 sram_ro_data[18]
port 713 nsew signal tristate
rlabel metal3 s 523200 44616 524400 44736 6 sram_ro_data[19]
port 714 nsew signal tristate
rlabel metal3 s 523200 17280 524400 17400 6 sram_ro_data[1]
port 715 nsew signal tristate
rlabel metal3 s 523200 46248 524400 46368 6 sram_ro_data[20]
port 716 nsew signal tristate
rlabel metal3 s 523200 47744 524400 47864 6 sram_ro_data[21]
port 717 nsew signal tristate
rlabel metal3 s 523200 49240 524400 49360 6 sram_ro_data[22]
port 718 nsew signal tristate
rlabel metal3 s 523200 50736 524400 50856 6 sram_ro_data[23]
port 719 nsew signal tristate
rlabel metal3 s 523200 52232 524400 52352 6 sram_ro_data[24]
port 720 nsew signal tristate
rlabel metal3 s 523200 53728 524400 53848 6 sram_ro_data[25]
port 721 nsew signal tristate
rlabel metal3 s 523200 55360 524400 55480 6 sram_ro_data[26]
port 722 nsew signal tristate
rlabel metal3 s 523200 56856 524400 56976 6 sram_ro_data[27]
port 723 nsew signal tristate
rlabel metal3 s 523200 58352 524400 58472 6 sram_ro_data[28]
port 724 nsew signal tristate
rlabel metal3 s 523200 59848 524400 59968 6 sram_ro_data[29]
port 725 nsew signal tristate
rlabel metal3 s 523200 18912 524400 19032 6 sram_ro_data[2]
port 726 nsew signal tristate
rlabel metal3 s 523200 61344 524400 61464 6 sram_ro_data[30]
port 727 nsew signal tristate
rlabel metal3 s 523200 62840 524400 62960 6 sram_ro_data[31]
port 728 nsew signal tristate
rlabel metal3 s 523200 20408 524400 20528 6 sram_ro_data[3]
port 729 nsew signal tristate
rlabel metal3 s 523200 21904 524400 22024 6 sram_ro_data[4]
port 730 nsew signal tristate
rlabel metal3 s 523200 23400 524400 23520 6 sram_ro_data[5]
port 731 nsew signal tristate
rlabel metal3 s 523200 24896 524400 25016 6 sram_ro_data[6]
port 732 nsew signal tristate
rlabel metal3 s 523200 26392 524400 26512 6 sram_ro_data[7]
port 733 nsew signal tristate
rlabel metal3 s 523200 28024 524400 28144 6 sram_ro_data[8]
port 734 nsew signal tristate
rlabel metal3 s 523200 29520 524400 29640 6 sram_ro_data[9]
port 735 nsew signal tristate
rlabel metal3 s 523200 70456 524400 70576 6 trap
port 736 nsew signal tristate
rlabel metal3 s 523200 88680 524400 88800 6 uart_enabled
port 737 nsew signal tristate
rlabel metal2 s 519358 163200 519414 164400 6 user_irq_ena[0]
port 738 nsew signal tristate
rlabel metal2 s 520186 163200 520242 164400 6 user_irq_ena[1]
port 739 nsew signal tristate
rlabel metal2 s 521014 163200 521070 164400 6 user_irq_ena[2]
port 740 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 524000 164000
<< end >>
