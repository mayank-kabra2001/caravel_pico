magic
tech sky130A
magscale 1 2
timestamp 1635525820
<< obsli1 >>
rect 1104 2159 169067 107729
<< obsm1 >>
rect 1104 2048 169079 107760
<< metal2 >>
rect 6550 109200 6606 110000
rect 19614 109200 19670 110000
rect 32678 109200 32734 110000
rect 45742 109200 45798 110000
rect 58806 109200 58862 110000
rect 71870 109200 71926 110000
rect 84934 109200 84990 110000
rect 98090 109200 98146 110000
rect 111154 109200 111210 110000
rect 124218 109200 124274 110000
rect 137282 109200 137338 110000
rect 150346 109200 150402 110000
rect 163410 109200 163466 110000
rect 85026 0 85082 800
<< obsm2 >>
rect 1400 109144 6494 109290
rect 6662 109144 19558 109290
rect 19726 109144 32622 109290
rect 32790 109144 45686 109290
rect 45854 109144 58750 109290
rect 58918 109144 71814 109290
rect 71982 109144 84878 109290
rect 85046 109144 98034 109290
rect 98202 109144 111098 109290
rect 111266 109144 124162 109290
rect 124330 109144 137226 109290
rect 137394 109144 150290 109290
rect 150458 109144 163354 109290
rect 163522 109144 168986 109290
rect 1400 856 168986 109144
rect 1400 734 84970 856
rect 85138 734 168986 856
<< metal3 >>
rect 0 108128 800 108248
rect 169200 108128 170000 108248
rect 0 104728 800 104848
rect 169200 104728 170000 104848
rect 0 101328 800 101448
rect 169200 101328 170000 101448
rect 0 97792 800 97912
rect 169200 97792 170000 97912
rect 0 94392 800 94512
rect 169200 94392 170000 94512
rect 0 90992 800 91112
rect 169200 90992 170000 91112
rect 0 87592 800 87712
rect 169200 87592 170000 87712
rect 0 84056 800 84176
rect 169200 84056 170000 84176
rect 0 80656 800 80776
rect 169200 80656 170000 80776
rect 0 77256 800 77376
rect 169200 77256 170000 77376
rect 0 73720 800 73840
rect 169200 73720 170000 73840
rect 0 70320 800 70440
rect 169200 70320 170000 70440
rect 0 66920 800 67040
rect 169200 66920 170000 67040
rect 0 63520 800 63640
rect 169200 63520 170000 63640
rect 0 59984 800 60104
rect 169200 59984 170000 60104
rect 0 56584 800 56704
rect 169200 56584 170000 56704
rect 0 53184 800 53304
rect 169200 53184 170000 53304
rect 0 49648 800 49768
rect 169200 49648 170000 49768
rect 0 46248 800 46368
rect 169200 46248 170000 46368
rect 0 42848 800 42968
rect 169200 42848 170000 42968
rect 0 39448 800 39568
rect 169200 39448 170000 39568
rect 0 35912 800 36032
rect 169200 35912 170000 36032
rect 0 32512 800 32632
rect 169200 32512 170000 32632
rect 0 29112 800 29232
rect 169200 29112 170000 29232
rect 0 25576 800 25696
rect 169200 25576 170000 25696
rect 0 22176 800 22296
rect 169200 22176 170000 22296
rect 0 18776 800 18896
rect 169200 18776 170000 18896
rect 0 15376 800 15496
rect 169200 15376 170000 15496
rect 0 11840 800 11960
rect 169200 11840 170000 11960
rect 0 8440 800 8560
rect 169200 8440 170000 8560
rect 0 5040 800 5160
rect 169200 5040 170000 5160
rect 0 1640 800 1760
rect 169200 1640 170000 1760
<< obsm3 >>
rect 880 108048 169120 108221
rect 800 104928 169200 108048
rect 880 104648 169120 104928
rect 800 101528 169200 104648
rect 880 101248 169120 101528
rect 800 97992 169200 101248
rect 880 97712 169120 97992
rect 800 94592 169200 97712
rect 880 94312 169120 94592
rect 800 91192 169200 94312
rect 880 90912 169120 91192
rect 800 87792 169200 90912
rect 880 87512 169120 87792
rect 800 84256 169200 87512
rect 880 83976 169120 84256
rect 800 80856 169200 83976
rect 880 80576 169120 80856
rect 800 77456 169200 80576
rect 880 77176 169120 77456
rect 800 73920 169200 77176
rect 880 73640 169120 73920
rect 800 70520 169200 73640
rect 880 70240 169120 70520
rect 800 67120 169200 70240
rect 880 66840 169120 67120
rect 800 63720 169200 66840
rect 880 63440 169120 63720
rect 800 60184 169200 63440
rect 880 59904 169120 60184
rect 800 56784 169200 59904
rect 880 56504 169120 56784
rect 800 53384 169200 56504
rect 880 53104 169120 53384
rect 800 49848 169200 53104
rect 880 49568 169120 49848
rect 800 46448 169200 49568
rect 880 46168 169120 46448
rect 800 43048 169200 46168
rect 880 42768 169120 43048
rect 800 39648 169200 42768
rect 880 39368 169120 39648
rect 800 36112 169200 39368
rect 880 35832 169120 36112
rect 800 32712 169200 35832
rect 880 32432 169120 32712
rect 800 29312 169200 32432
rect 880 29032 169120 29312
rect 800 25776 169200 29032
rect 880 25496 169120 25776
rect 800 22376 169200 25496
rect 880 22096 169120 22376
rect 800 18976 169200 22096
rect 880 18696 169120 18976
rect 800 15576 169200 18696
rect 880 15296 169120 15576
rect 800 12040 169200 15296
rect 880 11760 169120 12040
rect 800 8640 169200 11760
rect 880 8360 169120 8640
rect 800 5240 169200 8360
rect 880 4960 169120 5240
rect 800 1840 169200 4960
rect 880 1667 169120 1840
<< metal4 >>
rect 4208 2128 4528 107760
rect 19568 2128 19888 107760
rect 34928 2128 35248 107760
rect 50288 2128 50608 107760
rect 65648 2128 65968 107760
rect 81008 2128 81328 107760
rect 96368 2128 96688 107760
rect 111728 2128 112048 107760
rect 127088 2128 127408 107760
rect 142448 2128 142768 107760
rect 157808 2128 158128 107760
<< obsm4 >>
rect 5027 5203 19488 105637
rect 19968 5203 34848 105637
rect 35328 5203 50208 105637
rect 50688 5203 65568 105637
rect 66048 5203 80928 105637
rect 81408 5203 96288 105637
rect 96768 5203 111648 105637
rect 112128 5203 127008 105637
rect 127488 5203 142368 105637
rect 142848 5203 153949 105637
<< metal5 >>
rect 1104 97206 168820 97526
rect 1104 81888 168820 82208
rect 1104 66570 168820 66890
rect 1104 51252 168820 51572
rect 1104 35934 168820 36254
rect 1104 20616 168820 20936
rect 1104 5298 168820 5618
<< labels >>
rlabel metal2 s 6550 109200 6606 110000 6 A[0]
port 1 nsew signal input
rlabel metal2 s 19614 109200 19670 110000 6 A[1]
port 2 nsew signal input
rlabel metal2 s 32678 109200 32734 110000 6 A[2]
port 3 nsew signal input
rlabel metal2 s 45742 109200 45798 110000 6 A[3]
port 4 nsew signal input
rlabel metal2 s 58806 109200 58862 110000 6 A[4]
port 5 nsew signal input
rlabel metal2 s 71870 109200 71926 110000 6 A[5]
port 6 nsew signal input
rlabel metal2 s 84934 109200 84990 110000 6 A[6]
port 7 nsew signal input
rlabel metal2 s 98090 109200 98146 110000 6 A[7]
port 8 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 CLK
port 9 nsew signal input
rlabel metal3 s 169200 1640 170000 1760 6 Di[0]
port 10 nsew signal input
rlabel metal3 s 169200 35912 170000 36032 6 Di[10]
port 11 nsew signal input
rlabel metal3 s 169200 39448 170000 39568 6 Di[11]
port 12 nsew signal input
rlabel metal3 s 169200 42848 170000 42968 6 Di[12]
port 13 nsew signal input
rlabel metal3 s 169200 46248 170000 46368 6 Di[13]
port 14 nsew signal input
rlabel metal3 s 169200 49648 170000 49768 6 Di[14]
port 15 nsew signal input
rlabel metal3 s 169200 53184 170000 53304 6 Di[15]
port 16 nsew signal input
rlabel metal3 s 169200 56584 170000 56704 6 Di[16]
port 17 nsew signal input
rlabel metal3 s 169200 59984 170000 60104 6 Di[17]
port 18 nsew signal input
rlabel metal3 s 169200 63520 170000 63640 6 Di[18]
port 19 nsew signal input
rlabel metal3 s 169200 66920 170000 67040 6 Di[19]
port 20 nsew signal input
rlabel metal3 s 169200 5040 170000 5160 6 Di[1]
port 21 nsew signal input
rlabel metal3 s 169200 70320 170000 70440 6 Di[20]
port 22 nsew signal input
rlabel metal3 s 169200 73720 170000 73840 6 Di[21]
port 23 nsew signal input
rlabel metal3 s 169200 77256 170000 77376 6 Di[22]
port 24 nsew signal input
rlabel metal3 s 169200 80656 170000 80776 6 Di[23]
port 25 nsew signal input
rlabel metal3 s 169200 84056 170000 84176 6 Di[24]
port 26 nsew signal input
rlabel metal3 s 169200 87592 170000 87712 6 Di[25]
port 27 nsew signal input
rlabel metal3 s 169200 90992 170000 91112 6 Di[26]
port 28 nsew signal input
rlabel metal3 s 169200 94392 170000 94512 6 Di[27]
port 29 nsew signal input
rlabel metal3 s 169200 97792 170000 97912 6 Di[28]
port 30 nsew signal input
rlabel metal3 s 169200 101328 170000 101448 6 Di[29]
port 31 nsew signal input
rlabel metal3 s 169200 8440 170000 8560 6 Di[2]
port 32 nsew signal input
rlabel metal3 s 169200 104728 170000 104848 6 Di[30]
port 33 nsew signal input
rlabel metal3 s 169200 108128 170000 108248 6 Di[31]
port 34 nsew signal input
rlabel metal3 s 169200 11840 170000 11960 6 Di[3]
port 35 nsew signal input
rlabel metal3 s 169200 15376 170000 15496 6 Di[4]
port 36 nsew signal input
rlabel metal3 s 169200 18776 170000 18896 6 Di[5]
port 37 nsew signal input
rlabel metal3 s 169200 22176 170000 22296 6 Di[6]
port 38 nsew signal input
rlabel metal3 s 169200 25576 170000 25696 6 Di[7]
port 39 nsew signal input
rlabel metal3 s 169200 29112 170000 29232 6 Di[8]
port 40 nsew signal input
rlabel metal3 s 169200 32512 170000 32632 6 Di[9]
port 41 nsew signal input
rlabel metal3 s 0 1640 800 1760 6 Do[0]
port 42 nsew signal output
rlabel metal3 s 0 35912 800 36032 6 Do[10]
port 43 nsew signal output
rlabel metal3 s 0 39448 800 39568 6 Do[11]
port 44 nsew signal output
rlabel metal3 s 0 42848 800 42968 6 Do[12]
port 45 nsew signal output
rlabel metal3 s 0 46248 800 46368 6 Do[13]
port 46 nsew signal output
rlabel metal3 s 0 49648 800 49768 6 Do[14]
port 47 nsew signal output
rlabel metal3 s 0 53184 800 53304 6 Do[15]
port 48 nsew signal output
rlabel metal3 s 0 56584 800 56704 6 Do[16]
port 49 nsew signal output
rlabel metal3 s 0 59984 800 60104 6 Do[17]
port 50 nsew signal output
rlabel metal3 s 0 63520 800 63640 6 Do[18]
port 51 nsew signal output
rlabel metal3 s 0 66920 800 67040 6 Do[19]
port 52 nsew signal output
rlabel metal3 s 0 5040 800 5160 6 Do[1]
port 53 nsew signal output
rlabel metal3 s 0 70320 800 70440 6 Do[20]
port 54 nsew signal output
rlabel metal3 s 0 73720 800 73840 6 Do[21]
port 55 nsew signal output
rlabel metal3 s 0 77256 800 77376 6 Do[22]
port 56 nsew signal output
rlabel metal3 s 0 80656 800 80776 6 Do[23]
port 57 nsew signal output
rlabel metal3 s 0 84056 800 84176 6 Do[24]
port 58 nsew signal output
rlabel metal3 s 0 87592 800 87712 6 Do[25]
port 59 nsew signal output
rlabel metal3 s 0 90992 800 91112 6 Do[26]
port 60 nsew signal output
rlabel metal3 s 0 94392 800 94512 6 Do[27]
port 61 nsew signal output
rlabel metal3 s 0 97792 800 97912 6 Do[28]
port 62 nsew signal output
rlabel metal3 s 0 101328 800 101448 6 Do[29]
port 63 nsew signal output
rlabel metal3 s 0 8440 800 8560 6 Do[2]
port 64 nsew signal output
rlabel metal3 s 0 104728 800 104848 6 Do[30]
port 65 nsew signal output
rlabel metal3 s 0 108128 800 108248 6 Do[31]
port 66 nsew signal output
rlabel metal3 s 0 11840 800 11960 6 Do[3]
port 67 nsew signal output
rlabel metal3 s 0 15376 800 15496 6 Do[4]
port 68 nsew signal output
rlabel metal3 s 0 18776 800 18896 6 Do[5]
port 69 nsew signal output
rlabel metal3 s 0 22176 800 22296 6 Do[6]
port 70 nsew signal output
rlabel metal3 s 0 25576 800 25696 6 Do[7]
port 71 nsew signal output
rlabel metal3 s 0 29112 800 29232 6 Do[8]
port 72 nsew signal output
rlabel metal3 s 0 32512 800 32632 6 Do[9]
port 73 nsew signal output
rlabel metal2 s 163410 109200 163466 110000 6 EN
port 74 nsew signal input
rlabel metal5 s 1104 20616 168820 20936 6 VGND
port 75 nsew ground input
rlabel metal5 s 1104 51252 168820 51572 6 VGND
port 75 nsew ground input
rlabel metal5 s 1104 81888 168820 82208 6 VGND
port 75 nsew ground input
rlabel metal4 s 19568 2128 19888 107760 6 VGND
port 75 nsew ground input
rlabel metal4 s 50288 2128 50608 107760 6 VGND
port 75 nsew ground input
rlabel metal4 s 81008 2128 81328 107760 6 VGND
port 75 nsew ground input
rlabel metal4 s 111728 2128 112048 107760 6 VGND
port 75 nsew ground input
rlabel metal4 s 142448 2128 142768 107760 6 VGND
port 75 nsew ground input
rlabel metal5 s 1104 5298 168820 5618 6 VPWR
port 76 nsew power input
rlabel metal5 s 1104 35934 168820 36254 6 VPWR
port 76 nsew power input
rlabel metal5 s 1104 66570 168820 66890 6 VPWR
port 76 nsew power input
rlabel metal5 s 1104 97206 168820 97526 6 VPWR
port 76 nsew power input
rlabel metal4 s 4208 2128 4528 107760 6 VPWR
port 76 nsew power input
rlabel metal4 s 34928 2128 35248 107760 6 VPWR
port 76 nsew power input
rlabel metal4 s 65648 2128 65968 107760 6 VPWR
port 76 nsew power input
rlabel metal4 s 96368 2128 96688 107760 6 VPWR
port 76 nsew power input
rlabel metal4 s 127088 2128 127408 107760 6 VPWR
port 76 nsew power input
rlabel metal4 s 157808 2128 158128 107760 6 VPWR
port 76 nsew power input
rlabel metal2 s 111154 109200 111210 110000 6 WE[0]
port 77 nsew signal input
rlabel metal2 s 124218 109200 124274 110000 6 WE[1]
port 78 nsew signal input
rlabel metal2 s 137282 109200 137338 110000 6 WE[2]
port 79 nsew signal input
rlabel metal2 s 150346 109200 150402 110000 6 WE[3]
port 80 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 170000 110000
string LEFview TRUE
string GDS_FILE ../gds/DFFRAM.gds
string GDS_END 63571948
string GDS_START 252880
<< end >>

