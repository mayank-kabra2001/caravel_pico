magic
tech sky130A
magscale 1 2
timestamp 1637253870
<< metal1 >>
rect 43254 162596 43260 162648
rect 43312 162636 43318 162648
rect 151906 162636 151912 162648
rect 43312 162608 151912 162636
rect 43312 162596 43318 162608
rect 151906 162596 151912 162608
rect 151964 162596 151970 162648
rect 39850 162528 39856 162580
rect 39908 162568 39914 162580
rect 149422 162568 149428 162580
rect 39908 162540 149428 162568
rect 39908 162528 39914 162540
rect 149422 162528 149428 162540
rect 149480 162528 149486 162580
rect 108850 162460 108856 162512
rect 108908 162500 108914 162512
rect 202046 162500 202052 162512
rect 108908 162472 202052 162500
rect 108908 162460 108914 162472
rect 202046 162460 202052 162472
rect 202104 162460 202110 162512
rect 102134 162392 102140 162444
rect 102192 162432 102198 162444
rect 196894 162432 196900 162444
rect 102192 162404 196900 162432
rect 102192 162392 102198 162404
rect 196894 162392 196900 162404
rect 196952 162392 196958 162444
rect 95418 162324 95424 162376
rect 95476 162364 95482 162376
rect 190730 162364 190736 162376
rect 95476 162336 190736 162364
rect 95476 162324 95482 162336
rect 190730 162324 190736 162336
rect 190788 162324 190794 162376
rect 98730 162256 98736 162308
rect 98788 162296 98794 162308
rect 193398 162296 193404 162308
rect 98788 162268 193404 162296
rect 98788 162256 98794 162268
rect 193398 162256 193404 162268
rect 193456 162256 193462 162308
rect 92014 162188 92020 162240
rect 92072 162228 92078 162240
rect 189166 162228 189172 162240
rect 92072 162200 189172 162228
rect 92072 162188 92078 162200
rect 189166 162188 189172 162200
rect 189224 162188 189230 162240
rect 88702 162120 88708 162172
rect 88760 162160 88766 162172
rect 186314 162160 186320 162172
rect 88760 162132 186320 162160
rect 88760 162120 88766 162132
rect 186314 162120 186320 162132
rect 186372 162120 186378 162172
rect 81894 162052 81900 162104
rect 81952 162092 81958 162104
rect 181070 162092 181076 162104
rect 81952 162064 181076 162092
rect 81952 162052 81958 162064
rect 181070 162052 181076 162064
rect 181128 162052 181134 162104
rect 71866 161984 71872 162036
rect 71924 162024 71930 162036
rect 172698 162024 172704 162036
rect 71924 161996 172704 162024
rect 71924 161984 71930 161996
rect 172698 161984 172704 161996
rect 172756 161984 172762 162036
rect 78582 161916 78588 161968
rect 78640 161956 78646 161968
rect 178218 161956 178224 161968
rect 78640 161928 178224 161956
rect 78640 161916 78646 161928
rect 178218 161916 178224 161928
rect 178276 161916 178282 161968
rect 75178 161848 75184 161900
rect 75236 161888 75242 161900
rect 175550 161888 175556 161900
rect 75236 161860 175556 161888
rect 75236 161848 75242 161860
rect 175550 161848 175556 161860
rect 175608 161848 175614 161900
rect 68462 161780 68468 161832
rect 68520 161820 68526 161832
rect 171318 161820 171324 161832
rect 68520 161792 171324 161820
rect 68520 161780 68526 161792
rect 171318 161780 171324 161792
rect 171376 161780 171382 161832
rect 65150 161712 65156 161764
rect 65208 161752 65214 161764
rect 168466 161752 168472 161764
rect 65208 161724 168472 161752
rect 65208 161712 65214 161724
rect 168466 161712 168472 161724
rect 168524 161712 168530 161764
rect 56686 161644 56692 161696
rect 56744 161684 56750 161696
rect 161474 161684 161480 161696
rect 56744 161656 161480 161684
rect 56744 161644 56750 161656
rect 161474 161644 161480 161656
rect 161532 161644 161538 161696
rect 61746 161576 61752 161628
rect 61804 161616 61810 161628
rect 165614 161616 165620 161628
rect 61804 161588 165620 161616
rect 61804 161576 61810 161588
rect 165614 161576 165620 161588
rect 165672 161576 165678 161628
rect 115566 161508 115572 161560
rect 115624 161548 115630 161560
rect 207014 161548 207020 161560
rect 115624 161520 207020 161548
rect 115624 161508 115630 161520
rect 207014 161508 207020 161520
rect 207072 161508 207078 161560
rect 112254 161440 112260 161492
rect 112312 161480 112318 161492
rect 204254 161480 204260 161492
rect 112312 161452 204260 161480
rect 112312 161440 112318 161452
rect 204254 161440 204260 161452
rect 204312 161440 204318 161492
rect 114738 161372 114744 161424
rect 114796 161412 114802 161424
rect 206554 161412 206560 161424
rect 114796 161384 206560 161412
rect 114796 161372 114802 161384
rect 206554 161372 206560 161384
rect 206612 161372 206618 161424
rect 108022 161304 108028 161356
rect 108080 161344 108086 161356
rect 200298 161344 200304 161356
rect 108080 161316 200304 161344
rect 108080 161304 108086 161316
rect 200298 161304 200304 161316
rect 200356 161304 200362 161356
rect 101306 161236 101312 161288
rect 101364 161276 101370 161288
rect 196250 161276 196256 161288
rect 101364 161248 196256 161276
rect 101364 161236 101370 161248
rect 196250 161236 196256 161248
rect 196308 161236 196314 161288
rect 94590 161168 94596 161220
rect 94648 161208 94654 161220
rect 191098 161208 191104 161220
rect 94648 161180 191104 161208
rect 94648 161168 94654 161180
rect 191098 161168 191104 161180
rect 191156 161168 191162 161220
rect 205542 161168 205548 161220
rect 205600 161208 205606 161220
rect 275830 161208 275836 161220
rect 205600 161180 275836 161208
rect 205600 161168 205606 161180
rect 275830 161168 275836 161180
rect 275888 161168 275894 161220
rect 81066 161100 81072 161152
rect 81124 161140 81130 161152
rect 180886 161140 180892 161152
rect 81124 161112 180892 161140
rect 81124 161100 81130 161112
rect 180886 161100 180892 161112
rect 180944 161100 180950 161152
rect 198826 161100 198832 161152
rect 198884 161140 198890 161152
rect 270494 161140 270500 161152
rect 198884 161112 270500 161140
rect 198884 161100 198890 161112
rect 270494 161100 270500 161112
rect 270552 161100 270558 161152
rect 67634 161032 67640 161084
rect 67692 161072 67698 161084
rect 169846 161072 169852 161084
rect 67692 161044 169852 161072
rect 67692 161032 67698 161044
rect 169846 161032 169852 161044
rect 169904 161032 169910 161084
rect 183738 161032 183744 161084
rect 183796 161072 183802 161084
rect 258074 161072 258080 161084
rect 183796 161044 258080 161072
rect 183796 161032 183802 161044
rect 258074 161032 258080 161044
rect 258132 161032 258138 161084
rect 60918 160964 60924 161016
rect 60976 161004 60982 161016
rect 165430 161004 165436 161016
rect 60976 160976 165436 161004
rect 60976 160964 60982 160976
rect 165430 160964 165436 160976
rect 165488 160964 165494 161016
rect 175274 160964 175280 161016
rect 175332 161004 175338 161016
rect 252738 161004 252744 161016
rect 175332 160976 252744 161004
rect 175332 160964 175338 160976
rect 252738 160964 252744 160976
rect 252796 160964 252802 161016
rect 54202 160896 54208 160948
rect 54260 160936 54266 160948
rect 160278 160936 160284 160948
rect 54260 160908 160284 160936
rect 54260 160896 54266 160908
rect 160278 160896 160284 160908
rect 160336 160896 160342 160948
rect 161842 160896 161848 160948
rect 161900 160936 161906 160948
rect 242066 160936 242072 160948
rect 161900 160908 242072 160936
rect 161900 160896 161906 160908
rect 242066 160896 242072 160908
rect 242124 160896 242130 160948
rect 47486 160828 47492 160880
rect 47544 160868 47550 160880
rect 155034 160868 155040 160880
rect 47544 160840 155040 160868
rect 47544 160828 47550 160840
rect 155034 160828 155040 160840
rect 155092 160828 155098 160880
rect 166074 160828 166080 160880
rect 166132 160868 166138 160880
rect 245746 160868 245752 160880
rect 166132 160840 245752 160868
rect 166132 160828 166138 160840
rect 245746 160828 245752 160840
rect 245804 160828 245810 160880
rect 40678 160760 40684 160812
rect 40736 160800 40742 160812
rect 149146 160800 149152 160812
rect 40736 160772 149152 160800
rect 40736 160760 40742 160772
rect 149146 160760 149152 160772
rect 149204 160760 149210 160812
rect 155126 160760 155132 160812
rect 155184 160800 155190 160812
rect 237374 160800 237380 160812
rect 155184 160772 237380 160800
rect 155184 160760 155190 160772
rect 237374 160760 237380 160772
rect 237432 160760 237438 160812
rect 36538 160692 36544 160744
rect 36596 160732 36602 160744
rect 146846 160732 146852 160744
rect 36596 160704 146852 160732
rect 36596 160692 36602 160704
rect 146846 160692 146852 160704
rect 146904 160692 146910 160744
rect 148410 160692 148416 160744
rect 148468 160732 148474 160744
rect 231946 160732 231952 160744
rect 148468 160704 231952 160732
rect 148468 160692 148474 160704
rect 231946 160692 231952 160704
rect 232004 160692 232010 160744
rect 124858 160624 124864 160676
rect 124916 160664 124922 160676
rect 213914 160664 213920 160676
rect 124916 160636 213920 160664
rect 124916 160624 124922 160636
rect 213914 160624 213920 160636
rect 213972 160624 213978 160676
rect 141694 160556 141700 160608
rect 141752 160596 141758 160608
rect 227070 160596 227076 160608
rect 141752 160568 227076 160596
rect 141752 160556 141758 160568
rect 227070 160556 227076 160568
rect 227128 160556 227134 160608
rect 149238 160488 149244 160540
rect 149296 160528 149302 160540
rect 232866 160528 232872 160540
rect 149296 160500 232872 160528
rect 149296 160488 149302 160500
rect 232866 160488 232872 160500
rect 232924 160488 232930 160540
rect 93670 160012 93676 160064
rect 93728 160052 93734 160064
rect 165522 160052 165528 160064
rect 93728 160024 165528 160052
rect 93728 160012 93734 160024
rect 165522 160012 165528 160024
rect 165580 160012 165586 160064
rect 181162 160012 181168 160064
rect 181220 160052 181226 160064
rect 230750 160052 230756 160064
rect 181220 160024 230756 160052
rect 181220 160012 181226 160024
rect 230750 160012 230756 160024
rect 230808 160012 230814 160064
rect 240870 160012 240876 160064
rect 240928 160052 240934 160064
rect 263870 160052 263876 160064
rect 240928 160024 263876 160052
rect 240928 160012 240934 160024
rect 263870 160012 263876 160024
rect 263928 160012 263934 160064
rect 265342 160012 265348 160064
rect 265400 160052 265406 160064
rect 311066 160052 311072 160064
rect 265400 160024 311072 160052
rect 265400 160012 265406 160024
rect 311066 160012 311072 160024
rect 311124 160012 311130 160064
rect 318334 160012 318340 160064
rect 318392 160052 318398 160064
rect 336642 160052 336648 160064
rect 318392 160024 336648 160052
rect 318392 160012 318398 160024
rect 336642 160012 336648 160024
rect 336700 160012 336706 160064
rect 342714 160012 342720 160064
rect 342772 160052 342778 160064
rect 372614 160052 372620 160064
rect 342772 160024 372620 160052
rect 342772 160012 342778 160024
rect 372614 160012 372620 160024
rect 372672 160012 372678 160064
rect 409138 160012 409144 160064
rect 409196 160052 409202 160064
rect 409196 160024 422294 160052
rect 409196 160012 409202 160024
rect 86954 159944 86960 159996
rect 87012 159984 87018 159996
rect 158714 159984 158720 159996
rect 87012 159956 158720 159984
rect 87012 159944 87018 159956
rect 158714 159944 158720 159956
rect 158772 159944 158778 159996
rect 164326 159944 164332 159996
rect 164384 159984 164390 159996
rect 222010 159984 222016 159996
rect 164384 159956 222016 159984
rect 164384 159944 164390 159956
rect 222010 159944 222016 159956
rect 222068 159944 222074 159996
rect 234154 159944 234160 159996
rect 234212 159984 234218 159996
rect 255498 159984 255504 159996
rect 234212 159956 255504 159984
rect 234212 159944 234218 159956
rect 255498 159944 255504 159956
rect 255556 159944 255562 159996
rect 258534 159944 258540 159996
rect 258592 159984 258598 159996
rect 304994 159984 305000 159996
rect 258592 159956 305000 159984
rect 258592 159944 258598 159956
rect 304994 159944 305000 159956
rect 305052 159944 305058 159996
rect 311526 159944 311532 159996
rect 311584 159984 311590 159996
rect 330202 159984 330208 159996
rect 311584 159956 330208 159984
rect 311584 159944 311590 159956
rect 330202 159944 330208 159956
rect 330260 159944 330266 159996
rect 332594 159944 332600 159996
rect 332652 159984 332658 159996
rect 368566 159984 368572 159996
rect 332652 159956 368572 159984
rect 332652 159944 332658 159956
rect 368566 159944 368572 159956
rect 368624 159944 368630 159996
rect 386414 159944 386420 159996
rect 386472 159984 386478 159996
rect 412818 159984 412824 159996
rect 386472 159956 412824 159984
rect 386472 159944 386478 159956
rect 412818 159944 412824 159956
rect 412876 159944 412882 159996
rect 422266 159984 422294 160024
rect 425974 160012 425980 160064
rect 426032 160052 426038 160064
rect 426434 160052 426440 160064
rect 426032 160024 426440 160052
rect 426032 160012 426038 160024
rect 426434 160012 426440 160024
rect 426492 160012 426498 160064
rect 431218 159984 431224 159996
rect 422266 159956 431224 159984
rect 431218 159944 431224 159956
rect 431276 159944 431282 159996
rect 484854 159944 484860 159996
rect 484912 159984 484918 159996
rect 488994 159984 489000 159996
rect 484912 159956 489000 159984
rect 484912 159944 484918 159956
rect 488994 159944 489000 159956
rect 489052 159944 489058 159996
rect 76926 159876 76932 159928
rect 76984 159916 76990 159928
rect 147766 159916 147772 159928
rect 76984 159888 147772 159916
rect 76984 159876 76990 159888
rect 147766 159876 147772 159888
rect 147824 159876 147830 159928
rect 150894 159876 150900 159928
rect 150952 159916 150958 159928
rect 207106 159916 207112 159928
rect 150952 159888 207112 159916
rect 150952 159876 150958 159888
rect 207106 159876 207112 159888
rect 207164 159876 207170 159928
rect 208946 159876 208952 159928
rect 209004 159916 209010 159928
rect 220170 159916 220176 159928
rect 209004 159888 220176 159916
rect 209004 159876 209010 159888
rect 220170 159876 220176 159888
rect 220228 159876 220234 159928
rect 222378 159876 222384 159928
rect 222436 159916 222442 159928
rect 225690 159916 225696 159928
rect 222436 159888 225696 159916
rect 222436 159876 222442 159888
rect 225690 159876 225696 159888
rect 225748 159876 225754 159928
rect 230382 159916 230388 159928
rect 229066 159888 230388 159916
rect 70118 159808 70124 159860
rect 70176 159848 70182 159860
rect 140866 159848 140872 159860
rect 70176 159820 140872 159848
rect 70176 159808 70182 159820
rect 140866 159808 140872 159820
rect 140924 159808 140930 159860
rect 171134 159808 171140 159860
rect 171192 159848 171198 159860
rect 229066 159848 229094 159888
rect 230382 159876 230388 159888
rect 230440 159876 230446 159928
rect 238386 159876 238392 159928
rect 238444 159916 238450 159928
rect 288250 159916 288256 159928
rect 238444 159888 288256 159916
rect 238444 159876 238450 159888
rect 288250 159876 288256 159888
rect 288308 159876 288314 159928
rect 291378 159876 291384 159928
rect 291436 159916 291442 159928
rect 311894 159916 311900 159928
rect 291436 159888 311900 159916
rect 291436 159876 291442 159888
rect 311894 159876 311900 159888
rect 311952 159876 311958 159928
rect 325878 159876 325884 159928
rect 325936 159916 325942 159928
rect 362126 159916 362132 159928
rect 325936 159888 362132 159916
rect 325936 159876 325942 159888
rect 362126 159876 362132 159888
rect 362184 159876 362190 159928
rect 393130 159876 393136 159928
rect 393188 159916 393194 159928
rect 419074 159916 419080 159928
rect 393188 159888 419080 159916
rect 393188 159876 393194 159888
rect 419074 159876 419080 159888
rect 419132 159876 419138 159928
rect 171192 159820 229094 159848
rect 171192 159808 171198 159820
rect 231670 159808 231676 159860
rect 231728 159848 231734 159860
rect 284386 159848 284392 159860
rect 231728 159820 284392 159848
rect 231728 159808 231734 159820
rect 284386 159808 284392 159820
rect 284444 159808 284450 159860
rect 305638 159808 305644 159860
rect 305696 159848 305702 159860
rect 345934 159848 345940 159860
rect 305696 159820 345940 159848
rect 305696 159808 305702 159820
rect 345934 159808 345940 159820
rect 345992 159808 345998 159860
rect 375466 159808 375472 159860
rect 375524 159848 375530 159860
rect 405550 159848 405556 159860
rect 375524 159820 405556 159848
rect 375524 159808 375530 159820
rect 405550 159808 405556 159820
rect 405608 159808 405614 159860
rect 406654 159808 406660 159860
rect 406712 159848 406718 159860
rect 429378 159848 429384 159860
rect 406712 159820 429384 159848
rect 406712 159808 406718 159820
rect 429378 159808 429384 159820
rect 429436 159808 429442 159860
rect 472250 159808 472256 159860
rect 472308 159848 472314 159860
rect 479426 159848 479432 159860
rect 472308 159820 479432 159848
rect 472308 159808 472314 159820
rect 479426 159808 479432 159820
rect 479484 159808 479490 159860
rect 46566 159740 46572 159792
rect 46624 159780 46630 159792
rect 120166 159780 120172 159792
rect 46624 159752 120172 159780
rect 46624 159740 46630 159752
rect 120166 159740 120172 159752
rect 120224 159740 120230 159792
rect 124030 159740 124036 159792
rect 124088 159780 124094 159792
rect 187694 159780 187700 159792
rect 124088 159752 187700 159780
rect 124088 159740 124094 159752
rect 187694 159740 187700 159752
rect 187752 159740 187758 159792
rect 194686 159740 194692 159792
rect 194744 159780 194750 159792
rect 212626 159780 212632 159792
rect 194744 159752 212632 159780
rect 194744 159740 194750 159752
rect 212626 159740 212632 159752
rect 212684 159740 212690 159792
rect 218238 159740 218244 159792
rect 218296 159780 218302 159792
rect 272518 159780 272524 159792
rect 218296 159752 272524 159780
rect 218296 159740 218302 159752
rect 272518 159740 272524 159752
rect 272576 159740 272582 159792
rect 277946 159740 277952 159792
rect 278004 159780 278010 159792
rect 287054 159780 287060 159792
rect 278004 159752 287060 159780
rect 278004 159740 278010 159752
rect 287054 159740 287060 159752
rect 287112 159740 287118 159792
rect 287974 159740 287980 159792
rect 288032 159780 288038 159792
rect 288618 159780 288624 159792
rect 288032 159752 288624 159780
rect 288032 159740 288038 159752
rect 288618 159740 288624 159752
rect 288676 159740 288682 159792
rect 298922 159740 298928 159792
rect 298980 159780 298986 159792
rect 343634 159780 343640 159792
rect 298980 159752 343640 159780
rect 298980 159740 298986 159752
rect 343634 159740 343640 159752
rect 343692 159740 343698 159792
rect 368750 159740 368756 159792
rect 368808 159780 368814 159792
rect 400398 159780 400404 159792
rect 368808 159752 400404 159780
rect 368808 159740 368814 159752
rect 400398 159740 400404 159752
rect 400456 159740 400462 159792
rect 402422 159740 402428 159792
rect 402480 159780 402486 159792
rect 426158 159780 426164 159792
rect 402480 159752 426164 159780
rect 402480 159740 402486 159752
rect 426158 159740 426164 159752
rect 426216 159740 426222 159792
rect 481450 159740 481456 159792
rect 481508 159780 481514 159792
rect 485774 159780 485780 159792
rect 481508 159752 485780 159780
rect 481508 159740 481514 159752
rect 485774 159740 485780 159752
rect 485832 159740 485838 159792
rect 492398 159740 492404 159792
rect 492456 159780 492462 159792
rect 494790 159780 494796 159792
rect 492456 159752 494796 159780
rect 492456 159740 492462 159752
rect 494790 159740 494796 159752
rect 494848 159740 494854 159792
rect 53374 159672 53380 159724
rect 53432 159712 53438 159724
rect 128354 159712 128360 159724
rect 53432 159684 128360 159712
rect 53432 159672 53438 159684
rect 128354 159672 128360 159684
rect 128412 159672 128418 159724
rect 130746 159672 130752 159724
rect 130804 159712 130810 159724
rect 195238 159712 195244 159724
rect 130804 159684 195244 159712
rect 130804 159672 130810 159684
rect 195238 159672 195244 159684
rect 195296 159672 195302 159724
rect 211430 159672 211436 159724
rect 211488 159712 211494 159724
rect 268930 159712 268936 159724
rect 211488 159684 268936 159712
rect 211488 159672 211494 159684
rect 268930 159672 268936 159684
rect 268988 159672 268994 159724
rect 282086 159672 282092 159724
rect 282144 159712 282150 159724
rect 291102 159712 291108 159724
rect 282144 159684 291108 159712
rect 282144 159672 282150 159684
rect 291102 159672 291108 159684
rect 291160 159672 291166 159724
rect 292206 159672 292212 159724
rect 292264 159712 292270 159724
rect 338390 159712 338396 159724
rect 292264 159684 338396 159712
rect 292264 159672 292270 159684
rect 338390 159672 338396 159684
rect 338448 159672 338454 159724
rect 346026 159672 346032 159724
rect 346084 159712 346090 159724
rect 378318 159712 378324 159724
rect 346084 159684 378324 159712
rect 346084 159672 346090 159684
rect 378318 159672 378324 159684
rect 378376 159672 378382 159724
rect 382182 159672 382188 159724
rect 382240 159712 382246 159724
rect 408494 159712 408500 159724
rect 382240 159684 408500 159712
rect 382240 159672 382246 159684
rect 408494 159672 408500 159684
rect 408552 159672 408558 159724
rect 413370 159672 413376 159724
rect 413428 159712 413434 159724
rect 434438 159712 434444 159724
rect 413428 159684 434444 159712
rect 413428 159672 413434 159684
rect 434438 159672 434444 159684
rect 434496 159672 434502 159724
rect 478966 159672 478972 159724
rect 479024 159712 479030 159724
rect 484394 159712 484400 159724
rect 479024 159684 484400 159712
rect 479024 159672 479030 159684
rect 484394 159672 484400 159684
rect 484452 159672 484458 159724
rect 3694 159604 3700 159656
rect 3752 159644 3758 159656
rect 77202 159644 77208 159656
rect 3752 159616 77208 159644
rect 3752 159604 3758 159616
rect 77202 159604 77208 159616
rect 77260 159604 77266 159656
rect 80238 159604 80244 159656
rect 80296 159644 80302 159656
rect 156046 159644 156052 159656
rect 80296 159616 156052 159644
rect 80296 159604 80302 159616
rect 156046 159604 156052 159616
rect 156104 159604 156110 159656
rect 157610 159604 157616 159656
rect 157668 159644 157674 159656
rect 216858 159644 216864 159656
rect 157668 159616 216864 159644
rect 157668 159604 157674 159616
rect 216858 159604 216864 159616
rect 216916 159604 216922 159656
rect 224954 159604 224960 159656
rect 225012 159644 225018 159656
rect 281166 159644 281172 159656
rect 225012 159616 281172 159644
rect 225012 159604 225018 159616
rect 281166 159604 281172 159616
rect 281224 159604 281230 159656
rect 285490 159604 285496 159656
rect 285548 159644 285554 159656
rect 332594 159644 332600 159656
rect 285548 159616 332600 159644
rect 285548 159604 285554 159616
rect 332594 159604 332600 159616
rect 332652 159604 332658 159656
rect 352742 159604 352748 159656
rect 352800 159644 352806 159656
rect 385954 159644 385960 159656
rect 352800 159616 385960 159644
rect 352800 159604 352806 159616
rect 385954 159604 385960 159616
rect 386012 159604 386018 159656
rect 388990 159604 388996 159656
rect 389048 159644 389054 159656
rect 414290 159644 414296 159656
rect 389048 159616 414296 159644
rect 389048 159604 389054 159616
rect 414290 159604 414296 159616
rect 414348 159604 414354 159656
rect 420086 159604 420092 159656
rect 420144 159644 420150 159656
rect 435818 159644 435824 159656
rect 420144 159616 435824 159644
rect 420144 159604 420150 159616
rect 435818 159604 435824 159616
rect 435876 159604 435882 159656
rect 441062 159604 441068 159656
rect 441120 159644 441126 159656
rect 445478 159644 445484 159656
rect 441120 159616 445484 159644
rect 441120 159604 441126 159616
rect 445478 159604 445484 159616
rect 445536 159604 445542 159656
rect 478138 159604 478144 159656
rect 478196 159644 478202 159656
rect 483014 159644 483020 159656
rect 478196 159616 483020 159644
rect 478196 159604 478202 159616
rect 483014 159604 483020 159616
rect 483072 159604 483078 159656
rect 33962 159536 33968 159588
rect 34020 159576 34026 159588
rect 63494 159576 63500 159588
rect 34020 159548 63500 159576
rect 34020 159536 34026 159548
rect 63494 159536 63500 159548
rect 63552 159536 63558 159588
rect 66806 159536 66812 159588
rect 66864 159576 66870 159588
rect 144822 159576 144828 159588
rect 66864 159548 144828 159576
rect 66864 159536 66870 159548
rect 144822 159536 144828 159548
rect 144880 159536 144886 159588
rect 170214 159536 170220 159588
rect 170272 159576 170278 159588
rect 176654 159576 176660 159588
rect 170272 159548 176660 159576
rect 170272 159536 170278 159548
rect 176654 159536 176660 159548
rect 176712 159536 176718 159588
rect 197998 159536 198004 159588
rect 198056 159576 198062 159588
rect 260742 159576 260748 159588
rect 198056 159548 260748 159576
rect 198056 159536 198062 159548
rect 260742 159536 260748 159548
rect 260800 159536 260806 159588
rect 272058 159536 272064 159588
rect 272116 159576 272122 159588
rect 320726 159576 320732 159588
rect 272116 159548 320732 159576
rect 272116 159536 272122 159548
rect 320726 159536 320732 159548
rect 320784 159536 320790 159588
rect 339310 159536 339316 159588
rect 339368 159576 339374 159588
rect 377950 159576 377956 159588
rect 339368 159548 377956 159576
rect 339368 159536 339374 159548
rect 377950 159536 377956 159548
rect 378008 159536 378014 159588
rect 379698 159536 379704 159588
rect 379756 159576 379762 159588
rect 408770 159576 408776 159588
rect 379756 159548 408776 159576
rect 379756 159536 379762 159548
rect 408770 159536 408776 159548
rect 408828 159536 408834 159588
rect 431862 159536 431868 159588
rect 431920 159576 431926 159588
rect 436554 159576 436560 159588
rect 431920 159548 436560 159576
rect 431920 159536 431926 159548
rect 436554 159536 436560 159548
rect 436612 159536 436618 159588
rect 2866 159468 2872 159520
rect 2924 159508 2930 159520
rect 92474 159508 92480 159520
rect 2924 159480 92480 159508
rect 2924 159468 2930 159480
rect 92474 159468 92480 159480
rect 92532 159468 92538 159520
rect 100478 159468 100484 159520
rect 100536 159508 100542 159520
rect 169754 159508 169760 159520
rect 100536 159480 169760 159508
rect 100536 159468 100542 159480
rect 169754 159468 169760 159480
rect 169812 159468 169818 159520
rect 184566 159468 184572 159520
rect 184624 159508 184630 159520
rect 247218 159508 247224 159520
rect 184624 159480 247224 159508
rect 184624 159468 184630 159480
rect 247218 159468 247224 159480
rect 247276 159468 247282 159520
rect 251818 159468 251824 159520
rect 251876 159508 251882 159520
rect 301682 159508 301688 159520
rect 251876 159480 301688 159508
rect 251876 159468 251882 159480
rect 301682 159468 301688 159480
rect 301740 159468 301746 159520
rect 308214 159468 308220 159520
rect 308272 159508 308278 159520
rect 317782 159508 317788 159520
rect 308272 159480 317788 159508
rect 308272 159468 308278 159480
rect 317782 159468 317788 159480
rect 317840 159468 317846 159520
rect 319162 159468 319168 159520
rect 319220 159508 319226 159520
rect 361574 159508 361580 159520
rect 319220 159480 361580 159508
rect 319220 159468 319226 159480
rect 361574 159468 361580 159480
rect 361632 159468 361638 159520
rect 366266 159468 366272 159520
rect 366324 159508 366330 159520
rect 398466 159508 398472 159520
rect 366324 159480 398472 159508
rect 366324 159468 366330 159480
rect 398466 159468 398472 159480
rect 398524 159468 398530 159520
rect 399846 159468 399852 159520
rect 399904 159508 399910 159520
rect 424226 159508 424232 159520
rect 399904 159480 424232 159508
rect 399904 159468 399910 159480
rect 424226 159468 424232 159480
rect 424284 159468 424290 159520
rect 433518 159468 433524 159520
rect 433576 159508 433582 159520
rect 449802 159508 449808 159520
rect 433576 159480 449808 159508
rect 433576 159468 433582 159480
rect 449802 159468 449808 159480
rect 449860 159468 449866 159520
rect 451182 159468 451188 159520
rect 451240 159508 451246 159520
rect 455322 159508 455328 159520
rect 451240 159480 455328 159508
rect 451240 159468 451246 159480
rect 455322 159468 455328 159480
rect 455380 159468 455386 159520
rect 26418 159400 26424 159452
rect 26476 159440 26482 159452
rect 129826 159440 129832 159452
rect 26476 159412 129832 159440
rect 26476 159400 26482 159412
rect 129826 159400 129832 159412
rect 129884 159400 129890 159452
rect 139118 159400 139124 159452
rect 139176 159440 139182 159452
rect 157426 159440 157432 159452
rect 139176 159412 157432 159440
rect 139176 159400 139182 159412
rect 157426 159400 157432 159412
rect 157484 159400 157490 159452
rect 177850 159400 177856 159452
rect 177908 159440 177914 159452
rect 242434 159440 242440 159452
rect 177908 159412 242440 159440
rect 177908 159400 177914 159412
rect 242434 159400 242440 159412
rect 242492 159400 242498 159452
rect 245102 159400 245108 159452
rect 245160 159440 245166 159452
rect 299382 159440 299388 159452
rect 245160 159412 299388 159440
rect 245160 159400 245166 159412
rect 299382 159400 299388 159412
rect 299440 159400 299446 159452
rect 312446 159400 312452 159452
rect 312504 159440 312510 159452
rect 355686 159440 355692 159452
rect 312504 159412 355692 159440
rect 312504 159400 312510 159412
rect 355686 159400 355692 159412
rect 355744 159400 355750 159452
rect 359550 159400 359556 159452
rect 359608 159440 359614 159452
rect 393406 159440 393412 159452
rect 359608 159412 393412 159440
rect 359608 159400 359614 159412
rect 393406 159400 393412 159412
rect 393464 159400 393470 159452
rect 395706 159400 395712 159452
rect 395764 159440 395770 159452
rect 421098 159440 421104 159452
rect 395764 159412 421104 159440
rect 395764 159400 395770 159412
rect 421098 159400 421104 159412
rect 421156 159400 421162 159452
rect 432690 159400 432696 159452
rect 432748 159440 432754 159452
rect 447134 159440 447140 159452
rect 432748 159412 447140 159440
rect 432748 159400 432754 159412
rect 447134 159400 447140 159412
rect 447192 159400 447198 159452
rect 479794 159400 479800 159452
rect 479852 159440 479858 159452
rect 485222 159440 485228 159452
rect 479852 159412 485228 159440
rect 479852 159400 479858 159412
rect 485222 159400 485228 159412
rect 485280 159400 485286 159452
rect 496630 159400 496636 159452
rect 496688 159440 496694 159452
rect 498010 159440 498016 159452
rect 496688 159412 498016 159440
rect 496688 159400 496694 159412
rect 498010 159400 498016 159412
rect 498068 159400 498074 159452
rect 12986 159332 12992 159384
rect 13044 159372 13050 159384
rect 124122 159372 124128 159384
rect 13044 159344 124128 159372
rect 13044 159332 13050 159344
rect 124122 159332 124128 159344
rect 124180 159332 124186 159384
rect 132402 159332 132408 159384
rect 132460 159372 132466 159384
rect 135806 159372 135812 159384
rect 132460 159344 135812 159372
rect 132460 159332 132466 159344
rect 135806 159332 135812 159344
rect 135864 159332 135870 159384
rect 140774 159332 140780 159384
rect 140832 159372 140838 159384
rect 174906 159372 174912 159384
rect 140832 159344 174912 159372
rect 140832 159332 140838 159344
rect 174906 159332 174912 159344
rect 174964 159332 174970 159384
rect 191282 159332 191288 159384
rect 191340 159372 191346 159384
rect 256786 159372 256792 159384
rect 191340 159344 256792 159372
rect 191340 159332 191346 159344
rect 256786 159332 256792 159344
rect 256844 159332 256850 159384
rect 261938 159332 261944 159384
rect 261996 159372 262002 159384
rect 263502 159372 263508 159384
rect 261996 159344 263508 159372
rect 261996 159332 262002 159344
rect 263502 159332 263508 159344
rect 263560 159332 263566 159384
rect 287054 159332 287060 159384
rect 287112 159372 287118 159384
rect 291470 159372 291476 159384
rect 287112 159344 291476 159372
rect 287112 159332 287118 159344
rect 291470 159332 291476 159344
rect 291528 159332 291534 159384
rect 331766 159332 331772 159384
rect 331824 159372 331830 159384
rect 372062 159372 372068 159384
rect 331824 159344 372068 159372
rect 331824 159332 331830 159344
rect 372062 159332 372068 159344
rect 372120 159332 372126 159384
rect 372982 159332 372988 159384
rect 373040 159372 373046 159384
rect 403158 159372 403164 159384
rect 373040 159344 403164 159372
rect 373040 159332 373046 159344
rect 403158 159332 403164 159344
rect 403216 159332 403222 159384
rect 434346 159332 434352 159384
rect 434404 159372 434410 159384
rect 450078 159372 450084 159384
rect 434404 159344 450084 159372
rect 434404 159332 434410 159344
rect 450078 159332 450084 159344
rect 450136 159332 450142 159384
rect 461302 159332 461308 159384
rect 461360 159372 461366 159384
rect 464890 159372 464896 159384
rect 461360 159344 464896 159372
rect 461360 159332 461366 159344
rect 464890 159332 464896 159344
rect 464948 159332 464954 159384
rect 477310 159332 477316 159384
rect 477368 159372 477374 159384
rect 483290 159372 483296 159384
rect 477368 159344 483296 159372
rect 477368 159332 477374 159344
rect 483290 159332 483296 159344
rect 483348 159332 483354 159384
rect 497458 159332 497464 159384
rect 497516 159372 497522 159384
rect 498654 159372 498660 159384
rect 497516 159344 498660 159372
rect 497516 159332 497522 159344
rect 498654 159332 498660 159344
rect 498712 159332 498718 159384
rect 49970 159264 49976 159316
rect 50028 159304 50034 159316
rect 109218 159304 109224 159316
rect 50028 159276 109224 159304
rect 50028 159264 50034 159276
rect 109218 159264 109224 159276
rect 109276 159264 109282 159316
rect 110506 159264 110512 159316
rect 110564 159304 110570 159316
rect 179414 159304 179420 159316
rect 110564 159276 179420 159304
rect 110564 159264 110570 159276
rect 179414 159264 179420 159276
rect 179472 159264 179478 159316
rect 187878 159264 187884 159316
rect 187936 159304 187942 159316
rect 210878 159304 210884 159316
rect 187936 159276 210884 159304
rect 187936 159264 187942 159276
rect 210878 159264 210884 159276
rect 210936 159264 210942 159316
rect 214834 159264 214840 159316
rect 214892 159304 214898 159316
rect 223942 159304 223948 159316
rect 214892 159276 223948 159304
rect 214892 159264 214898 159276
rect 223942 159264 223948 159276
rect 224000 159264 224006 159316
rect 227438 159264 227444 159316
rect 227496 159304 227502 159316
rect 247034 159304 247040 159316
rect 227496 159276 247040 159304
rect 227496 159264 227502 159276
rect 247034 159264 247040 159276
rect 247092 159264 247098 159316
rect 261110 159264 261116 159316
rect 261168 159304 261174 159316
rect 269022 159304 269028 159316
rect 261168 159276 269028 159304
rect 261168 159264 261174 159276
rect 269022 159264 269028 159276
rect 269080 159264 269086 159316
rect 271230 159264 271236 159316
rect 271288 159304 271294 159316
rect 296806 159304 296812 159316
rect 271288 159276 296812 159304
rect 271288 159264 271294 159276
rect 296806 159264 296812 159276
rect 296864 159264 296870 159316
rect 298094 159264 298100 159316
rect 298152 159304 298158 159316
rect 311986 159304 311992 159316
rect 298152 159276 311992 159304
rect 298152 159264 298158 159276
rect 311986 159264 311992 159276
rect 312044 159264 312050 159316
rect 325050 159264 325056 159316
rect 325108 159304 325114 159316
rect 352006 159304 352012 159316
rect 325108 159276 352012 159304
rect 325108 159264 325114 159276
rect 352006 159264 352012 159276
rect 352064 159264 352070 159316
rect 480622 159264 480628 159316
rect 480680 159304 480686 159316
rect 485866 159304 485872 159316
rect 480680 159276 485872 159304
rect 480680 159264 480686 159276
rect 485866 159264 485872 159276
rect 485924 159264 485930 159316
rect 494974 159264 494980 159316
rect 495032 159304 495038 159316
rect 496722 159304 496728 159316
rect 495032 159276 496728 159304
rect 495032 159264 495038 159276
rect 496722 159264 496728 159276
rect 496780 159264 496786 159316
rect 76006 159196 76012 159248
rect 76064 159236 76070 159248
rect 79962 159236 79968 159248
rect 76064 159208 79968 159236
rect 76064 159196 76070 159208
rect 79962 159196 79968 159208
rect 80020 159196 80026 159248
rect 120626 159196 120632 159248
rect 120684 159236 120690 159248
rect 184842 159236 184848 159248
rect 120684 159208 184848 159236
rect 120684 159196 120690 159208
rect 184842 159196 184848 159208
rect 184900 159196 184906 159248
rect 208118 159196 208124 159248
rect 208176 159236 208182 159248
rect 222102 159236 222108 159248
rect 208176 159208 222108 159236
rect 208176 159196 208182 159208
rect 222102 159196 222108 159208
rect 222160 159196 222166 159248
rect 228266 159196 228272 159248
rect 228324 159236 228330 159248
rect 239950 159236 239956 159248
rect 228324 159208 239956 159236
rect 228324 159196 228330 159208
rect 239950 159196 239956 159208
rect 240008 159196 240014 159248
rect 250990 159196 250996 159248
rect 251048 159236 251054 159248
rect 274634 159236 274640 159248
rect 251048 159208 274640 159236
rect 251048 159196 251054 159208
rect 274634 159196 274640 159208
rect 274692 159196 274698 159248
rect 284662 159196 284668 159248
rect 284720 159236 284726 159248
rect 305454 159236 305460 159248
rect 284720 159208 305460 159236
rect 284720 159196 284726 159208
rect 305454 159196 305460 159208
rect 305512 159196 305518 159248
rect 489914 159196 489920 159248
rect 489972 159236 489978 159248
rect 492674 159236 492680 159248
rect 489972 159208 492680 159236
rect 489972 159196 489978 159208
rect 492674 159196 492680 159208
rect 492732 159196 492738 159248
rect 37366 159128 37372 159180
rect 37424 159168 37430 159180
rect 38562 159168 38568 159180
rect 37424 159140 38568 159168
rect 37424 159128 37430 159140
rect 38562 159128 38568 159140
rect 38620 159128 38626 159180
rect 127342 159128 127348 159180
rect 127400 159168 127406 159180
rect 143074 159168 143080 159180
rect 127400 159140 143080 159168
rect 127400 159128 127406 159140
rect 143074 159128 143080 159140
rect 143132 159128 143138 159180
rect 144178 159128 144184 159180
rect 144236 159168 144242 159180
rect 193122 159168 193128 159180
rect 144236 159140 193128 159168
rect 144236 159128 144242 159140
rect 193122 159128 193128 159140
rect 193180 159128 193186 159180
rect 201402 159128 201408 159180
rect 201460 159168 201466 159180
rect 212350 159168 212356 159180
rect 201460 159140 212356 159168
rect 201460 159128 201466 159140
rect 212350 159128 212356 159140
rect 212408 159128 212414 159180
rect 237558 159128 237564 159180
rect 237616 159168 237622 159180
rect 251726 159168 251732 159180
rect 237616 159140 251732 159168
rect 237616 159128 237622 159140
rect 251726 159128 251732 159140
rect 251784 159128 251790 159180
rect 257706 159128 257712 159180
rect 257764 159168 257770 159180
rect 279878 159168 279884 159180
rect 257764 159140 279884 159168
rect 257764 159128 257770 159140
rect 279878 159128 279884 159140
rect 279936 159128 279942 159180
rect 304810 159128 304816 159180
rect 304868 159168 304874 159180
rect 324314 159168 324320 159180
rect 304868 159140 324320 159168
rect 304868 159128 304874 159140
rect 324314 159128 324320 159140
rect 324372 159128 324378 159180
rect 493226 159128 493232 159180
rect 493284 159168 493290 159180
rect 495434 159168 495440 159180
rect 493284 159140 495440 159168
rect 493284 159128 493290 159140
rect 495434 159128 495440 159140
rect 495492 159128 495498 159180
rect 91186 159060 91192 159112
rect 91244 159100 91250 159112
rect 92382 159100 92388 159112
rect 91244 159072 92388 159100
rect 91244 159060 91250 159072
rect 92382 159060 92388 159072
rect 92440 159060 92446 159112
rect 155954 159060 155960 159112
rect 156012 159100 156018 159112
rect 197354 159100 197360 159112
rect 156012 159072 197360 159100
rect 156012 159060 156018 159072
rect 197354 159060 197360 159072
rect 197412 159060 197418 159112
rect 214006 159060 214012 159112
rect 214064 159100 214070 159112
rect 216674 159100 216680 159112
rect 214064 159072 216680 159100
rect 214064 159060 214070 159072
rect 216674 159060 216680 159072
rect 216732 159060 216738 159112
rect 217318 159060 217324 159112
rect 217376 159100 217382 159112
rect 223482 159100 223488 159112
rect 217376 159072 223488 159100
rect 217376 159060 217382 159072
rect 223482 159060 223488 159072
rect 223540 159060 223546 159112
rect 247678 159060 247684 159112
rect 247736 159100 247742 159112
rect 262122 159100 262128 159112
rect 247736 159072 262128 159100
rect 247736 159060 247742 159072
rect 262122 159060 262128 159072
rect 262180 159060 262186 159112
rect 264422 159060 264428 159112
rect 264480 159100 264486 159112
rect 284294 159100 284300 159112
rect 264480 159072 284300 159100
rect 264480 159060 264486 159072
rect 284294 159060 284300 159072
rect 284352 159060 284358 159112
rect 426802 159060 426808 159112
rect 426860 159100 426866 159112
rect 433058 159100 433064 159112
rect 426860 159072 433064 159100
rect 426860 159060 426866 159072
rect 433058 159060 433064 159072
rect 433116 159060 433122 159112
rect 471422 159060 471428 159112
rect 471480 159100 471486 159112
rect 477678 159100 477684 159112
rect 471480 159072 477684 159100
rect 471480 159060 471486 159072
rect 477678 159060 477684 159072
rect 477736 159060 477742 159112
rect 484026 159060 484032 159112
rect 484084 159100 484090 159112
rect 488442 159100 488448 159112
rect 484084 159072 488448 159100
rect 484084 159060 484090 159072
rect 488442 159060 488448 159072
rect 488500 159060 488506 159112
rect 174446 158992 174452 159044
rect 174504 159032 174510 159044
rect 204162 159032 204168 159044
rect 174504 159004 204168 159032
rect 174504 158992 174510 159004
rect 204162 158992 204168 159004
rect 204220 158992 204226 159044
rect 210602 158992 210608 159044
rect 210660 159032 210666 159044
rect 215018 159032 215024 159044
rect 210660 159004 215024 159032
rect 210660 158992 210666 159004
rect 215018 158992 215024 159004
rect 215076 158992 215082 159044
rect 267826 158992 267832 159044
rect 267884 159032 267890 159044
rect 279510 159032 279516 159044
rect 267884 159004 279516 159032
rect 267884 158992 267890 159004
rect 279510 158992 279516 159004
rect 279568 158992 279574 159044
rect 390646 158992 390652 159044
rect 390704 159032 390710 159044
rect 391842 159032 391848 159044
rect 390704 159004 391848 159032
rect 390704 158992 390710 159004
rect 391842 158992 391848 159004
rect 391900 158992 391906 159044
rect 453758 158992 453764 159044
rect 453816 159032 453822 159044
rect 458174 159032 458180 159044
rect 453816 159004 458180 159032
rect 453816 158992 453822 159004
rect 458174 158992 458180 159004
rect 458232 158992 458238 159044
rect 473078 158992 473084 159044
rect 473136 159032 473142 159044
rect 478966 159032 478972 159044
rect 473136 159004 478972 159032
rect 473136 158992 473142 159004
rect 478966 158992 478972 159004
rect 479024 158992 479030 159044
rect 486510 158992 486516 159044
rect 486568 159032 486574 159044
rect 490282 159032 490288 159044
rect 486568 159004 490288 159032
rect 486568 158992 486574 159004
rect 490282 158992 490288 159004
rect 490340 158992 490346 159044
rect 118970 158924 118976 158976
rect 119028 158964 119034 158976
rect 125502 158964 125508 158976
rect 119028 158936 125508 158964
rect 119028 158924 119034 158936
rect 125502 158924 125508 158936
rect 125560 158924 125566 158976
rect 224126 158924 224132 158976
rect 224184 158964 224190 158976
rect 227714 158964 227720 158976
rect 224184 158936 227720 158964
rect 224184 158924 224190 158936
rect 227714 158924 227720 158936
rect 227772 158924 227778 158976
rect 278774 158924 278780 158976
rect 278832 158964 278838 158976
rect 278832 158936 316034 158964
rect 278832 158924 278838 158936
rect 275370 158856 275376 158908
rect 275428 158896 275434 158908
rect 278682 158896 278688 158908
rect 275428 158868 278688 158896
rect 275428 158856 275434 158868
rect 278682 158856 278688 158868
rect 278740 158856 278746 158908
rect 316006 158896 316034 158936
rect 327534 158924 327540 158976
rect 327592 158964 327598 158976
rect 328362 158964 328368 158976
rect 327592 158936 328368 158964
rect 327592 158924 327598 158936
rect 328362 158924 328368 158936
rect 328420 158924 328426 158976
rect 362034 158924 362040 158976
rect 362092 158964 362098 158976
rect 366818 158964 366824 158976
rect 362092 158936 366824 158964
rect 362092 158924 362098 158936
rect 366818 158924 366824 158936
rect 366876 158924 366882 158976
rect 372154 158924 372160 158976
rect 372212 158964 372218 158976
rect 374270 158964 374276 158976
rect 372212 158936 374276 158964
rect 372212 158924 372218 158936
rect 374270 158924 374276 158936
rect 374328 158924 374334 158976
rect 437750 158924 437756 158976
rect 437808 158964 437814 158976
rect 444282 158964 444288 158976
rect 437808 158936 444288 158964
rect 437808 158924 437814 158936
rect 444282 158924 444288 158936
rect 444340 158924 444346 158976
rect 447870 158924 447876 158976
rect 447928 158964 447934 158976
rect 452470 158964 452476 158976
rect 447928 158936 452476 158964
rect 447928 158924 447934 158936
rect 452470 158924 452476 158936
rect 452528 158924 452534 158976
rect 463786 158924 463792 158976
rect 463844 158964 463850 158976
rect 471790 158964 471796 158976
rect 463844 158936 471796 158964
rect 463844 158924 463850 158936
rect 471790 158924 471796 158936
rect 471848 158924 471854 158976
rect 475562 158924 475568 158976
rect 475620 158964 475626 158976
rect 481634 158964 481640 158976
rect 475620 158936 481640 158964
rect 475620 158924 475626 158936
rect 481634 158924 481640 158936
rect 481692 158924 481698 158976
rect 487338 158924 487344 158976
rect 487396 158964 487402 158976
rect 489914 158964 489920 158976
rect 487396 158936 489920 158964
rect 487396 158924 487402 158936
rect 489914 158924 489920 158936
rect 489972 158924 489978 158976
rect 491570 158924 491576 158976
rect 491628 158964 491634 158976
rect 494146 158964 494152 158976
rect 491628 158936 494152 158964
rect 491628 158924 491634 158936
rect 494146 158924 494152 158936
rect 494204 158924 494210 158976
rect 331766 158896 331772 158908
rect 316006 158868 331772 158896
rect 331766 158856 331772 158868
rect 331824 158856 331830 158908
rect 473906 158856 473912 158908
rect 473964 158896 473970 158908
rect 480254 158896 480260 158908
rect 473964 158868 480260 158896
rect 473964 158856 473970 158868
rect 480254 158856 480260 158868
rect 480312 158856 480318 158908
rect 482278 158856 482284 158908
rect 482336 158896 482342 158908
rect 487154 158896 487160 158908
rect 482336 158868 487160 158896
rect 482336 158856 482342 158868
rect 487154 158856 487160 158868
rect 487212 158856 487218 158908
rect 489086 158856 489092 158908
rect 489144 158896 489150 158908
rect 491294 158896 491300 158908
rect 489144 158868 491300 158896
rect 489144 158856 489150 158868
rect 491294 158856 491300 158868
rect 491352 158856 491358 158908
rect 121454 158788 121460 158840
rect 121512 158828 121518 158840
rect 122742 158828 122748 158840
rect 121512 158800 122748 158828
rect 121512 158788 121518 158800
rect 122742 158788 122748 158800
rect 122800 158788 122806 158840
rect 128998 158788 129004 158840
rect 129056 158828 129062 158840
rect 132126 158828 132132 158840
rect 129056 158800 132132 158828
rect 129056 158788 129062 158800
rect 132126 158788 132132 158800
rect 132184 158788 132190 158840
rect 145834 158788 145840 158840
rect 145892 158828 145898 158840
rect 150434 158828 150440 158840
rect 145892 158800 150440 158828
rect 145892 158788 145898 158800
rect 150434 158788 150440 158800
rect 150492 158788 150498 158840
rect 241790 158788 241796 158840
rect 241848 158828 241854 158840
rect 244550 158828 244556 158840
rect 241848 158800 244556 158828
rect 241848 158788 241854 158800
rect 244550 158788 244556 158800
rect 244608 158788 244614 158840
rect 315758 158788 315764 158840
rect 315816 158828 315822 158840
rect 318702 158828 318708 158840
rect 315816 158800 318708 158828
rect 315816 158788 315822 158800
rect 318702 158788 318708 158800
rect 318760 158788 318766 158840
rect 378870 158788 378876 158840
rect 378928 158828 378934 158840
rect 380986 158828 380992 158840
rect 378928 158800 380992 158828
rect 378928 158788 378934 158800
rect 380986 158788 380992 158800
rect 381044 158788 381050 158840
rect 389818 158788 389824 158840
rect 389876 158828 389882 158840
rect 391566 158828 391572 158840
rect 389876 158800 391572 158828
rect 389876 158788 389882 158800
rect 391566 158788 391572 158800
rect 391624 158788 391630 158840
rect 405734 158788 405740 158840
rect 405792 158828 405798 158840
rect 406930 158828 406936 158840
rect 405792 158800 406936 158828
rect 405792 158788 405798 158800
rect 406930 158788 406936 158800
rect 406988 158788 406994 158840
rect 436094 158788 436100 158840
rect 436152 158828 436158 158840
rect 438854 158828 438860 158840
rect 436152 158800 438860 158828
rect 436152 158788 436158 158800
rect 438854 158788 438860 158800
rect 438912 158788 438918 158840
rect 449526 158788 449532 158840
rect 449584 158828 449590 158840
rect 453942 158828 453948 158840
rect 449584 158800 453948 158828
rect 449584 158788 449590 158800
rect 453942 158788 453948 158800
rect 454000 158788 454006 158840
rect 474734 158788 474740 158840
rect 474792 158828 474798 158840
rect 481358 158828 481364 158840
rect 474792 158800 481364 158828
rect 474792 158788 474798 158800
rect 481358 158788 481364 158800
rect 481416 158788 481422 158840
rect 483198 158788 483204 158840
rect 483256 158828 483262 158840
rect 487522 158828 487528 158840
rect 483256 158800 487528 158828
rect 483256 158788 483262 158800
rect 487522 158788 487528 158800
rect 487580 158788 487586 158840
rect 488166 158788 488172 158840
rect 488224 158828 488230 158840
rect 491570 158828 491576 158840
rect 488224 158800 491576 158828
rect 488224 158788 488230 158800
rect 491570 158788 491576 158800
rect 491628 158788 491634 158840
rect 382 158720 388 158772
rect 440 158760 446 158772
rect 2038 158760 2044 158772
rect 440 158732 2044 158760
rect 440 158720 446 158732
rect 2038 158720 2044 158732
rect 2096 158720 2102 158772
rect 64230 158720 64236 158772
rect 64288 158760 64294 158772
rect 64782 158760 64788 158772
rect 64288 158732 64788 158760
rect 64288 158720 64294 158732
rect 64782 158720 64788 158732
rect 64840 158720 64846 158772
rect 65978 158720 65984 158772
rect 66036 158760 66042 158772
rect 66036 158732 66300 158760
rect 66036 158720 66042 158732
rect 66272 158692 66300 158732
rect 71038 158720 71044 158772
rect 71096 158760 71102 158772
rect 71682 158760 71688 158772
rect 71096 158732 71688 158760
rect 71096 158720 71102 158732
rect 71682 158720 71688 158732
rect 71740 158720 71746 158772
rect 77754 158720 77760 158772
rect 77812 158760 77818 158772
rect 78582 158760 78588 158772
rect 77812 158732 78588 158760
rect 77812 158720 77818 158732
rect 78582 158720 78588 158732
rect 78640 158720 78646 158772
rect 84470 158720 84476 158772
rect 84528 158760 84534 158772
rect 85482 158760 85488 158772
rect 84528 158732 85488 158760
rect 84528 158720 84534 158732
rect 85482 158720 85488 158732
rect 85540 158720 85546 158772
rect 103790 158720 103796 158772
rect 103848 158760 103854 158772
rect 109034 158760 109040 158772
rect 103848 158732 109040 158760
rect 103848 158720 103854 158732
rect 109034 158720 109040 158732
rect 109092 158720 109098 158772
rect 116394 158720 116400 158772
rect 116452 158760 116458 158772
rect 119522 158760 119528 158772
rect 116452 158732 119528 158760
rect 116452 158720 116458 158732
rect 119522 158720 119528 158732
rect 119580 158720 119586 158772
rect 131574 158720 131580 158772
rect 131632 158760 131638 158772
rect 132402 158760 132408 158772
rect 131632 158732 132408 158760
rect 131632 158720 131638 158732
rect 132402 158720 132408 158732
rect 132460 158720 132466 158772
rect 145006 158720 145012 158772
rect 145064 158760 145070 158772
rect 146202 158760 146208 158772
rect 145064 158732 146208 158760
rect 145064 158720 145070 158732
rect 146202 158720 146208 158732
rect 146260 158720 146266 158772
rect 152550 158720 152556 158772
rect 152608 158760 152614 158772
rect 153102 158760 153108 158772
rect 152608 158732 153108 158760
rect 152608 158720 152614 158732
rect 153102 158720 153108 158732
rect 153160 158720 153166 158772
rect 165246 158720 165252 158772
rect 165304 158760 165310 158772
rect 167638 158760 167644 158772
rect 165304 158732 167644 158760
rect 165304 158720 165310 158732
rect 167638 158720 167644 158732
rect 167696 158720 167702 158772
rect 196342 158720 196348 158772
rect 196400 158760 196406 158772
rect 198734 158760 198740 158772
rect 196400 158732 198740 158760
rect 196400 158720 196406 158732
rect 198734 158720 198740 158732
rect 198792 158720 198798 158772
rect 202230 158720 202236 158772
rect 202288 158760 202294 158772
rect 202782 158760 202788 158772
rect 202288 158732 202788 158760
rect 202288 158720 202294 158732
rect 202782 158720 202788 158732
rect 202840 158720 202846 158772
rect 203058 158720 203064 158772
rect 203116 158760 203122 158772
rect 208486 158760 208492 158772
rect 203116 158732 208492 158760
rect 203116 158720 203122 158732
rect 208486 158720 208492 158732
rect 208544 158720 208550 158772
rect 220722 158720 220728 158772
rect 220780 158760 220786 158772
rect 227898 158760 227904 158772
rect 220780 158732 227904 158760
rect 220780 158720 220786 158732
rect 227898 158720 227904 158732
rect 227956 158720 227962 158772
rect 230842 158720 230848 158772
rect 230900 158760 230906 158772
rect 238018 158760 238024 158772
rect 230900 158732 238024 158760
rect 230900 158720 230906 158732
rect 238018 158720 238024 158732
rect 238076 158720 238082 158772
rect 248506 158720 248512 158772
rect 248564 158760 248570 158772
rect 249610 158760 249616 158772
rect 248564 158732 249616 158760
rect 248564 158720 248570 158732
rect 249610 158720 249616 158732
rect 249668 158720 249674 158772
rect 256878 158720 256884 158772
rect 256936 158760 256942 158772
rect 257982 158760 257988 158772
rect 256936 158732 257988 158760
rect 256936 158720 256942 158732
rect 257982 158720 257988 158732
rect 258040 158720 258046 158772
rect 268654 158720 268660 158772
rect 268712 158760 268718 158772
rect 271690 158760 271696 158772
rect 268712 158732 271696 158760
rect 268712 158720 268718 158732
rect 271690 158720 271696 158732
rect 271748 158720 271754 158772
rect 286318 158720 286324 158772
rect 286376 158760 286382 158772
rect 286870 158760 286876 158772
rect 286376 158732 286876 158760
rect 286376 158720 286382 158732
rect 286870 158720 286876 158732
rect 286928 158720 286934 158772
rect 288894 158720 288900 158772
rect 288952 158760 288958 158772
rect 292298 158760 292304 158772
rect 288952 158732 292304 158760
rect 288952 158720 288958 158732
rect 292298 158720 292304 158732
rect 292356 158720 292362 158772
rect 301498 158720 301504 158772
rect 301556 158760 301562 158772
rect 304810 158760 304816 158772
rect 301556 158732 304816 158760
rect 301556 158720 301562 158732
rect 304810 158720 304816 158732
rect 304868 158720 304874 158772
rect 335998 158720 336004 158772
rect 336056 158760 336062 158772
rect 337746 158760 337752 158772
rect 336056 158732 337752 158760
rect 336056 158720 336062 158732
rect 337746 158720 337752 158732
rect 337804 158720 337810 158772
rect 385586 158720 385592 158772
rect 385644 158760 385650 158772
rect 389082 158760 389088 158772
rect 385644 158732 389088 158760
rect 385644 158720 385650 158732
rect 389082 158720 389088 158732
rect 389140 158720 389146 158772
rect 430206 158720 430212 158772
rect 430264 158760 430270 158772
rect 433242 158760 433248 158772
rect 430264 158732 433248 158760
rect 430264 158720 430270 158732
rect 433242 158720 433248 158732
rect 433300 158720 433306 158772
rect 458726 158720 458732 158772
rect 458784 158760 458790 158772
rect 463326 158760 463332 158772
rect 458784 158732 463332 158760
rect 458784 158720 458790 158732
rect 463326 158720 463332 158732
rect 463384 158720 463390 158772
rect 476390 158720 476396 158772
rect 476448 158760 476454 158772
rect 482646 158760 482652 158772
rect 476448 158732 482652 158760
rect 476448 158720 476454 158732
rect 482646 158720 482652 158732
rect 482704 158720 482710 158772
rect 485682 158720 485688 158772
rect 485740 158760 485746 158772
rect 488626 158760 488632 158772
rect 485740 158732 488632 158760
rect 485740 158720 485746 158732
rect 488626 158720 488632 158732
rect 488684 158720 488690 158772
rect 490742 158720 490748 158772
rect 490800 158760 490806 158772
rect 493502 158760 493508 158772
rect 490800 158732 493508 158760
rect 490800 158720 490806 158732
rect 493502 158720 493508 158732
rect 493560 158720 493566 158772
rect 494054 158720 494060 158772
rect 494112 158760 494118 158772
rect 495710 158760 495716 158772
rect 494112 158732 495716 158760
rect 494112 158720 494118 158732
rect 495710 158720 495716 158732
rect 495768 158720 495774 158772
rect 495802 158720 495808 158772
rect 495860 158760 495866 158772
rect 496998 158760 497004 158772
rect 495860 158732 497004 158760
rect 495860 158720 495866 158732
rect 496998 158720 497004 158732
rect 497056 158720 497062 158772
rect 499666 158720 499672 158772
rect 499724 158760 499730 158772
rect 500586 158760 500592 158772
rect 499724 158732 500592 158760
rect 499724 158720 499730 158732
rect 500586 158720 500592 158732
rect 500644 158720 500650 158772
rect 504450 158720 504456 158772
rect 504508 158760 504514 158772
rect 505002 158760 505008 158772
rect 504508 158732 505008 158760
rect 504508 158720 504514 158732
rect 505002 158720 505008 158732
rect 505060 158720 505066 158772
rect 66272 158664 74534 158692
rect 74506 158624 74534 158664
rect 86126 158652 86132 158704
rect 86184 158692 86190 158704
rect 183554 158692 183560 158704
rect 86184 158664 183560 158692
rect 86184 158652 86190 158664
rect 183554 158652 183560 158664
rect 183612 158652 183618 158704
rect 195238 158652 195244 158704
rect 195296 158692 195302 158704
rect 218698 158692 218704 158704
rect 195296 158664 218704 158692
rect 195296 158652 195302 158664
rect 218698 158652 218704 158664
rect 218756 158652 218762 158704
rect 220170 158652 220176 158704
rect 220228 158692 220234 158704
rect 277946 158692 277952 158704
rect 220228 158664 277952 158692
rect 220228 158652 220234 158664
rect 277946 158652 277952 158664
rect 278004 158652 278010 158704
rect 321646 158652 321652 158704
rect 321704 158692 321710 158704
rect 359458 158692 359464 158704
rect 321704 158664 359464 158692
rect 321704 158652 321710 158664
rect 359458 158652 359464 158664
rect 359516 158652 359522 158704
rect 168374 158624 168380 158636
rect 74506 158596 168380 158624
rect 168374 158584 168380 158596
rect 168432 158584 168438 158636
rect 169754 158584 169760 158636
rect 169812 158624 169818 158636
rect 194594 158624 194600 158636
rect 169812 158596 194600 158624
rect 169812 158584 169818 158596
rect 194594 158584 194600 158596
rect 194652 158584 194658 158636
rect 200574 158584 200580 158636
rect 200632 158624 200638 158636
rect 272058 158624 272064 158636
rect 200632 158596 272064 158624
rect 200632 158584 200638 158596
rect 272058 158584 272064 158596
rect 272116 158584 272122 158636
rect 279602 158584 279608 158636
rect 279660 158624 279666 158636
rect 331306 158624 331312 158636
rect 279660 158596 331312 158624
rect 279660 158584 279666 158596
rect 331306 158584 331312 158596
rect 331364 158584 331370 158636
rect 351914 158584 351920 158636
rect 351972 158624 351978 158636
rect 386506 158624 386512 158636
rect 351972 158596 386512 158624
rect 351972 158584 351978 158596
rect 386506 158584 386512 158596
rect 386564 158584 386570 158636
rect 62574 158516 62580 158568
rect 62632 158556 62638 158568
rect 166718 158556 166724 158568
rect 62632 158528 166724 158556
rect 62632 158516 62638 158528
rect 166718 158516 166724 158528
rect 166776 158516 166782 158568
rect 190454 158516 190460 158568
rect 190512 158556 190518 158568
rect 263778 158556 263784 158568
rect 190512 158528 263784 158556
rect 190512 158516 190518 158528
rect 263778 158516 263784 158528
rect 263836 158516 263842 158568
rect 274542 158516 274548 158568
rect 274600 158556 274606 158568
rect 328546 158556 328552 158568
rect 274600 158528 328552 158556
rect 274600 158516 274606 158528
rect 328546 158516 328552 158528
rect 328604 158516 328610 158568
rect 351086 158516 351092 158568
rect 351144 158556 351150 158568
rect 386966 158556 386972 158568
rect 351144 158528 386972 158556
rect 351144 158516 351150 158528
rect 386966 158516 386972 158528
rect 387024 158516 387030 158568
rect 29822 158448 29828 158500
rect 29880 158488 29886 158500
rect 55766 158488 55772 158500
rect 29880 158460 55772 158488
rect 29880 158448 29886 158460
rect 55766 158448 55772 158460
rect 55824 158448 55830 158500
rect 59262 158448 59268 158500
rect 59320 158488 59326 158500
rect 163038 158488 163044 158500
rect 59320 158460 163044 158488
rect 59320 158448 59326 158460
rect 163038 158448 163044 158460
rect 163096 158448 163102 158500
rect 165522 158448 165528 158500
rect 165580 158488 165586 158500
rect 190546 158488 190552 158500
rect 165580 158460 190552 158488
rect 165580 158448 165586 158460
rect 190546 158448 190552 158460
rect 190604 158448 190610 158500
rect 197170 158448 197176 158500
rect 197228 158488 197234 158500
rect 269390 158488 269396 158500
rect 197228 158460 269396 158488
rect 197228 158448 197234 158460
rect 269390 158448 269396 158460
rect 269448 158448 269454 158500
rect 272886 158448 272892 158500
rect 272944 158488 272950 158500
rect 327074 158488 327080 158500
rect 272944 158460 327080 158488
rect 272944 158448 272950 158460
rect 327074 158448 327080 158460
rect 327132 158448 327138 158500
rect 338482 158448 338488 158500
rect 338540 158488 338546 158500
rect 376846 158488 376852 158500
rect 338540 158460 376852 158488
rect 338540 158448 338546 158460
rect 376846 158448 376852 158460
rect 376904 158448 376910 158500
rect 377214 158448 377220 158500
rect 377272 158488 377278 158500
rect 406838 158488 406844 158500
rect 377272 158460 406844 158488
rect 377272 158448 377278 158460
rect 406838 158448 406844 158460
rect 406896 158448 406902 158500
rect 52454 158380 52460 158432
rect 52512 158420 52518 158432
rect 52512 158392 155172 158420
rect 52512 158380 52518 158392
rect 45738 158312 45744 158364
rect 45796 158352 45802 158364
rect 153378 158352 153384 158364
rect 45796 158324 153384 158352
rect 45796 158312 45802 158324
rect 153378 158312 153384 158324
rect 153436 158312 153442 158364
rect 155144 158352 155172 158392
rect 158714 158380 158720 158432
rect 158772 158420 158778 158432
rect 185026 158420 185032 158432
rect 158772 158392 185032 158420
rect 158772 158380 158778 158392
rect 185026 158380 185032 158392
rect 185084 158380 185090 158432
rect 187050 158380 187056 158432
rect 187108 158420 187114 158432
rect 260834 158420 260840 158432
rect 187108 158392 260840 158420
rect 187108 158380 187114 158392
rect 260834 158380 260840 158392
rect 260892 158380 260898 158432
rect 266170 158380 266176 158432
rect 266228 158420 266234 158432
rect 322106 158420 322112 158432
rect 266228 158392 322112 158420
rect 266228 158380 266234 158392
rect 322106 158380 322112 158392
rect 322164 158380 322170 158432
rect 330110 158380 330116 158432
rect 330168 158420 330174 158432
rect 370866 158420 370872 158432
rect 330168 158392 370872 158420
rect 330168 158380 330174 158392
rect 370866 158380 370872 158392
rect 370924 158380 370930 158432
rect 158990 158352 158996 158364
rect 155144 158324 158996 158352
rect 158990 158312 158996 158324
rect 159048 158312 159054 158364
rect 177022 158312 177028 158364
rect 177080 158352 177086 158364
rect 254026 158352 254032 158364
rect 177080 158324 254032 158352
rect 177080 158312 177086 158324
rect 254026 158312 254032 158324
rect 254084 158312 254090 158364
rect 256050 158312 256056 158364
rect 256108 158352 256114 158364
rect 314378 158352 314384 158364
rect 256108 158324 314384 158352
rect 256108 158312 256114 158324
rect 314378 158312 314384 158324
rect 314436 158312 314442 158364
rect 320818 158312 320824 158364
rect 320876 158352 320882 158364
rect 363506 158352 363512 158364
rect 320876 158324 363512 158352
rect 320876 158312 320882 158324
rect 363506 158312 363512 158324
rect 363564 158312 363570 158364
rect 378042 158312 378048 158364
rect 378100 158352 378106 158364
rect 407390 158352 407396 158364
rect 378100 158324 407396 158352
rect 378100 158312 378106 158324
rect 407390 158312 407396 158324
rect 407448 158312 407454 158364
rect 42426 158244 42432 158296
rect 42484 158284 42490 158296
rect 150526 158284 150532 158296
rect 42484 158256 150532 158284
rect 42484 158244 42490 158256
rect 150526 158244 150532 158256
rect 150584 158244 150590 158296
rect 173618 158244 173624 158296
rect 173676 158284 173682 158296
rect 251450 158284 251456 158296
rect 173676 158256 251456 158284
rect 173676 158244 173682 158256
rect 251450 158244 251456 158256
rect 251508 158244 251514 158296
rect 252646 158244 252652 158296
rect 252704 158284 252710 158296
rect 310606 158284 310612 158296
rect 252704 158256 310612 158284
rect 252704 158244 252710 158256
rect 310606 158244 310612 158256
rect 310664 158244 310670 158296
rect 317414 158244 317420 158296
rect 317472 158284 317478 158296
rect 360194 158284 360200 158296
rect 317472 158256 360200 158284
rect 317472 158244 317478 158256
rect 360194 158244 360200 158256
rect 360252 158244 360258 158296
rect 367094 158244 367100 158296
rect 367152 158284 367158 158296
rect 399110 158284 399116 158296
rect 367152 158256 399116 158284
rect 367152 158244 367158 158256
rect 399110 158244 399116 158256
rect 399168 158244 399174 158296
rect 426434 158244 426440 158296
rect 426492 158284 426498 158296
rect 442994 158284 443000 158296
rect 426492 158256 443000 158284
rect 426492 158244 426498 158256
rect 442994 158244 443000 158256
rect 443052 158244 443058 158296
rect 31478 158176 31484 158228
rect 31536 158216 31542 158228
rect 139486 158216 139492 158228
rect 31536 158188 139492 158216
rect 31536 158176 31542 158188
rect 139486 158176 139492 158188
rect 139544 158176 139550 158228
rect 163498 158176 163504 158228
rect 163556 158216 163562 158228
rect 242894 158216 242900 158228
rect 163556 158188 242900 158216
rect 163556 158176 163562 158188
rect 242894 158176 242900 158188
rect 242952 158176 242958 158228
rect 245930 158176 245936 158228
rect 245988 158216 245994 158228
rect 306374 158216 306380 158228
rect 245988 158188 306380 158216
rect 245988 158176 245994 158188
rect 306374 158176 306380 158188
rect 306432 158176 306438 158228
rect 314102 158176 314108 158228
rect 314160 158216 314166 158228
rect 357618 158216 357624 158228
rect 314160 158188 357624 158216
rect 314160 158176 314166 158188
rect 357618 158176 357624 158188
rect 357676 158176 357682 158228
rect 361206 158176 361212 158228
rect 361264 158216 361270 158228
rect 394694 158216 394700 158228
rect 361264 158188 394700 158216
rect 361264 158176 361270 158188
rect 394694 158176 394700 158188
rect 394752 158176 394758 158228
rect 404906 158176 404912 158228
rect 404964 158216 404970 158228
rect 427998 158216 428004 158228
rect 404964 158188 428004 158216
rect 404964 158176 404970 158188
rect 427998 158176 428004 158188
rect 428056 158176 428062 158228
rect 439406 158176 439412 158228
rect 439464 158216 439470 158228
rect 454402 158216 454408 158228
rect 439464 158188 454408 158216
rect 439464 158176 439470 158188
rect 454402 158176 454408 158188
rect 454460 158176 454466 158228
rect 32306 158108 32312 158160
rect 32364 158148 32370 158160
rect 143626 158148 143632 158160
rect 32364 158120 143632 158148
rect 32364 158108 32370 158120
rect 143626 158108 143632 158120
rect 143684 158108 143690 158160
rect 153470 158108 153476 158160
rect 153528 158148 153534 158160
rect 236086 158148 236092 158160
rect 153528 158120 236092 158148
rect 153528 158108 153534 158120
rect 236086 158108 236092 158120
rect 236144 158108 236150 158160
rect 242618 158108 242624 158160
rect 242676 158148 242682 158160
rect 304074 158148 304080 158160
rect 242676 158120 304080 158148
rect 242676 158108 242682 158120
rect 304074 158108 304080 158120
rect 304132 158108 304138 158160
rect 307386 158108 307392 158160
rect 307444 158148 307450 158160
rect 353294 158148 353300 158160
rect 307444 158120 353300 158148
rect 307444 158108 307450 158120
rect 353294 158108 353300 158120
rect 353352 158108 353358 158160
rect 358630 158108 358636 158160
rect 358688 158148 358694 158160
rect 391934 158148 391940 158160
rect 358688 158120 391940 158148
rect 358688 158108 358694 158120
rect 391934 158108 391940 158120
rect 391992 158108 391998 158160
rect 404078 158108 404084 158160
rect 404136 158148 404142 158160
rect 427354 158148 427360 158160
rect 404136 158120 427360 158148
rect 404136 158108 404142 158120
rect 427354 158108 427360 158120
rect 427412 158108 427418 158160
rect 428458 158108 428464 158160
rect 428516 158148 428522 158160
rect 445754 158148 445760 158160
rect 428516 158120 445760 158148
rect 428516 158108 428522 158120
rect 445754 158108 445760 158120
rect 445812 158108 445818 158160
rect 448698 158108 448704 158160
rect 448756 158148 448762 158160
rect 461394 158148 461400 158160
rect 448756 158120 461400 158148
rect 448756 158108 448762 158120
rect 461394 158108 461400 158120
rect 461452 158108 461458 158160
rect 18874 158040 18880 158092
rect 18932 158080 18938 158092
rect 132494 158080 132500 158092
rect 18932 158052 132500 158080
rect 18932 158040 18938 158052
rect 132494 158040 132500 158052
rect 132552 158040 132558 158092
rect 139946 158040 139952 158092
rect 140004 158080 140010 158092
rect 224954 158080 224960 158092
rect 140004 158052 224960 158080
rect 140004 158040 140010 158052
rect 224954 158040 224960 158052
rect 225012 158040 225018 158092
rect 229094 158040 229100 158092
rect 229152 158080 229158 158092
rect 292758 158080 292764 158092
rect 229152 158052 292764 158080
rect 229152 158040 229158 158052
rect 292758 158040 292764 158052
rect 292816 158040 292822 158092
rect 293034 158040 293040 158092
rect 293092 158080 293098 158092
rect 342254 158080 342260 158092
rect 293092 158052 342260 158080
rect 293092 158040 293098 158052
rect 342254 158040 342260 158052
rect 342312 158040 342318 158092
rect 350258 158040 350264 158092
rect 350316 158080 350322 158092
rect 385218 158080 385224 158092
rect 350316 158052 385224 158080
rect 350316 158040 350322 158052
rect 385218 158040 385224 158052
rect 385276 158040 385282 158092
rect 393958 158040 393964 158092
rect 394016 158080 394022 158092
rect 419534 158080 419540 158092
rect 394016 158052 419540 158080
rect 394016 158040 394022 158052
rect 419534 158040 419540 158052
rect 419592 158040 419598 158092
rect 420914 158040 420920 158092
rect 420972 158080 420978 158092
rect 440326 158080 440332 158092
rect 420972 158052 440332 158080
rect 420972 158040 420978 158052
rect 440326 158040 440332 158052
rect 440384 158040 440390 158092
rect 443638 158040 443644 158092
rect 443696 158080 443702 158092
rect 456794 158080 456800 158092
rect 443696 158052 456800 158080
rect 443696 158040 443702 158052
rect 456794 158040 456800 158052
rect 456852 158040 456858 158092
rect 466362 158040 466368 158092
rect 466420 158080 466426 158092
rect 474918 158080 474924 158092
rect 466420 158052 474924 158080
rect 466420 158040 466426 158052
rect 474918 158040 474924 158052
rect 474976 158040 474982 158092
rect 2130 157972 2136 158024
rect 2188 158012 2194 158024
rect 120074 158012 120080 158024
rect 2188 157984 120080 158012
rect 2188 157972 2194 157984
rect 120074 157972 120080 157984
rect 120132 157972 120138 158024
rect 133230 157972 133236 158024
rect 133288 158012 133294 158024
rect 220630 158012 220636 158024
rect 133288 157984 220636 158012
rect 133288 157972 133294 157984
rect 220630 157972 220636 157984
rect 220688 157972 220694 158024
rect 225690 157972 225696 158024
rect 225748 158012 225754 158024
rect 288434 158012 288440 158024
rect 225748 157984 288440 158012
rect 225748 157972 225754 157984
rect 288434 157972 288440 157984
rect 288492 157972 288498 158024
rect 289722 157972 289728 158024
rect 289780 158012 289786 158024
rect 340046 158012 340052 158024
rect 289780 157984 340052 158012
rect 289780 157972 289786 157984
rect 340046 157972 340052 157984
rect 340104 157972 340110 158024
rect 340138 157972 340144 158024
rect 340196 158012 340202 158024
rect 378594 158012 378600 158024
rect 340196 157984 378600 158012
rect 340196 157972 340202 157984
rect 378594 157972 378600 157984
rect 378652 157972 378658 158024
rect 388070 157972 388076 158024
rect 388128 158012 388134 158024
rect 414566 158012 414572 158024
rect 388128 157984 414572 158012
rect 388128 157972 388134 157984
rect 414566 157972 414572 157984
rect 414624 157972 414630 158024
rect 415026 157972 415032 158024
rect 415084 158012 415090 158024
rect 434714 158012 434720 158024
rect 415084 157984 434720 158012
rect 415084 157972 415090 157984
rect 434714 157972 434720 157984
rect 434772 157972 434778 158024
rect 435174 157972 435180 158024
rect 435232 158012 435238 158024
rect 451090 158012 451096 158024
rect 435232 157984 451096 158012
rect 435232 157972 435238 157984
rect 451090 157972 451096 157984
rect 451148 157972 451154 158024
rect 457898 157972 457904 158024
rect 457956 158012 457962 158024
rect 468478 158012 468484 158024
rect 457956 157984 468484 158012
rect 457956 157972 457962 157984
rect 468478 157972 468484 157984
rect 468536 157972 468542 158024
rect 99558 157904 99564 157956
rect 99616 157944 99622 157956
rect 194962 157944 194968 157956
rect 99616 157916 194968 157944
rect 99616 157904 99622 157916
rect 194962 157904 194968 157916
rect 195020 157904 195026 157956
rect 207106 157904 207112 157956
rect 207164 157944 207170 157956
rect 233234 157944 233240 157956
rect 207164 157916 233240 157944
rect 207164 157904 207170 157916
rect 233234 157904 233240 157916
rect 233292 157904 233298 157956
rect 239214 157904 239220 157956
rect 239272 157944 239278 157956
rect 256694 157944 256700 157956
rect 239272 157916 256700 157944
rect 239272 157904 239278 157916
rect 256694 157904 256700 157916
rect 256752 157904 256758 157956
rect 262766 157904 262772 157956
rect 262824 157944 262830 157956
rect 319530 157944 319536 157956
rect 262824 157916 319536 157944
rect 262824 157904 262830 157916
rect 319530 157904 319536 157916
rect 319588 157904 319594 157956
rect 324314 157904 324320 157956
rect 324372 157944 324378 157956
rect 350534 157944 350540 157956
rect 324372 157916 350540 157944
rect 324372 157904 324378 157916
rect 350534 157904 350540 157916
rect 350592 157904 350598 157956
rect 106366 157836 106372 157888
rect 106424 157876 106430 157888
rect 200114 157876 200120 157888
rect 106424 157848 200120 157876
rect 106424 157836 106430 157848
rect 200114 157836 200120 157848
rect 200172 157836 200178 157888
rect 221550 157836 221556 157888
rect 221608 157876 221614 157888
rect 245654 157876 245660 157888
rect 221608 157848 245660 157876
rect 221608 157836 221614 157848
rect 245654 157836 245660 157848
rect 245712 157836 245718 157888
rect 259454 157836 259460 157888
rect 259512 157876 259518 157888
rect 316954 157876 316960 157888
rect 259512 157848 316960 157876
rect 259512 157836 259518 157848
rect 316954 157836 316960 157848
rect 317012 157836 317018 157888
rect 123110 157768 123116 157820
rect 123168 157808 123174 157820
rect 207106 157808 207112 157820
rect 123168 157780 207112 157808
rect 123168 157768 123174 157780
rect 207106 157768 207112 157780
rect 207164 157768 207170 157820
rect 269482 157768 269488 157820
rect 269540 157808 269546 157820
rect 324682 157808 324688 157820
rect 269540 157780 324688 157808
rect 269540 157768 269546 157780
rect 324682 157768 324688 157780
rect 324740 157768 324746 157820
rect 144822 157700 144828 157752
rect 144880 157740 144886 157752
rect 169938 157740 169944 157752
rect 144880 157712 169944 157740
rect 144880 157700 144886 157712
rect 169938 157700 169944 157712
rect 169996 157700 170002 157752
rect 201310 157700 201316 157752
rect 201368 157740 201374 157752
rect 223850 157740 223856 157752
rect 201368 157712 223856 157740
rect 201368 157700 201374 157712
rect 223850 157700 223856 157712
rect 223908 157700 223914 157752
rect 311894 157700 311900 157752
rect 311952 157740 311958 157752
rect 341334 157740 341340 157752
rect 311952 157712 341340 157740
rect 311952 157700 311958 157712
rect 341334 157700 341340 157712
rect 341392 157700 341398 157752
rect 79962 157292 79968 157344
rect 80020 157332 80026 157344
rect 177022 157332 177028 157344
rect 80020 157304 177028 157332
rect 80020 157292 80026 157304
rect 177022 157292 177028 157304
rect 177080 157292 177086 157344
rect 193766 157292 193772 157344
rect 193824 157332 193830 157344
rect 266906 157332 266912 157344
rect 193824 157304 266912 157332
rect 193824 157292 193830 157304
rect 266906 157292 266912 157304
rect 266964 157292 266970 157344
rect 296438 157292 296444 157344
rect 296496 157332 296502 157344
rect 345014 157332 345020 157344
rect 296496 157304 345020 157332
rect 296496 157292 296502 157304
rect 345014 157292 345020 157304
rect 345072 157292 345078 157344
rect 356146 157292 356152 157344
rect 356204 157332 356210 157344
rect 358906 157332 358912 157344
rect 356204 157304 358912 157332
rect 356204 157292 356210 157304
rect 358906 157292 358912 157304
rect 358964 157292 358970 157344
rect 69290 157224 69296 157276
rect 69348 157264 69354 157276
rect 171134 157264 171140 157276
rect 69348 157236 171140 157264
rect 69348 157224 69354 157236
rect 171134 157224 171140 157236
rect 171192 157224 171198 157276
rect 179506 157224 179512 157276
rect 179564 157264 179570 157276
rect 255866 157264 255872 157276
rect 179564 157236 255872 157264
rect 179564 157224 179570 157236
rect 255866 157224 255872 157236
rect 255924 157224 255930 157276
rect 276198 157224 276204 157276
rect 276256 157264 276262 157276
rect 329834 157264 329840 157276
rect 276256 157236 329840 157264
rect 276256 157224 276262 157236
rect 329834 157224 329840 157236
rect 329892 157224 329898 157276
rect 352006 157224 352012 157276
rect 352064 157264 352070 157276
rect 365898 157264 365904 157276
rect 352064 157236 365904 157264
rect 352064 157224 352070 157236
rect 365898 157224 365904 157236
rect 365956 157224 365962 157276
rect 4522 157156 4528 157208
rect 4580 157196 4586 157208
rect 109126 157196 109132 157208
rect 4580 157168 109132 157196
rect 4580 157156 4586 157168
rect 109126 157156 109132 157168
rect 109184 157156 109190 157208
rect 113082 157156 113088 157208
rect 113140 157196 113146 157208
rect 205266 157196 205272 157208
rect 113140 157168 205272 157196
rect 113140 157156 113146 157168
rect 205266 157156 205272 157168
rect 205324 157156 205330 157208
rect 209774 157156 209780 157208
rect 209832 157196 209838 157208
rect 278774 157196 278780 157208
rect 209832 157168 278780 157196
rect 209832 157156 209838 157168
rect 278774 157156 278780 157168
rect 278832 157156 278838 157208
rect 288618 157156 288624 157208
rect 288676 157196 288682 157208
rect 338666 157196 338672 157208
rect 288676 157168 338672 157196
rect 288676 157156 288682 157168
rect 338666 157156 338672 157168
rect 338724 157156 338730 157208
rect 347774 157156 347780 157208
rect 347832 157196 347838 157208
rect 383654 157196 383660 157208
rect 347832 157168 383660 157196
rect 347832 157156 347838 157168
rect 383654 157156 383660 157168
rect 383712 157156 383718 157208
rect 55858 157088 55864 157140
rect 55916 157128 55922 157140
rect 161566 157128 161572 157140
rect 55916 157100 161572 157128
rect 55916 157088 55922 157100
rect 161566 157088 161572 157100
rect 161624 157088 161630 157140
rect 172790 157088 172796 157140
rect 172848 157128 172854 157140
rect 250806 157128 250812 157140
rect 172848 157100 250812 157128
rect 172848 157088 172854 157100
rect 250806 157088 250812 157100
rect 250864 157088 250870 157140
rect 260282 157088 260288 157140
rect 260340 157128 260346 157140
rect 317414 157128 317420 157140
rect 260340 157100 317420 157128
rect 260340 157088 260346 157100
rect 317414 157088 317420 157100
rect 317472 157088 317478 157140
rect 346854 157088 346860 157140
rect 346912 157128 346918 157140
rect 383746 157128 383752 157140
rect 346912 157100 383752 157128
rect 346912 157088 346918 157100
rect 383746 157088 383752 157100
rect 383804 157088 383810 157140
rect 49142 157020 49148 157072
rect 49200 157060 49206 157072
rect 156414 157060 156420 157072
rect 49200 157032 156420 157060
rect 49200 157020 49206 157032
rect 156414 157020 156420 157032
rect 156472 157020 156478 157072
rect 176102 157020 176108 157072
rect 176160 157060 176166 157072
rect 252554 157060 252560 157072
rect 176160 157032 252560 157060
rect 176160 157020 176166 157032
rect 252554 157020 252560 157032
rect 252612 157020 252618 157072
rect 254394 157020 254400 157072
rect 254452 157060 254458 157072
rect 311894 157060 311900 157072
rect 254452 157032 311900 157060
rect 254452 157020 254458 157032
rect 311894 157020 311900 157032
rect 311952 157020 311958 157072
rect 336826 157020 336832 157072
rect 336884 157060 336890 157072
rect 376018 157060 376024 157072
rect 336884 157032 376024 157060
rect 336884 157020 336890 157032
rect 376018 157020 376024 157032
rect 376076 157020 376082 157072
rect 383102 157020 383108 157072
rect 383160 157060 383166 157072
rect 411346 157060 411352 157072
rect 383160 157032 411352 157060
rect 383160 157020 383166 157032
rect 411346 157020 411352 157032
rect 411404 157020 411410 157072
rect 39022 156952 39028 157004
rect 39080 156992 39086 157004
rect 147674 156992 147680 157004
rect 39080 156964 147680 156992
rect 39080 156952 39086 156964
rect 147674 156952 147680 156964
rect 147732 156952 147738 157004
rect 169386 156952 169392 157004
rect 169444 156992 169450 157004
rect 247126 156992 247132 157004
rect 169444 156964 247132 156992
rect 169444 156952 169450 156964
rect 247126 156952 247132 156964
rect 247184 156952 247190 157004
rect 253566 156952 253572 157004
rect 253624 156992 253630 157004
rect 307018 156992 307024 157004
rect 253624 156964 307024 156992
rect 253624 156952 253630 156964
rect 307018 156952 307024 156964
rect 307076 156952 307082 157004
rect 330938 156952 330944 157004
rect 330996 156992 331002 157004
rect 371234 156992 371240 157004
rect 330996 156964 371240 156992
rect 330996 156952 331002 156964
rect 371234 156952 371240 156964
rect 371292 156952 371298 157004
rect 374638 156952 374644 157004
rect 374696 156992 374702 157004
rect 404446 156992 404452 157004
rect 374696 156964 404452 156992
rect 374696 156952 374702 156964
rect 404446 156952 404452 156964
rect 404504 156952 404510 157004
rect 423398 156952 423404 157004
rect 423456 156992 423462 157004
rect 442166 156992 442172 157004
rect 423456 156964 442172 156992
rect 423456 156952 423462 156964
rect 442166 156952 442172 156964
rect 442224 156952 442230 157004
rect 464890 156952 464896 157004
rect 464948 156992 464954 157004
rect 471054 156992 471060 157004
rect 464948 156964 471060 156992
rect 464948 156952 464954 156964
rect 471054 156952 471060 156964
rect 471112 156952 471118 157004
rect 28074 156884 28080 156936
rect 28132 156924 28138 156936
rect 139394 156924 139400 156936
rect 28132 156896 139400 156924
rect 28132 156884 28138 156896
rect 139394 156884 139400 156896
rect 139452 156884 139458 156936
rect 160186 156884 160192 156936
rect 160244 156924 160250 156936
rect 240134 156924 240140 156936
rect 160244 156896 240140 156924
rect 160244 156884 160250 156896
rect 240134 156884 240140 156896
rect 240192 156884 240198 156936
rect 249334 156884 249340 156936
rect 249392 156924 249398 156936
rect 306374 156924 306380 156936
rect 249392 156896 306380 156924
rect 249392 156884 249398 156896
rect 306374 156884 306380 156896
rect 306432 156884 306438 156936
rect 307294 156924 307300 156936
rect 306484 156896 307300 156924
rect 24762 156816 24768 156868
rect 24820 156856 24826 156868
rect 137830 156856 137836 156868
rect 24820 156828 137836 156856
rect 24820 156816 24826 156828
rect 137830 156816 137836 156828
rect 137888 156816 137894 156868
rect 150066 156816 150072 156868
rect 150124 156856 150130 156868
rect 233510 156856 233516 156868
rect 150124 156828 233516 156856
rect 150124 156816 150130 156828
rect 233510 156816 233516 156828
rect 233568 156816 233574 156868
rect 246758 156816 246764 156868
rect 246816 156856 246822 156868
rect 306484 156856 306512 156896
rect 307294 156884 307300 156896
rect 307352 156884 307358 156936
rect 310698 156884 310704 156936
rect 310756 156924 310762 156936
rect 356146 156924 356152 156936
rect 310756 156896 356152 156924
rect 310756 156884 310762 156896
rect 356146 156884 356152 156896
rect 356204 156884 356210 156936
rect 373810 156884 373816 156936
rect 373868 156924 373874 156936
rect 404078 156924 404084 156936
rect 373868 156896 404084 156924
rect 373868 156884 373874 156896
rect 404078 156884 404084 156896
rect 404136 156884 404142 156936
rect 411622 156884 411628 156936
rect 411680 156924 411686 156936
rect 433150 156924 433156 156936
rect 411680 156896 433156 156924
rect 411680 156884 411686 156896
rect 433150 156884 433156 156896
rect 433208 156884 433214 156936
rect 436554 156884 436560 156936
rect 436612 156924 436618 156936
rect 448606 156924 448612 156936
rect 436612 156896 448612 156924
rect 436612 156884 436618 156896
rect 448606 156884 448612 156896
rect 448664 156884 448670 156936
rect 246816 156828 306512 156856
rect 246816 156816 246822 156828
rect 306650 156816 306656 156868
rect 306708 156856 306714 156868
rect 351914 156856 351920 156868
rect 306708 156828 351920 156856
rect 306708 156816 306714 156828
rect 351914 156816 351920 156828
rect 351972 156816 351978 156868
rect 363690 156816 363696 156868
rect 363748 156856 363754 156868
rect 396534 156856 396540 156868
rect 363748 156828 396540 156856
rect 363748 156816 363754 156828
rect 396534 156816 396540 156828
rect 396592 156816 396598 156868
rect 400766 156816 400772 156868
rect 400824 156856 400830 156868
rect 423766 156856 423772 156868
rect 400824 156828 423772 156856
rect 400824 156816 400830 156828
rect 423766 156816 423772 156828
rect 423824 156816 423830 156868
rect 433242 156816 433248 156868
rect 433300 156856 433306 156868
rect 447318 156856 447324 156868
rect 433300 156828 447324 156856
rect 433300 156816 433306 156828
rect 447318 156816 447324 156828
rect 447376 156816 447382 156868
rect 18046 156748 18052 156800
rect 18104 156788 18110 156800
rect 132678 156788 132684 156800
rect 18104 156760 132684 156788
rect 18104 156748 18110 156760
rect 132678 156748 132684 156760
rect 132736 156748 132742 156800
rect 136634 156748 136640 156800
rect 136692 156788 136698 156800
rect 222746 156788 222752 156800
rect 136692 156760 222752 156788
rect 136692 156748 136698 156760
rect 222746 156748 222752 156760
rect 222804 156748 222810 156800
rect 240042 156748 240048 156800
rect 240100 156788 240106 156800
rect 302234 156788 302240 156800
rect 240100 156760 302240 156788
rect 240100 156748 240106 156760
rect 302234 156748 302240 156760
rect 302292 156748 302298 156800
rect 303154 156748 303160 156800
rect 303212 156788 303218 156800
rect 349246 156788 349252 156800
rect 303212 156760 349252 156788
rect 303212 156748 303218 156760
rect 349246 156748 349252 156760
rect 349304 156748 349310 156800
rect 357802 156748 357808 156800
rect 357860 156788 357866 156800
rect 392118 156788 392124 156800
rect 357860 156760 392124 156788
rect 357860 156748 357866 156760
rect 392118 156748 392124 156760
rect 392176 156748 392182 156800
rect 401594 156748 401600 156800
rect 401652 156788 401658 156800
rect 425146 156788 425152 156800
rect 401652 156760 425152 156788
rect 401652 156748 401658 156760
rect 425146 156748 425152 156760
rect 425204 156748 425210 156800
rect 427630 156748 427636 156800
rect 427688 156788 427694 156800
rect 444374 156788 444380 156800
rect 427688 156760 444380 156788
rect 427688 156748 427694 156760
rect 444374 156748 444380 156760
rect 444432 156748 444438 156800
rect 11238 156680 11244 156732
rect 11296 156720 11302 156732
rect 125686 156720 125692 156732
rect 11296 156692 125692 156720
rect 11296 156680 11302 156692
rect 125686 156680 125692 156692
rect 125744 156680 125750 156732
rect 126514 156680 126520 156732
rect 126572 156720 126578 156732
rect 215478 156720 215484 156732
rect 126572 156692 215484 156720
rect 126572 156680 126578 156692
rect 215478 156680 215484 156692
rect 215536 156680 215542 156732
rect 216674 156680 216680 156732
rect 216732 156720 216738 156732
rect 282086 156720 282092 156732
rect 216732 156692 282092 156720
rect 216732 156680 216738 156692
rect 282086 156680 282092 156692
rect 282144 156680 282150 156732
rect 283006 156680 283012 156732
rect 283064 156720 283070 156732
rect 334894 156720 334900 156732
rect 283064 156692 334900 156720
rect 283064 156680 283070 156692
rect 334894 156680 334900 156692
rect 334952 156680 334958 156732
rect 341886 156680 341892 156732
rect 341944 156720 341950 156732
rect 379882 156720 379888 156732
rect 341944 156692 379888 156720
rect 341944 156680 341950 156692
rect 379882 156680 379888 156692
rect 379940 156680 379946 156732
rect 384758 156680 384764 156732
rect 384816 156720 384822 156732
rect 412634 156720 412640 156732
rect 384816 156692 412640 156720
rect 384816 156680 384822 156692
rect 412634 156680 412640 156692
rect 412692 156680 412698 156732
rect 419258 156680 419264 156732
rect 419316 156720 419322 156732
rect 438946 156720 438952 156732
rect 419316 156692 438952 156720
rect 419316 156680 419322 156692
rect 438946 156680 438952 156692
rect 439004 156680 439010 156732
rect 446122 156680 446128 156732
rect 446180 156720 446186 156732
rect 459462 156720 459468 156732
rect 446180 156692 459468 156720
rect 446180 156680 446186 156692
rect 459462 156680 459468 156692
rect 459520 156680 459526 156732
rect 14642 156612 14648 156664
rect 14700 156652 14706 156664
rect 129734 156652 129740 156664
rect 14700 156624 129740 156652
rect 14700 156612 14706 156624
rect 129734 156612 129740 156624
rect 129792 156612 129798 156664
rect 129918 156612 129924 156664
rect 129976 156652 129982 156664
rect 218054 156652 218060 156664
rect 129976 156624 218060 156652
rect 129976 156612 129982 156624
rect 218054 156612 218060 156624
rect 218112 156612 218118 156664
rect 236730 156612 236736 156664
rect 236788 156652 236794 156664
rect 299658 156652 299664 156664
rect 236788 156624 299664 156652
rect 236788 156612 236794 156624
rect 299658 156612 299664 156624
rect 299716 156612 299722 156664
rect 299750 156612 299756 156664
rect 299808 156652 299814 156664
rect 347774 156652 347780 156664
rect 299808 156624 347780 156652
rect 299808 156612 299814 156624
rect 347774 156612 347780 156624
rect 347832 156612 347838 156664
rect 348602 156612 348608 156664
rect 348660 156652 348666 156664
rect 385034 156652 385040 156664
rect 348660 156624 385040 156652
rect 348660 156612 348666 156624
rect 385034 156612 385040 156624
rect 385092 156612 385098 156664
rect 387242 156612 387248 156664
rect 387300 156652 387306 156664
rect 414106 156652 414112 156664
rect 387300 156624 414112 156652
rect 387300 156612 387306 156624
rect 414106 156612 414112 156624
rect 414164 156612 414170 156664
rect 414198 156612 414204 156664
rect 414256 156652 414262 156664
rect 435082 156652 435088 156664
rect 414256 156624 435088 156652
rect 414256 156612 414262 156624
rect 435082 156612 435088 156624
rect 435140 156612 435146 156664
rect 445294 156612 445300 156664
rect 445352 156652 445358 156664
rect 445352 156624 451274 156652
rect 445352 156612 445358 156624
rect 96246 156544 96252 156596
rect 96304 156584 96310 156596
rect 192386 156584 192392 156596
rect 96304 156556 192392 156584
rect 96304 156544 96310 156556
rect 192386 156544 192392 156556
rect 192444 156544 192450 156596
rect 215018 156544 215024 156596
rect 215076 156584 215082 156596
rect 279326 156584 279332 156596
rect 215076 156556 279332 156584
rect 215076 156544 215082 156556
rect 279326 156544 279332 156556
rect 279384 156544 279390 156596
rect 303982 156544 303988 156596
rect 304040 156584 304046 156596
rect 350994 156584 351000 156596
rect 304040 156556 351000 156584
rect 304040 156544 304046 156556
rect 350994 156544 351000 156556
rect 351052 156544 351058 156596
rect 451246 156584 451274 156624
rect 458174 156612 458180 156664
rect 458232 156652 458238 156664
rect 465258 156652 465264 156664
rect 458232 156624 465264 156652
rect 458232 156612 458238 156624
rect 465258 156612 465264 156624
rect 465316 156612 465322 156664
rect 458358 156584 458364 156596
rect 451246 156556 458364 156584
rect 458358 156544 458364 156556
rect 458416 156544 458422 156596
rect 109678 156476 109684 156528
rect 109736 156516 109742 156528
rect 194318 156516 194324 156528
rect 109736 156488 194324 156516
rect 109736 156476 109742 156488
rect 194318 156476 194324 156488
rect 194376 156476 194382 156528
rect 227714 156476 227720 156528
rect 227772 156516 227778 156528
rect 289998 156516 290004 156528
rect 227772 156488 290004 156516
rect 227772 156476 227778 156488
rect 289998 156476 290004 156488
rect 290056 156476 290062 156528
rect 307018 156476 307024 156528
rect 307076 156516 307082 156528
rect 312446 156516 312452 156528
rect 307076 156488 312452 156516
rect 307076 156476 307082 156488
rect 312446 156476 312452 156488
rect 312504 156476 312510 156528
rect 317782 156476 317788 156528
rect 317840 156516 317846 156528
rect 354214 156516 354220 156528
rect 317840 156488 354220 156516
rect 317840 156476 317846 156488
rect 354214 156476 354220 156488
rect 354272 156476 354278 156528
rect 133414 156408 133420 156460
rect 133472 156448 133478 156460
rect 164418 156448 164424 156460
rect 133472 156420 164424 156448
rect 133472 156408 133478 156420
rect 164418 156408 164424 156420
rect 164476 156408 164482 156460
rect 176654 156408 176660 156460
rect 176712 156448 176718 156460
rect 248874 156448 248880 156460
rect 176712 156420 248880 156448
rect 176712 156408 176718 156420
rect 248874 156408 248880 156420
rect 248932 156408 248938 156460
rect 251726 156408 251732 156460
rect 251784 156448 251790 156460
rect 299474 156448 299480 156460
rect 251784 156420 299480 156448
rect 251784 156408 251790 156420
rect 299474 156408 299480 156420
rect 299532 156408 299538 156460
rect 306374 156408 306380 156460
rect 306432 156448 306438 156460
rect 309226 156448 309232 156460
rect 306432 156420 309232 156448
rect 306432 156408 306438 156420
rect 309226 156408 309232 156420
rect 309284 156408 309290 156460
rect 311986 156408 311992 156460
rect 312044 156448 312050 156460
rect 346486 156448 346492 156460
rect 312044 156420 346492 156448
rect 312044 156408 312050 156420
rect 346486 156408 346492 156420
rect 346544 156408 346550 156460
rect 140866 156340 140872 156392
rect 140924 156380 140930 156392
rect 172514 156380 172520 156392
rect 140924 156352 172520 156380
rect 140924 156340 140930 156352
rect 172514 156340 172520 156352
rect 172572 156340 172578 156392
rect 279510 156340 279516 156392
rect 279568 156380 279574 156392
rect 323394 156380 323400 156392
rect 279568 156352 323400 156380
rect 279568 156340 279574 156352
rect 323394 156340 323400 156352
rect 323452 156340 323458 156392
rect 89530 155864 89536 155916
rect 89588 155904 89594 155916
rect 187234 155904 187240 155916
rect 89588 155876 187240 155904
rect 89588 155864 89594 155876
rect 187234 155864 187240 155876
rect 187292 155864 187298 155916
rect 203886 155864 203892 155916
rect 203944 155904 203950 155916
rect 273438 155904 273444 155916
rect 203944 155876 273444 155904
rect 203944 155864 203950 155876
rect 273438 155864 273444 155876
rect 273496 155864 273502 155916
rect 324222 155864 324228 155916
rect 324280 155904 324286 155916
rect 366266 155904 366272 155916
rect 324280 155876 366272 155904
rect 324280 155864 324286 155876
rect 366266 155864 366272 155876
rect 366324 155864 366330 155916
rect 85298 155796 85304 155848
rect 85356 155836 85362 155848
rect 184014 155836 184020 155848
rect 85356 155808 184020 155836
rect 85356 155796 85362 155808
rect 184014 155796 184020 155808
rect 184072 155796 184078 155848
rect 206462 155796 206468 155848
rect 206520 155836 206526 155848
rect 276474 155836 276480 155848
rect 206520 155808 276480 155836
rect 206520 155796 206526 155808
rect 276474 155796 276480 155808
rect 276532 155796 276538 155848
rect 287146 155796 287152 155848
rect 287204 155836 287210 155848
rect 296622 155836 296628 155848
rect 287204 155808 296628 155836
rect 287204 155796 287210 155808
rect 296622 155796 296628 155808
rect 296680 155796 296686 155848
rect 297266 155796 297272 155848
rect 297324 155836 297330 155848
rect 345842 155836 345848 155848
rect 297324 155808 345848 155836
rect 297324 155796 297330 155808
rect 345842 155796 345848 155808
rect 345900 155796 345906 155848
rect 345934 155796 345940 155848
rect 345992 155836 345998 155848
rect 352282 155836 352288 155848
rect 345992 155808 352288 155836
rect 345992 155796 345998 155808
rect 352282 155796 352288 155808
rect 352340 155796 352346 155848
rect 72694 155728 72700 155780
rect 72752 155768 72758 155780
rect 174446 155768 174452 155780
rect 72752 155740 174452 155768
rect 72752 155728 72758 155740
rect 174446 155728 174452 155740
rect 174504 155728 174510 155780
rect 199654 155728 199660 155780
rect 199712 155768 199718 155780
rect 271046 155768 271052 155780
rect 199712 155740 271052 155768
rect 199712 155728 199718 155740
rect 271046 155728 271052 155740
rect 271104 155728 271110 155780
rect 280430 155728 280436 155780
rect 280488 155768 280494 155780
rect 333054 155768 333060 155780
rect 280488 155740 333060 155768
rect 280488 155728 280494 155740
rect 333054 155728 333060 155740
rect 333112 155728 333118 155780
rect 336642 155728 336648 155780
rect 336700 155768 336706 155780
rect 361942 155768 361948 155780
rect 336700 155740 361948 155768
rect 336700 155728 336706 155740
rect 361942 155728 361948 155740
rect 362000 155728 362006 155780
rect 362126 155728 362132 155780
rect 362184 155768 362190 155780
rect 367646 155768 367652 155780
rect 362184 155740 367652 155768
rect 362184 155728 362190 155740
rect 367646 155728 367652 155740
rect 367704 155728 367710 155780
rect 370406 155728 370412 155780
rect 370464 155768 370470 155780
rect 401686 155768 401692 155780
rect 370464 155740 401692 155768
rect 370464 155728 370470 155740
rect 401686 155728 401692 155740
rect 401744 155728 401750 155780
rect 55030 155660 55036 155712
rect 55088 155700 55094 155712
rect 157334 155700 157340 155712
rect 55088 155672 157340 155700
rect 55088 155660 55094 155672
rect 157334 155660 157340 155672
rect 157392 155660 157398 155712
rect 192938 155660 192944 155712
rect 192996 155700 193002 155712
rect 265158 155700 265164 155712
rect 192996 155672 265164 155700
rect 192996 155660 193002 155672
rect 265158 155660 265164 155672
rect 265216 155660 265222 155712
rect 273714 155660 273720 155712
rect 273772 155700 273778 155712
rect 327902 155700 327908 155712
rect 273772 155672 327908 155700
rect 273772 155660 273778 155672
rect 327902 155660 327908 155672
rect 327960 155660 327966 155712
rect 328362 155660 328368 155712
rect 328420 155700 328426 155712
rect 368934 155700 368940 155712
rect 328420 155672 368940 155700
rect 328420 155660 328426 155672
rect 368934 155660 368940 155672
rect 368992 155660 368998 155712
rect 369578 155660 369584 155712
rect 369636 155700 369642 155712
rect 400214 155700 400220 155712
rect 369636 155672 400220 155700
rect 369636 155660 369642 155672
rect 400214 155660 400220 155672
rect 400272 155660 400278 155712
rect 48314 155592 48320 155644
rect 48372 155632 48378 155644
rect 154666 155632 154672 155644
rect 48372 155604 154672 155632
rect 48372 155592 48378 155604
rect 154666 155592 154672 155604
rect 154724 155592 154730 155644
rect 186222 155592 186228 155644
rect 186280 155632 186286 155644
rect 261110 155632 261116 155644
rect 186280 155604 261116 155632
rect 186280 155592 186286 155604
rect 261110 155592 261116 155604
rect 261168 155592 261174 155644
rect 277118 155592 277124 155644
rect 277176 155632 277182 155644
rect 330478 155632 330484 155644
rect 277176 155604 330484 155632
rect 277176 155592 277182 155604
rect 330478 155592 330484 155604
rect 330536 155592 330542 155644
rect 334250 155592 334256 155644
rect 334308 155632 334314 155644
rect 374086 155632 374092 155644
rect 334308 155604 374092 155632
rect 334308 155592 334314 155604
rect 374086 155592 374092 155604
rect 374144 155592 374150 155644
rect 378318 155592 378324 155644
rect 378376 155632 378382 155644
rect 383102 155632 383108 155644
rect 378376 155604 383108 155632
rect 378376 155592 378382 155604
rect 383102 155592 383108 155604
rect 383160 155592 383166 155644
rect 41598 155524 41604 155576
rect 41656 155564 41662 155576
rect 150618 155564 150624 155576
rect 41656 155536 150624 155564
rect 41656 155524 41662 155536
rect 150618 155524 150624 155536
rect 150676 155524 150682 155576
rect 156782 155524 156788 155576
rect 156840 155564 156846 155576
rect 237926 155564 237932 155576
rect 156840 155536 237932 155564
rect 156840 155524 156846 155536
rect 237926 155524 237932 155536
rect 237984 155524 237990 155576
rect 238018 155524 238024 155576
rect 238076 155564 238082 155576
rect 238076 155536 291424 155564
rect 238076 155524 238082 155536
rect 23934 155456 23940 155508
rect 23992 155496 23998 155508
rect 136726 155496 136732 155508
rect 23992 155468 136732 155496
rect 23992 155456 23998 155468
rect 136726 155456 136732 155468
rect 136784 155456 136790 155508
rect 138290 155456 138296 155508
rect 138348 155496 138354 155508
rect 221734 155496 221740 155508
rect 138348 155468 221740 155496
rect 138348 155456 138354 155468
rect 221734 155456 221740 155468
rect 221792 155456 221798 155508
rect 225782 155456 225788 155508
rect 225840 155496 225846 155508
rect 291286 155496 291292 155508
rect 225840 155468 291292 155496
rect 225840 155456 225846 155468
rect 291286 155456 291292 155468
rect 291344 155456 291350 155508
rect 22186 155388 22192 155440
rect 22244 155428 22250 155440
rect 135898 155428 135904 155440
rect 22244 155400 135904 155428
rect 22244 155388 22250 155400
rect 135898 155388 135904 155400
rect 135956 155388 135962 155440
rect 146662 155388 146668 155440
rect 146720 155428 146726 155440
rect 230934 155428 230940 155440
rect 146720 155400 230940 155428
rect 146720 155388 146726 155400
rect 230934 155388 230940 155400
rect 230992 155388 230998 155440
rect 232498 155388 232504 155440
rect 232556 155428 232562 155440
rect 291396 155428 291424 155536
rect 294782 155524 294788 155576
rect 294840 155564 294846 155576
rect 343910 155564 343916 155576
rect 294840 155536 343916 155564
rect 294840 155524 294846 155536
rect 343910 155524 343916 155536
rect 343968 155524 343974 155576
rect 364518 155524 364524 155576
rect 364576 155564 364582 155576
rect 396166 155564 396172 155576
rect 364576 155536 396172 155564
rect 364576 155524 364582 155536
rect 396166 155524 396172 155536
rect 396224 155524 396230 155576
rect 293862 155456 293868 155508
rect 293920 155496 293926 155508
rect 343266 155496 343272 155508
rect 293920 155468 343272 155496
rect 293920 155456 293926 155468
rect 343266 155456 343272 155468
rect 343324 155456 343330 155508
rect 353662 155456 353668 155508
rect 353720 155496 353726 155508
rect 388346 155496 388352 155508
rect 353720 155468 388352 155496
rect 353720 155456 353726 155468
rect 388346 155456 388352 155468
rect 388404 155456 388410 155508
rect 408310 155456 408316 155508
rect 408368 155496 408374 155508
rect 430574 155496 430580 155508
rect 408368 155468 430580 155496
rect 408368 155456 408374 155468
rect 430574 155456 430580 155468
rect 430632 155456 430638 155508
rect 433058 155456 433064 155508
rect 433116 155496 433122 155508
rect 444742 155496 444748 155508
rect 433116 155468 444748 155496
rect 433116 155456 433122 155468
rect 444742 155456 444748 155468
rect 444800 155456 444806 155508
rect 295150 155428 295156 155440
rect 232556 155400 291332 155428
rect 291396 155400 295156 155428
rect 232556 155388 232562 155400
rect 15470 155320 15476 155372
rect 15528 155360 15534 155372
rect 130286 155360 130292 155372
rect 15528 155332 130292 155360
rect 15528 155320 15534 155332
rect 130286 155320 130292 155332
rect 130344 155320 130350 155372
rect 135806 155320 135812 155372
rect 135864 155360 135870 155372
rect 219526 155360 219532 155372
rect 135864 155332 219532 155360
rect 135864 155320 135870 155332
rect 219526 155320 219532 155332
rect 219584 155320 219590 155372
rect 223206 155320 223212 155372
rect 223264 155360 223270 155372
rect 289354 155360 289360 155372
rect 223264 155332 289360 155360
rect 223264 155320 223270 155332
rect 289354 155320 289360 155332
rect 289412 155320 289418 155372
rect 291304 155360 291332 155400
rect 295150 155388 295156 155400
rect 295208 155388 295214 155440
rect 300670 155388 300676 155440
rect 300728 155428 300734 155440
rect 348418 155428 348424 155440
rect 300728 155400 348424 155428
rect 300728 155388 300734 155400
rect 348418 155388 348424 155400
rect 348476 155388 348482 155440
rect 354490 155388 354496 155440
rect 354548 155428 354554 155440
rect 389542 155428 389548 155440
rect 354548 155400 389548 155428
rect 354548 155388 354554 155400
rect 389542 155388 389548 155400
rect 389600 155388 389606 155440
rect 394878 155388 394884 155440
rect 394936 155428 394942 155440
rect 420362 155428 420368 155440
rect 394936 155400 420368 155428
rect 394936 155388 394942 155400
rect 420362 155388 420368 155400
rect 420420 155388 420426 155440
rect 429286 155388 429292 155440
rect 429344 155428 429350 155440
rect 446674 155428 446680 155440
rect 429344 155400 446680 155428
rect 429344 155388 429350 155400
rect 446674 155388 446680 155400
rect 446732 155388 446738 155440
rect 296438 155360 296444 155372
rect 291304 155332 296444 155360
rect 296438 155320 296444 155332
rect 296496 155320 296502 155372
rect 339586 155360 339592 155372
rect 296548 155332 339592 155360
rect 8754 155252 8760 155304
rect 8812 155292 8818 155304
rect 125594 155292 125600 155304
rect 8812 155264 125600 155292
rect 8812 155252 8818 155264
rect 125594 155252 125600 155264
rect 125652 155252 125658 155304
rect 125778 155252 125784 155304
rect 125836 155292 125842 155304
rect 214834 155292 214840 155304
rect 125836 155264 214840 155292
rect 125836 155252 125842 155264
rect 214834 155252 214840 155264
rect 214892 155252 214898 155304
rect 219066 155252 219072 155304
rect 219124 155292 219130 155304
rect 286134 155292 286140 155304
rect 219124 155264 286140 155292
rect 219124 155252 219130 155264
rect 286134 155252 286140 155264
rect 286192 155252 286198 155304
rect 290550 155252 290556 155304
rect 290608 155292 290614 155304
rect 296548 155292 296576 155332
rect 339586 155320 339592 155332
rect 339644 155320 339650 155372
rect 345198 155320 345204 155372
rect 345256 155360 345262 155372
rect 382274 155360 382280 155372
rect 345256 155332 382280 155360
rect 345256 155320 345262 155332
rect 382274 155320 382280 155332
rect 382332 155320 382338 155372
rect 397362 155320 397368 155372
rect 397420 155360 397426 155372
rect 422294 155360 422300 155372
rect 397420 155332 422300 155360
rect 397420 155320 397426 155332
rect 422294 155320 422300 155332
rect 422352 155320 422358 155372
rect 424318 155320 424324 155372
rect 424376 155360 424382 155372
rect 441706 155360 441712 155372
rect 424376 155332 441712 155360
rect 424376 155320 424382 155332
rect 441706 155320 441712 155332
rect 441764 155320 441770 155372
rect 444466 155320 444472 155372
rect 444524 155360 444530 155372
rect 458174 155360 458180 155372
rect 444524 155332 458180 155360
rect 444524 155320 444530 155332
rect 458174 155320 458180 155332
rect 458232 155320 458238 155372
rect 290608 155264 296576 155292
rect 290608 155252 290614 155264
rect 296622 155252 296628 155304
rect 296680 155292 296686 155304
rect 338114 155292 338120 155304
rect 296680 155264 338120 155292
rect 296680 155252 296686 155264
rect 338114 155252 338120 155264
rect 338172 155252 338178 155304
rect 344370 155252 344376 155304
rect 344428 155292 344434 155304
rect 381446 155292 381452 155304
rect 344428 155264 381452 155292
rect 344428 155252 344434 155264
rect 381446 155252 381452 155264
rect 381504 155252 381510 155304
rect 383930 155252 383936 155304
rect 383988 155292 383994 155304
rect 411990 155292 411996 155304
rect 383988 155264 411996 155292
rect 383988 155252 383994 155264
rect 411990 155252 411996 155264
rect 412048 155252 412054 155304
rect 421742 155252 421748 155304
rect 421800 155292 421806 155304
rect 440878 155292 440884 155304
rect 421800 155264 440884 155292
rect 421800 155252 421806 155264
rect 440878 155252 440884 155264
rect 440936 155252 440942 155304
rect 441982 155252 441988 155304
rect 442040 155292 442046 155304
rect 442040 155264 453252 155292
rect 442040 155252 442046 155264
rect 1210 155184 1216 155236
rect 1268 155224 1274 155236
rect 118786 155224 118792 155236
rect 1268 155196 118792 155224
rect 1268 155184 1274 155196
rect 118786 155184 118792 155196
rect 118844 155184 118850 155236
rect 119522 155184 119528 155236
rect 119580 155224 119586 155236
rect 207566 155224 207572 155236
rect 119580 155196 207572 155224
rect 119580 155184 119586 155196
rect 207566 155184 207572 155196
rect 207624 155184 207630 155236
rect 216490 155184 216496 155236
rect 216548 155224 216554 155236
rect 283098 155224 283104 155236
rect 216548 155196 283104 155224
rect 216548 155184 216554 155196
rect 283098 155184 283104 155196
rect 283156 155184 283162 155236
rect 283834 155184 283840 155236
rect 283892 155224 283898 155236
rect 335538 155224 335544 155236
rect 283892 155196 335544 155224
rect 283892 155184 283898 155196
rect 335538 155184 335544 155196
rect 335596 155184 335602 155236
rect 343542 155184 343548 155236
rect 343600 155224 343606 155236
rect 380894 155224 380900 155236
rect 343600 155196 380900 155224
rect 343600 155184 343606 155196
rect 380894 155184 380900 155196
rect 380952 155184 380958 155236
rect 381354 155184 381360 155236
rect 381412 155224 381418 155236
rect 410058 155224 410064 155236
rect 381412 155196 410064 155224
rect 381412 155184 381418 155196
rect 410058 155184 410064 155196
rect 410116 155184 410122 155236
rect 410794 155184 410800 155236
rect 410852 155224 410858 155236
rect 432046 155224 432052 155236
rect 410852 155196 432052 155224
rect 410852 155184 410858 155196
rect 432046 155184 432052 155196
rect 432104 155184 432110 155236
rect 442810 155184 442816 155236
rect 442868 155224 442874 155236
rect 453224 155224 453252 155264
rect 456242 155252 456248 155304
rect 456300 155292 456306 155304
rect 467098 155292 467104 155304
rect 456300 155264 467104 155292
rect 456300 155252 456306 155264
rect 467098 155252 467104 155264
rect 467156 155252 467162 155304
rect 456334 155224 456340 155236
rect 442868 155196 451274 155224
rect 453224 155196 456340 155224
rect 442868 155184 442874 155196
rect 92474 155116 92480 155168
rect 92532 155156 92538 155168
rect 121086 155156 121092 155168
rect 92532 155128 121092 155156
rect 92532 155116 92538 155128
rect 121086 155116 121092 155128
rect 121144 155116 121150 155168
rect 150434 155116 150440 155168
rect 150492 155156 150498 155168
rect 229186 155156 229192 155168
rect 150492 155128 229192 155156
rect 150492 155116 150498 155128
rect 229186 155116 229192 155128
rect 229244 155116 229250 155168
rect 230014 155116 230020 155168
rect 230072 155156 230078 155168
rect 294046 155156 294052 155168
rect 230072 155128 294052 155156
rect 230072 155116 230078 155128
rect 294046 155116 294052 155128
rect 294104 155116 294110 155168
rect 330202 155116 330208 155168
rect 330260 155156 330266 155168
rect 356790 155156 356796 155168
rect 330260 155128 356796 155156
rect 330260 155116 330266 155128
rect 356790 155116 356796 155128
rect 356848 155116 356854 155168
rect 451246 155156 451274 155196
rect 456334 155184 456340 155196
rect 456392 155184 456398 155236
rect 456978 155156 456984 155168
rect 451246 155128 456984 155156
rect 456978 155116 456984 155128
rect 457036 155116 457042 155168
rect 128170 155048 128176 155100
rect 128228 155088 128234 155100
rect 198090 155088 198096 155100
rect 128228 155060 198096 155088
rect 128228 155048 128234 155060
rect 198090 155048 198096 155060
rect 198148 155048 198154 155100
rect 226610 155048 226616 155100
rect 226668 155088 226674 155100
rect 291194 155088 291200 155100
rect 226668 155060 291200 155088
rect 226668 155048 226674 155060
rect 291194 155048 291200 155060
rect 291252 155048 291258 155100
rect 291470 155048 291476 155100
rect 291528 155088 291534 155100
rect 330018 155088 330024 155100
rect 291528 155060 330024 155088
rect 291528 155048 291534 155060
rect 330018 155048 330024 155060
rect 330076 155048 330082 155100
rect 134886 154980 134892 155032
rect 134944 155020 134950 155032
rect 201862 155020 201868 155032
rect 134944 154992 201868 155020
rect 134944 154980 134950 154992
rect 201862 154980 201868 154992
rect 201920 154980 201926 155032
rect 269022 154980 269028 155032
rect 269080 155020 269086 155032
rect 317966 155020 317972 155032
rect 269080 154992 317972 155020
rect 269080 154980 269086 154992
rect 317966 154980 317972 154992
rect 318024 154980 318030 155032
rect 118142 154912 118148 154964
rect 118200 154952 118206 154964
rect 144822 154952 144828 154964
rect 118200 154924 144828 154952
rect 118200 154912 118206 154924
rect 144822 154912 144828 154924
rect 144880 154912 144886 154964
rect 157426 154912 157432 154964
rect 157484 154952 157490 154964
rect 225138 154952 225144 154964
rect 157484 154924 225144 154952
rect 157484 154912 157490 154924
rect 225138 154912 225144 154924
rect 225196 154912 225202 154964
rect 262122 154912 262128 154964
rect 262180 154952 262186 154964
rect 307938 154952 307944 154964
rect 262180 154924 307944 154952
rect 262180 154912 262186 154924
rect 307938 154912 307944 154924
rect 307996 154912 308002 154964
rect 105446 154504 105452 154556
rect 105504 154544 105510 154556
rect 199470 154544 199476 154556
rect 105504 154516 199476 154544
rect 105504 154504 105510 154516
rect 199470 154504 199476 154516
rect 199528 154504 199534 154556
rect 215662 154504 215668 154556
rect 215720 154544 215726 154556
rect 283558 154544 283564 154556
rect 215720 154516 283564 154544
rect 215720 154504 215726 154516
rect 283558 154504 283564 154516
rect 283616 154504 283622 154556
rect 284294 154504 284300 154556
rect 284352 154544 284358 154556
rect 320910 154544 320916 154556
rect 284352 154516 320916 154544
rect 284352 154504 284358 154516
rect 320910 154504 320916 154516
rect 320968 154504 320974 154556
rect 338390 154504 338396 154556
rect 338448 154544 338454 154556
rect 341978 154544 341984 154556
rect 338448 154516 341984 154544
rect 338448 154504 338454 154516
rect 341978 154504 341984 154516
rect 342036 154504 342042 154556
rect 463326 154504 463332 154556
rect 463384 154544 463390 154556
rect 468938 154544 468944 154556
rect 463384 154516 468944 154544
rect 463384 154504 463390 154516
rect 468938 154504 468944 154516
rect 468996 154504 469002 154556
rect 471790 154504 471796 154556
rect 471848 154544 471854 154556
rect 472986 154544 472992 154556
rect 471848 154516 472992 154544
rect 471848 154504 471854 154516
rect 472986 154504 472992 154516
rect 473044 154504 473050 154556
rect 103422 154436 103428 154488
rect 103480 154476 103486 154488
rect 197538 154476 197544 154488
rect 103480 154448 197544 154476
rect 103480 154436 103486 154448
rect 197538 154436 197544 154448
rect 197596 154436 197602 154488
rect 213178 154436 213184 154488
rect 213236 154476 213242 154488
rect 281626 154476 281632 154488
rect 213236 154448 281632 154476
rect 213236 154436 213242 154448
rect 281626 154436 281632 154448
rect 281684 154436 281690 154488
rect 313274 154436 313280 154488
rect 313332 154476 313338 154488
rect 358078 154476 358084 154488
rect 313332 154448 358084 154476
rect 313332 154436 313338 154448
rect 358078 154436 358084 154448
rect 358136 154436 358142 154488
rect 366818 154436 366824 154488
rect 366876 154476 366882 154488
rect 395338 154476 395344 154488
rect 366876 154448 395344 154476
rect 366876 154436 366882 154448
rect 395338 154436 395344 154448
rect 395396 154436 395402 154488
rect 92842 154368 92848 154420
rect 92900 154408 92906 154420
rect 189810 154408 189816 154420
rect 92900 154380 189816 154408
rect 92900 154368 92906 154380
rect 189810 154368 189816 154380
rect 189868 154368 189874 154420
rect 198734 154368 198740 154420
rect 198792 154408 198798 154420
rect 268838 154408 268844 154420
rect 198792 154380 268844 154408
rect 198792 154368 198798 154380
rect 268838 154368 268844 154380
rect 268896 154368 268902 154420
rect 281534 154368 281540 154420
rect 281592 154408 281598 154420
rect 333698 154408 333704 154420
rect 281592 154380 333704 154408
rect 281592 154368 281598 154380
rect 333698 154368 333704 154380
rect 333756 154368 333762 154420
rect 335078 154368 335084 154420
rect 335136 154408 335142 154420
rect 338942 154408 338948 154420
rect 335136 154380 338948 154408
rect 335136 154368 335142 154380
rect 338942 154368 338948 154380
rect 339000 154368 339006 154420
rect 340966 154368 340972 154420
rect 341024 154408 341030 154420
rect 379238 154408 379244 154420
rect 341024 154380 379244 154408
rect 341024 154368 341030 154380
rect 379238 154368 379244 154380
rect 379296 154368 379302 154420
rect 58342 154300 58348 154352
rect 58400 154340 58406 154352
rect 163498 154340 163504 154352
rect 58400 154312 163504 154340
rect 58400 154300 58406 154312
rect 163498 154300 163504 154312
rect 163556 154300 163562 154352
rect 192110 154300 192116 154352
rect 192168 154340 192174 154352
rect 265710 154340 265716 154352
rect 192168 154312 265716 154340
rect 192168 154300 192174 154312
rect 265710 154300 265716 154312
rect 265768 154300 265774 154352
rect 270310 154300 270316 154352
rect 270368 154340 270374 154352
rect 325326 154340 325332 154352
rect 270368 154312 325332 154340
rect 270368 154300 270374 154312
rect 325326 154300 325332 154312
rect 325384 154300 325390 154352
rect 333422 154300 333428 154352
rect 333480 154340 333486 154352
rect 373442 154340 373448 154352
rect 333480 154312 373448 154340
rect 333480 154300 333486 154312
rect 373442 154300 373448 154312
rect 373500 154300 373506 154352
rect 51626 154232 51632 154284
rect 51684 154272 51690 154284
rect 155954 154272 155960 154284
rect 51684 154244 155960 154272
rect 51684 154232 51690 154244
rect 155954 154232 155960 154244
rect 156012 154232 156018 154284
rect 188798 154232 188804 154284
rect 188856 154272 188862 154284
rect 263042 154272 263048 154284
rect 188856 154244 263048 154272
rect 188856 154232 188862 154244
rect 263042 154232 263048 154244
rect 263100 154232 263106 154284
rect 266998 154232 267004 154284
rect 267056 154272 267062 154284
rect 322842 154272 322848 154284
rect 267056 154244 322848 154272
rect 267056 154232 267062 154244
rect 322842 154232 322848 154244
rect 322900 154232 322906 154284
rect 326982 154232 326988 154284
rect 327040 154272 327046 154284
rect 368290 154272 368296 154284
rect 327040 154244 368296 154272
rect 327040 154232 327046 154244
rect 368290 154232 368296 154244
rect 368348 154232 368354 154284
rect 44910 154164 44916 154216
rect 44968 154204 44974 154216
rect 153194 154204 153200 154216
rect 44968 154176 153200 154204
rect 44968 154164 44974 154176
rect 153194 154164 153200 154176
rect 153252 154164 153258 154216
rect 154298 154164 154304 154216
rect 154356 154204 154362 154216
rect 182358 154204 182364 154216
rect 154356 154176 182364 154204
rect 154356 154164 154362 154176
rect 182358 154164 182364 154176
rect 182416 154164 182422 154216
rect 185394 154164 185400 154216
rect 185452 154204 185458 154216
rect 260466 154204 260472 154216
rect 185452 154176 260472 154204
rect 185452 154164 185458 154176
rect 260466 154164 260472 154176
rect 260524 154164 260530 154216
rect 263594 154164 263600 154216
rect 263652 154204 263658 154216
rect 320174 154204 320180 154216
rect 263652 154176 320180 154204
rect 263652 154164 263658 154176
rect 320174 154164 320180 154176
rect 320232 154164 320238 154216
rect 323302 154164 323308 154216
rect 323360 154204 323366 154216
rect 365714 154204 365720 154216
rect 323360 154176 365720 154204
rect 323360 154164 323366 154176
rect 365714 154164 365720 154176
rect 365772 154164 365778 154216
rect 371326 154164 371332 154216
rect 371384 154204 371390 154216
rect 402330 154204 402336 154216
rect 371384 154176 402336 154204
rect 371384 154164 371390 154176
rect 402330 154164 402336 154176
rect 402388 154164 402394 154216
rect 422570 154164 422576 154216
rect 422628 154204 422634 154216
rect 422628 154176 430068 154204
rect 422628 154164 422634 154176
rect 34790 154096 34796 154148
rect 34848 154136 34854 154148
rect 145558 154136 145564 154148
rect 34848 154108 145564 154136
rect 34848 154096 34854 154108
rect 145558 154096 145564 154108
rect 145616 154096 145622 154148
rect 147766 154096 147772 154148
rect 147824 154136 147830 154148
rect 177666 154136 177672 154148
rect 147824 154108 177672 154136
rect 147824 154096 147830 154108
rect 177666 154096 177672 154108
rect 177724 154096 177730 154148
rect 181990 154096 181996 154148
rect 182048 154136 182054 154148
rect 257890 154136 257896 154148
rect 182048 154108 257896 154136
rect 182048 154096 182054 154108
rect 257890 154096 257896 154108
rect 257948 154096 257954 154148
rect 257982 154096 257988 154148
rect 258040 154136 258046 154148
rect 315022 154136 315028 154148
rect 258040 154108 315028 154136
rect 258040 154096 258046 154108
rect 315022 154096 315028 154108
rect 315080 154096 315086 154148
rect 319990 154096 319996 154148
rect 320048 154136 320054 154148
rect 363230 154136 363236 154148
rect 320048 154108 363236 154136
rect 320048 154096 320054 154108
rect 363230 154096 363236 154108
rect 363288 154096 363294 154148
rect 368382 154096 368388 154148
rect 368440 154136 368446 154148
rect 399754 154136 399760 154148
rect 368440 154108 399760 154136
rect 368440 154096 368446 154108
rect 399754 154096 399760 154108
rect 399812 154096 399818 154148
rect 407482 154096 407488 154148
rect 407540 154136 407546 154148
rect 429930 154136 429936 154148
rect 407540 154108 429936 154136
rect 407540 154096 407546 154108
rect 429930 154096 429936 154108
rect 429988 154096 429994 154148
rect 25590 154028 25596 154080
rect 25648 154068 25654 154080
rect 138474 154068 138480 154080
rect 25648 154040 138480 154068
rect 25648 154028 25654 154040
rect 138474 154028 138480 154040
rect 138532 154028 138538 154080
rect 172422 154028 172428 154080
rect 172480 154068 172486 154080
rect 250162 154068 250168 154080
rect 172480 154040 250168 154068
rect 172480 154028 172486 154040
rect 250162 154028 250168 154040
rect 250220 154028 250226 154080
rect 250254 154028 250260 154080
rect 250312 154068 250318 154080
rect 309870 154068 309876 154080
rect 250312 154040 309876 154068
rect 250312 154028 250318 154040
rect 309870 154028 309876 154040
rect 309928 154028 309934 154080
rect 316586 154028 316592 154080
rect 316644 154068 316650 154080
rect 360654 154068 360660 154080
rect 316644 154040 360660 154068
rect 316644 154028 316650 154040
rect 360654 154028 360660 154040
rect 360712 154028 360718 154080
rect 394050 154068 394056 154080
rect 360764 154040 394056 154068
rect 20530 153960 20536 154012
rect 20588 154000 20594 154012
rect 134610 154000 134616 154012
rect 20588 153972 134616 154000
rect 20588 153960 20594 153972
rect 134610 153960 134616 153972
rect 134668 153960 134674 154012
rect 143350 153960 143356 154012
rect 143408 154000 143414 154012
rect 228358 154000 228364 154012
rect 143408 153972 228364 154000
rect 143408 153960 143414 153972
rect 228358 153960 228364 153972
rect 228416 153960 228422 154012
rect 243446 153960 243452 154012
rect 243504 154000 243510 154012
rect 304718 154000 304724 154012
rect 243504 153972 304724 154000
rect 243504 153960 243510 153972
rect 304718 153960 304724 153972
rect 304776 153960 304782 154012
rect 304810 153960 304816 154012
rect 304868 154000 304874 154012
rect 349062 154000 349068 154012
rect 304868 153972 349068 154000
rect 304868 153960 304874 153972
rect 349062 153960 349068 153972
rect 349120 153960 349126 154012
rect 360378 153960 360384 154012
rect 360436 154000 360442 154012
rect 360764 154000 360792 154040
rect 394050 154028 394056 154040
rect 394108 154028 394114 154080
rect 398190 154028 398196 154080
rect 398248 154068 398254 154080
rect 422938 154068 422944 154080
rect 398248 154040 422944 154068
rect 398248 154028 398254 154040
rect 422938 154028 422944 154040
rect 422996 154028 423002 154080
rect 430040 154068 430068 154176
rect 438854 154164 438860 154216
rect 438912 154204 438918 154216
rect 451826 154204 451832 154216
rect 438912 154176 451832 154204
rect 438912 154164 438918 154176
rect 451826 154164 451832 154176
rect 451884 154164 451890 154216
rect 431034 154096 431040 154148
rect 431092 154136 431098 154148
rect 447962 154136 447968 154148
rect 431092 154108 447968 154136
rect 431092 154096 431098 154108
rect 447962 154096 447968 154108
rect 448020 154096 448026 154148
rect 441430 154068 441436 154080
rect 430040 154040 441436 154068
rect 441430 154028 441436 154040
rect 441488 154028 441494 154080
rect 391474 154000 391480 154012
rect 360436 153972 360792 154000
rect 360948 153972 391480 154000
rect 360436 153960 360442 153972
rect 17126 153892 17132 153944
rect 17184 153932 17190 153944
rect 132034 153932 132040 153944
rect 17184 153904 132040 153932
rect 17184 153892 17190 153904
rect 132034 153892 132040 153904
rect 132092 153892 132098 153944
rect 132126 153892 132132 153944
rect 132184 153932 132190 153944
rect 217410 153932 217416 153944
rect 132184 153904 217416 153932
rect 132184 153892 132190 153904
rect 217410 153892 217416 153904
rect 217468 153892 217474 153944
rect 219894 153892 219900 153944
rect 219952 153932 219958 153944
rect 286778 153932 286784 153944
rect 219952 153904 286784 153932
rect 219952 153892 219958 153904
rect 286778 153892 286784 153904
rect 286836 153892 286842 153944
rect 286870 153892 286876 153944
rect 286928 153932 286934 153944
rect 337470 153932 337476 153944
rect 286928 153904 337476 153932
rect 286928 153892 286934 153904
rect 337470 153892 337476 153904
rect 337528 153892 337534 153944
rect 338022 153892 338028 153944
rect 338080 153932 338086 153944
rect 360838 153932 360844 153944
rect 338080 153904 360844 153932
rect 338080 153892 338086 153904
rect 360838 153892 360844 153904
rect 360896 153892 360902 153944
rect 13814 153824 13820 153876
rect 13872 153864 13878 153876
rect 129458 153864 129464 153876
rect 13872 153836 129464 153864
rect 13872 153824 13878 153836
rect 129458 153824 129464 153836
rect 129516 153824 129522 153876
rect 135714 153824 135720 153876
rect 135772 153864 135778 153876
rect 222562 153864 222568 153876
rect 135772 153836 222568 153864
rect 135772 153824 135778 153836
rect 222562 153824 222568 153836
rect 222620 153824 222626 153876
rect 233326 153824 233332 153876
rect 233384 153864 233390 153876
rect 297082 153864 297088 153876
rect 233384 153836 297088 153864
rect 233384 153824 233390 153836
rect 297082 153824 297088 153836
rect 297140 153824 297146 153876
rect 309962 153824 309968 153876
rect 310020 153864 310026 153876
rect 355502 153864 355508 153876
rect 310020 153836 355508 153864
rect 310020 153824 310026 153836
rect 355502 153824 355508 153836
rect 355560 153824 355566 153876
rect 357342 153824 357348 153876
rect 357400 153864 357406 153876
rect 360948 153864 360976 153972
rect 391474 153960 391480 153972
rect 391532 153960 391538 154012
rect 391842 153960 391848 154012
rect 391900 154000 391906 154012
rect 417142 154000 417148 154012
rect 391900 153972 417148 154000
rect 391900 153960 391906 153972
rect 417142 153960 417148 153972
rect 417200 153960 417206 154012
rect 425238 153960 425244 154012
rect 425296 154000 425302 154012
rect 443454 154000 443460 154012
rect 425296 153972 443460 154000
rect 425296 153960 425302 153972
rect 443454 153960 443460 153972
rect 443512 153960 443518 154012
rect 361022 153892 361028 153944
rect 361080 153932 361086 153944
rect 376570 153932 376576 153944
rect 361080 153904 376576 153932
rect 361080 153892 361086 153904
rect 376570 153892 376576 153904
rect 376628 153892 376634 153944
rect 380802 153892 380808 153944
rect 380860 153932 380866 153944
rect 409414 153932 409420 153944
rect 380860 153904 409420 153932
rect 380860 153892 380866 153904
rect 409414 153892 409420 153904
rect 409472 153892 409478 153944
rect 417510 153892 417516 153944
rect 417568 153932 417574 153944
rect 417568 153904 417924 153932
rect 417568 153892 417574 153904
rect 390186 153864 390192 153876
rect 357400 153836 360976 153864
rect 364306 153836 390192 153864
rect 357400 153824 357406 153836
rect 63402 153756 63408 153808
rect 63460 153796 63466 153808
rect 118694 153796 118700 153808
rect 63460 153768 118700 153796
rect 63460 153756 63466 153768
rect 118694 153756 118700 153768
rect 118752 153756 118758 153808
rect 119798 153756 119804 153808
rect 119856 153796 119862 153808
rect 208394 153796 208400 153808
rect 119856 153768 208400 153796
rect 119856 153756 119862 153768
rect 208394 153756 208400 153768
rect 208452 153756 208458 153808
rect 244274 153756 244280 153808
rect 244332 153796 244338 153808
rect 305362 153796 305368 153808
rect 244332 153768 305368 153796
rect 244332 153756 244338 153768
rect 305362 153756 305368 153768
rect 305420 153756 305426 153808
rect 305454 153756 305460 153808
rect 305512 153796 305518 153808
rect 336182 153796 336188 153808
rect 305512 153768 336188 153796
rect 305512 153756 305518 153768
rect 336182 153756 336188 153768
rect 336240 153756 336246 153808
rect 355318 153756 355324 153808
rect 355376 153796 355382 153808
rect 364306 153796 364334 153836
rect 390186 153824 390192 153836
rect 390244 153824 390250 153876
rect 391750 153824 391756 153876
rect 391808 153864 391814 153876
rect 417786 153864 417792 153876
rect 391808 153836 417792 153864
rect 391808 153824 391814 153836
rect 417786 153824 417792 153836
rect 417844 153824 417850 153876
rect 417896 153864 417924 153904
rect 418430 153892 418436 153944
rect 418488 153932 418494 153944
rect 438302 153932 438308 153944
rect 418488 153904 438308 153932
rect 418488 153892 418494 153904
rect 438302 153892 438308 153904
rect 438360 153892 438366 153944
rect 440234 153892 440240 153944
rect 440292 153932 440298 153944
rect 455046 153932 455052 153944
rect 440292 153904 455052 153932
rect 440292 153892 440298 153904
rect 455046 153892 455052 153904
rect 455104 153892 455110 153944
rect 437658 153864 437664 153876
rect 417896 153836 437664 153864
rect 437658 153824 437664 153836
rect 437716 153824 437722 153876
rect 453942 153824 453948 153876
rect 454000 153864 454006 153876
rect 462038 153864 462044 153876
rect 454000 153836 462044 153864
rect 454000 153824 454006 153836
rect 462038 153824 462044 153836
rect 462096 153824 462102 153876
rect 355376 153768 364334 153796
rect 355376 153756 355382 153768
rect 438578 153756 438584 153808
rect 438636 153796 438642 153808
rect 453758 153796 453764 153808
rect 438636 153768 453764 153796
rect 438636 153756 438642 153768
rect 453758 153756 453764 153768
rect 453816 153756 453822 153808
rect 77202 153688 77208 153740
rect 77260 153728 77266 153740
rect 121730 153728 121736 153740
rect 77260 153700 121736 153728
rect 77260 153688 77266 153700
rect 121730 153688 121736 153700
rect 121788 153688 121794 153740
rect 122650 153688 122656 153740
rect 122708 153728 122714 153740
rect 212258 153728 212264 153740
rect 122708 153700 212264 153728
rect 122708 153688 122714 153700
rect 212258 153688 212264 153700
rect 212316 153688 212322 153740
rect 263594 153688 263600 153740
rect 263652 153728 263658 153740
rect 263778 153728 263784 153740
rect 263652 153700 263784 153728
rect 263652 153688 263658 153700
rect 263778 153688 263784 153700
rect 263836 153688 263842 153740
rect 274634 153688 274640 153740
rect 274692 153728 274698 153740
rect 310514 153728 310520 153740
rect 274692 153700 310520 153728
rect 274692 153688 274698 153700
rect 310514 153688 310520 153700
rect 310572 153688 310578 153740
rect 128354 153620 128360 153672
rect 128412 153660 128418 153672
rect 159634 153660 159640 153672
rect 128412 153632 159640 153660
rect 128412 153620 128418 153632
rect 159634 153620 159640 153632
rect 159692 153620 159698 153672
rect 208486 153620 208492 153672
rect 208544 153660 208550 153672
rect 273898 153660 273904 153672
rect 208544 153632 273904 153660
rect 208544 153620 208550 153632
rect 273898 153620 273904 153632
rect 273956 153620 273962 153672
rect 279878 153620 279884 153672
rect 279936 153660 279942 153672
rect 315666 153660 315672 153672
rect 279936 153632 315672 153660
rect 279936 153620 279942 153632
rect 315666 153620 315672 153632
rect 315724 153620 315730 153672
rect 168558 153552 168564 153604
rect 168616 153592 168622 153604
rect 216214 153592 216220 153604
rect 168616 153564 216220 153592
rect 168616 153552 168622 153564
rect 216214 153552 216220 153564
rect 216272 153552 216278 153604
rect 296806 153552 296812 153604
rect 296864 153592 296870 153604
rect 325970 153592 325976 153604
rect 296864 153564 325976 153592
rect 296864 153552 296870 153564
rect 325970 153552 325976 153564
rect 326028 153552 326034 153604
rect 197354 153484 197360 153536
rect 197412 153524 197418 153536
rect 237834 153524 237840 153536
rect 197412 153496 237840 153524
rect 197412 153484 197418 153496
rect 237834 153484 237840 153496
rect 237892 153484 237898 153536
rect 237466 153212 237472 153264
rect 237524 153252 237530 153264
rect 240594 153252 240600 153264
rect 237524 153224 240600 153252
rect 237524 153212 237530 153224
rect 240594 153212 240600 153224
rect 240652 153212 240658 153264
rect 455322 153212 455328 153264
rect 455380 153252 455386 153264
rect 463326 153252 463332 153264
rect 455380 153224 463332 153252
rect 455380 153212 455386 153224
rect 463326 153212 463332 153224
rect 463384 153212 463390 153264
rect 118694 153144 118700 153196
rect 118752 153184 118758 153196
rect 167362 153184 167368 153196
rect 118752 153156 167368 153184
rect 118752 153144 118758 153156
rect 167362 153144 167368 153156
rect 167420 153144 167426 153196
rect 167730 153144 167736 153196
rect 167788 153184 167794 153196
rect 246942 153184 246948 153196
rect 167788 153156 246948 153184
rect 167788 153144 167794 153156
rect 246942 153144 246948 153156
rect 247000 153144 247006 153196
rect 247218 153144 247224 153196
rect 247276 153184 247282 153196
rect 259822 153184 259828 153196
rect 247276 153156 259828 153184
rect 247276 153144 247282 153156
rect 259822 153144 259828 153156
rect 259880 153144 259886 153196
rect 268930 153144 268936 153196
rect 268988 153184 268994 153196
rect 280338 153184 280344 153196
rect 268988 153156 280344 153184
rect 268988 153144 268994 153156
rect 280338 153144 280344 153156
rect 280396 153144 280402 153196
rect 281166 153144 281172 153196
rect 281224 153184 281230 153196
rect 290642 153184 290648 153196
rect 281224 153156 290648 153184
rect 281224 153144 281230 153156
rect 290642 153144 290648 153156
rect 290700 153144 290706 153196
rect 291102 153144 291108 153196
rect 291160 153184 291166 153196
rect 334342 153184 334348 153196
rect 291160 153156 334348 153184
rect 291160 153144 291166 153156
rect 334342 153144 334348 153156
rect 334400 153144 334406 153196
rect 338942 153144 338948 153196
rect 339000 153184 339006 153196
rect 339000 153156 345014 153184
rect 339000 153144 339006 153156
rect 63494 153076 63500 153128
rect 63552 153116 63558 153128
rect 144914 153116 144920 153128
rect 63552 153088 144920 153116
rect 63552 153076 63558 153088
rect 144914 153076 144920 153088
rect 144972 153076 144978 153128
rect 155954 153076 155960 153128
rect 156012 153116 156018 153128
rect 158346 153116 158352 153128
rect 156012 153088 158352 153116
rect 156012 153076 156018 153088
rect 158346 153076 158352 153088
rect 158404 153076 158410 153128
rect 161382 153076 161388 153128
rect 161440 153116 161446 153128
rect 241882 153116 241888 153128
rect 161440 153088 241888 153116
rect 161440 153076 161446 153088
rect 241882 153076 241888 153088
rect 241940 153076 241946 153128
rect 245654 153076 245660 153128
rect 245712 153116 245718 153128
rect 288066 153116 288072 153128
rect 245712 153088 288072 153116
rect 245712 153076 245718 153088
rect 288066 153076 288072 153088
rect 288124 153076 288130 153128
rect 292298 153076 292304 153128
rect 292356 153116 292362 153128
rect 339402 153116 339408 153128
rect 292356 153088 339408 153116
rect 292356 153076 292362 153088
rect 339402 153076 339408 153088
rect 339460 153076 339466 153128
rect 344986 153116 345014 153156
rect 355686 153144 355692 153196
rect 355744 153184 355750 153196
rect 357434 153184 357440 153196
rect 355744 153156 357440 153184
rect 355744 153144 355750 153156
rect 357434 153144 357440 153156
rect 357492 153144 357498 153196
rect 368566 153144 368572 153196
rect 368624 153184 368630 153196
rect 372798 153184 372804 153196
rect 368624 153156 372804 153184
rect 368624 153144 368630 153156
rect 372798 153144 372804 153156
rect 372856 153144 372862 153196
rect 385954 153144 385960 153196
rect 386012 153184 386018 153196
rect 388254 153184 388260 153196
rect 386012 153156 388260 153184
rect 386012 153144 386018 153156
rect 388254 153144 388260 153156
rect 388312 153144 388318 153196
rect 408494 153144 408500 153196
rect 408552 153184 408558 153196
rect 410702 153184 410708 153196
rect 408552 153156 410708 153184
rect 408552 153144 408558 153156
rect 410702 153144 410708 153156
rect 410760 153144 410766 153196
rect 435818 153144 435824 153196
rect 435876 153184 435882 153196
rect 439590 153184 439596 153196
rect 435876 153156 439596 153184
rect 435876 153144 435882 153156
rect 439590 153144 439596 153156
rect 439648 153144 439654 153196
rect 447134 153144 447140 153196
rect 447192 153184 447198 153196
rect 449250 153184 449256 153196
rect 447192 153156 449256 153184
rect 447192 153144 447198 153156
rect 449250 153144 449256 153156
rect 449308 153144 449314 153196
rect 452470 153144 452476 153196
rect 452528 153184 452534 153196
rect 460658 153184 460664 153196
rect 452528 153156 460664 153184
rect 452528 153144 452534 153156
rect 460658 153144 460664 153156
rect 460716 153144 460722 153196
rect 498286 153144 498292 153196
rect 498344 153184 498350 153196
rect 499298 153184 499304 153196
rect 498344 153156 499304 153184
rect 498344 153144 498350 153156
rect 499298 153144 499304 153156
rect 499356 153144 499362 153196
rect 505830 153144 505836 153196
rect 505888 153184 505894 153196
rect 506750 153184 506756 153196
rect 505888 153156 506756 153184
rect 505888 153144 505894 153156
rect 506750 153144 506756 153156
rect 506808 153144 506814 153196
rect 509694 153144 509700 153196
rect 509752 153184 509758 153196
rect 511718 153184 511724 153196
rect 509752 153156 511724 153184
rect 509752 153144 509758 153156
rect 511718 153144 511724 153156
rect 511776 153144 511782 153196
rect 512270 153144 512276 153196
rect 512328 153184 512334 153196
rect 514846 153184 514852 153196
rect 512328 153156 514852 153184
rect 512328 153144 512334 153156
rect 514846 153144 514852 153156
rect 514904 153144 514910 153196
rect 374730 153116 374736 153128
rect 344986 153088 374736 153116
rect 374730 153076 374736 153088
rect 374788 153076 374794 153128
rect 465534 153076 465540 153128
rect 465592 153116 465598 153128
rect 474274 153116 474280 153128
rect 465592 153088 474280 153116
rect 465592 153076 465598 153088
rect 474274 153076 474280 153088
rect 474332 153076 474338 153128
rect 506382 153076 506388 153128
rect 506440 153116 506446 153128
rect 507578 153116 507584 153128
rect 506440 153088 507584 153116
rect 506440 153076 506446 153088
rect 507578 153076 507584 153088
rect 507636 153076 507642 153128
rect 510982 153076 510988 153128
rect 511040 153116 511046 153128
rect 513466 153116 513472 153128
rect 511040 153088 513472 153116
rect 511040 153076 511046 153088
rect 513466 153076 513472 153088
rect 513524 153076 513530 153128
rect 514202 153076 514208 153128
rect 514260 153116 514266 153128
rect 517606 153116 517612 153128
rect 514260 153088 517612 153116
rect 514260 153076 514266 153088
rect 517606 153076 517612 153088
rect 517664 153076 517670 153128
rect 109034 153008 109040 153060
rect 109092 153048 109098 153060
rect 197998 153048 198004 153060
rect 109092 153020 198004 153048
rect 109092 153008 109098 153020
rect 197998 153008 198004 153020
rect 198056 153008 198062 153060
rect 198090 153008 198096 153060
rect 198148 153048 198154 153060
rect 216766 153048 216772 153060
rect 198148 153020 216772 153048
rect 198148 153008 198154 153020
rect 216766 153008 216772 153020
rect 216824 153008 216830 153060
rect 216858 153008 216864 153060
rect 216916 153048 216922 153060
rect 239306 153048 239312 153060
rect 216916 153020 239312 153048
rect 216916 153008 216922 153020
rect 239306 153008 239312 153020
rect 239364 153008 239370 153060
rect 239950 153008 239956 153060
rect 240008 153048 240014 153060
rect 293218 153048 293224 153060
rect 240008 153020 293224 153048
rect 240008 153008 240014 153020
rect 293218 153008 293224 153020
rect 293276 153008 293282 153060
rect 299382 153008 299388 153060
rect 299440 153048 299446 153060
rect 306006 153048 306012 153060
rect 299440 153020 306012 153048
rect 299440 153008 299446 153020
rect 306006 153008 306012 153020
rect 306064 153008 306070 153060
rect 318702 153008 318708 153060
rect 318760 153048 318766 153060
rect 360010 153048 360016 153060
rect 318760 153020 360016 153048
rect 318760 153008 318766 153020
rect 360010 153008 360016 153020
rect 360068 153008 360074 153060
rect 409966 153008 409972 153060
rect 410024 153048 410030 153060
rect 431862 153048 431868 153060
rect 410024 153020 431868 153048
rect 410024 153008 410030 153020
rect 431862 153008 431868 153020
rect 431920 153008 431926 153060
rect 462130 153008 462136 153060
rect 462188 153048 462194 153060
rect 471698 153048 471704 153060
rect 462188 153020 471704 153048
rect 462188 153008 462194 153020
rect 471698 153008 471704 153020
rect 471756 153008 471762 153060
rect 512914 153008 512920 153060
rect 512972 153048 512978 153060
rect 515950 153048 515956 153060
rect 512972 153020 515956 153048
rect 512972 153008 512978 153020
rect 515950 153008 515956 153020
rect 516008 153008 516014 153060
rect 117222 152940 117228 152992
rect 117280 152980 117286 152992
rect 208486 152980 208492 152992
rect 117280 152952 208492 152980
rect 117280 152940 117286 152952
rect 208486 152940 208492 152952
rect 208544 152940 208550 152992
rect 212626 152940 212632 152992
rect 212684 152980 212690 152992
rect 267550 152980 267556 152992
rect 212684 152952 267556 152980
rect 212684 152940 212690 152952
rect 267550 152940 267556 152952
rect 267608 152940 267614 152992
rect 271690 152940 271696 152992
rect 271748 152980 271754 152992
rect 324038 152980 324044 152992
rect 271748 152952 324044 152980
rect 271748 152940 271754 152952
rect 324038 152940 324044 152952
rect 324096 152940 324102 152992
rect 337746 152940 337752 152992
rect 337804 152980 337810 152992
rect 375374 152980 375380 152992
rect 337804 152952 375380 152980
rect 337804 152940 337810 152952
rect 375374 152940 375380 152952
rect 375432 152940 375438 152992
rect 389082 152940 389088 152992
rect 389140 152980 389146 152992
rect 413278 152980 413284 152992
rect 389140 152952 413284 152980
rect 389140 152940 389146 152952
rect 413278 152940 413284 152952
rect 413336 152940 413342 152992
rect 415854 152940 415860 152992
rect 415912 152980 415918 152992
rect 436370 152980 436376 152992
rect 415912 152952 436376 152980
rect 415912 152940 415918 152952
rect 436370 152940 436376 152952
rect 436428 152940 436434 152992
rect 454586 152940 454592 152992
rect 454644 152980 454650 152992
rect 454644 152952 456012 152980
rect 454644 152940 454650 152952
rect 113910 152872 113916 152924
rect 113968 152912 113974 152924
rect 205910 152912 205916 152924
rect 113968 152884 205916 152912
rect 113968 152872 113974 152884
rect 205910 152872 205916 152884
rect 205968 152872 205974 152924
rect 210878 152872 210884 152924
rect 210936 152912 210942 152924
rect 262398 152912 262404 152924
rect 210936 152884 262404 152912
rect 210936 152872 210942 152884
rect 262398 152872 262404 152884
rect 262456 152872 262462 152924
rect 263502 152872 263508 152924
rect 263560 152912 263566 152924
rect 318886 152912 318892 152924
rect 263560 152884 318892 152912
rect 263560 152872 263566 152884
rect 318886 152872 318892 152884
rect 318944 152872 318950 152924
rect 328270 152872 328276 152924
rect 328328 152912 328334 152924
rect 369578 152912 369584 152924
rect 328328 152884 369584 152912
rect 328328 152872 328334 152884
rect 369578 152872 369584 152884
rect 369636 152872 369642 152924
rect 372614 152872 372620 152924
rect 372672 152912 372678 152924
rect 380526 152912 380532 152924
rect 372672 152884 380532 152912
rect 372672 152872 372678 152884
rect 380526 152872 380532 152884
rect 380584 152872 380590 152924
rect 380986 152872 380992 152924
rect 381044 152912 381050 152924
rect 408126 152912 408132 152924
rect 381044 152884 408132 152912
rect 381044 152872 381050 152884
rect 408126 152872 408132 152884
rect 408184 152872 408190 152924
rect 412542 152872 412548 152924
rect 412600 152912 412606 152924
rect 433794 152912 433800 152924
rect 412600 152884 433800 152912
rect 412600 152872 412606 152884
rect 433794 152872 433800 152884
rect 433852 152872 433858 152924
rect 452838 152872 452844 152924
rect 452896 152912 452902 152924
rect 452896 152884 455920 152912
rect 452896 152872 452902 152884
rect 107470 152804 107476 152856
rect 107528 152844 107534 152856
rect 200758 152844 200764 152856
rect 107528 152816 200764 152844
rect 107528 152804 107534 152816
rect 200758 152804 200764 152816
rect 200816 152804 200822 152856
rect 207106 152804 207112 152856
rect 207164 152844 207170 152856
rect 212902 152844 212908 152856
rect 207164 152816 212908 152844
rect 207164 152804 207170 152816
rect 212902 152804 212908 152816
rect 212960 152804 212966 152856
rect 221734 152804 221740 152856
rect 221792 152844 221798 152856
rect 224494 152844 224500 152856
rect 221792 152816 224500 152844
rect 221792 152804 221798 152816
rect 224494 152804 224500 152816
rect 224552 152804 224558 152856
rect 224586 152804 224592 152856
rect 224644 152844 224650 152856
rect 244366 152844 244372 152856
rect 224644 152816 244372 152844
rect 224644 152804 224650 152816
rect 244366 152804 244372 152816
rect 244424 152804 244430 152856
rect 244550 152804 244556 152856
rect 244608 152844 244614 152856
rect 303522 152844 303528 152856
rect 244608 152816 303528 152844
rect 244608 152804 244614 152816
rect 303522 152804 303528 152816
rect 303580 152804 303586 152856
rect 304994 152804 305000 152856
rect 305052 152844 305058 152856
rect 316310 152844 316316 152856
rect 305052 152816 316316 152844
rect 305052 152804 305058 152816
rect 316310 152804 316316 152816
rect 316368 152804 316374 152856
rect 322750 152804 322756 152856
rect 322808 152844 322814 152856
rect 365162 152844 365168 152856
rect 322808 152816 365168 152844
rect 322808 152804 322814 152816
rect 365162 152804 365168 152816
rect 365220 152804 365226 152856
rect 374270 152804 374276 152856
rect 374328 152844 374334 152856
rect 402974 152844 402980 152856
rect 374328 152816 402980 152844
rect 374328 152804 374334 152816
rect 402974 152804 402980 152816
rect 403032 152804 403038 152856
rect 403250 152804 403256 152856
rect 403308 152844 403314 152856
rect 426802 152844 426808 152856
rect 403308 152816 426808 152844
rect 403308 152804 403314 152816
rect 426802 152804 426808 152816
rect 426860 152804 426866 152856
rect 97074 152736 97080 152788
rect 97132 152776 97138 152788
rect 193030 152776 193036 152788
rect 97132 152748 193036 152776
rect 97132 152736 97138 152748
rect 193030 152736 193036 152748
rect 193088 152736 193094 152788
rect 193122 152736 193128 152788
rect 193180 152776 193186 152788
rect 229002 152776 229008 152788
rect 193180 152748 229008 152776
rect 193180 152736 193186 152748
rect 229002 152736 229008 152748
rect 229060 152736 229066 152788
rect 230382 152736 230388 152788
rect 230440 152776 230446 152788
rect 249518 152776 249524 152788
rect 230440 152748 249524 152776
rect 230440 152736 230446 152748
rect 249518 152736 249524 152748
rect 249576 152736 249582 152788
rect 249610 152736 249616 152788
rect 249668 152776 249674 152788
rect 308582 152776 308588 152788
rect 249668 152748 308588 152776
rect 249668 152736 249674 152748
rect 308582 152736 308588 152748
rect 308640 152736 308646 152788
rect 309042 152736 309048 152788
rect 309100 152776 309106 152788
rect 354858 152776 354864 152788
rect 309100 152748 354864 152776
rect 309100 152736 309106 152748
rect 354858 152736 354864 152748
rect 354916 152736 354922 152788
rect 358906 152736 358912 152788
rect 358964 152776 358970 152788
rect 390830 152776 390836 152788
rect 358964 152748 390836 152776
rect 358964 152736 358970 152748
rect 390830 152736 390836 152748
rect 390888 152736 390894 152788
rect 391566 152736 391572 152788
rect 391624 152776 391630 152788
rect 416498 152776 416504 152788
rect 391624 152748 416504 152776
rect 391624 152736 391630 152748
rect 416498 152736 416504 152748
rect 416556 152736 416562 152788
rect 416682 152736 416688 152788
rect 416740 152776 416746 152788
rect 437014 152776 437020 152788
rect 416740 152748 437020 152776
rect 416740 152736 416746 152748
rect 437014 152736 437020 152748
rect 437072 152736 437078 152788
rect 444282 152736 444288 152788
rect 444340 152776 444346 152788
rect 453114 152776 453120 152788
rect 444340 152748 453120 152776
rect 444340 152736 444346 152748
rect 453114 152736 453120 152748
rect 453172 152736 453178 152788
rect 455414 152736 455420 152788
rect 455472 152776 455478 152788
rect 455892 152776 455920 152884
rect 455984 152844 456012 152952
rect 460842 152940 460848 152992
rect 460900 152980 460906 152992
rect 470318 152980 470324 152992
rect 460900 152952 470324 152980
rect 460900 152940 460906 152952
rect 470318 152940 470324 152952
rect 470376 152940 470382 152992
rect 514846 152940 514852 152992
rect 514904 152980 514910 152992
rect 518526 152980 518532 152992
rect 514904 152952 518532 152980
rect 514904 152940 514910 152952
rect 518526 152940 518532 152952
rect 518584 152940 518590 152992
rect 457070 152872 457076 152924
rect 457128 152912 457134 152924
rect 467834 152912 467840 152924
rect 457128 152884 467840 152912
rect 457128 152872 457134 152884
rect 467834 152872 467840 152884
rect 467892 152872 467898 152924
rect 469122 152872 469128 152924
rect 469180 152912 469186 152924
rect 476850 152912 476856 152924
rect 469180 152884 476856 152912
rect 469180 152872 469186 152884
rect 476850 152872 476856 152884
rect 476908 152872 476914 152924
rect 465902 152844 465908 152856
rect 455984 152816 465908 152844
rect 465902 152804 465908 152816
rect 465960 152804 465966 152856
rect 469674 152804 469680 152856
rect 469732 152844 469738 152856
rect 477494 152844 477500 152856
rect 469732 152816 477500 152844
rect 469732 152804 469738 152816
rect 477494 152804 477500 152816
rect 477552 152804 477558 152856
rect 510338 152804 510344 152856
rect 510396 152844 510402 152856
rect 511994 152844 512000 152856
rect 510396 152816 512000 152844
rect 510396 152804 510402 152816
rect 511994 152804 512000 152816
rect 512052 152804 512058 152856
rect 518066 152804 518072 152856
rect 518124 152844 518130 152856
rect 522666 152844 522672 152856
rect 518124 152816 522672 152844
rect 518124 152804 518130 152816
rect 522666 152804 522672 152816
rect 522724 152804 522730 152856
rect 464614 152776 464620 152788
rect 455472 152748 455828 152776
rect 455892 152748 464620 152776
rect 455472 152736 455478 152748
rect 90358 152668 90364 152720
rect 90416 152708 90422 152720
rect 187878 152708 187884 152720
rect 90416 152680 187884 152708
rect 90416 152668 90422 152680
rect 187878 152668 187884 152680
rect 187936 152668 187942 152720
rect 201862 152668 201868 152720
rect 201920 152708 201926 152720
rect 221918 152708 221924 152720
rect 201920 152680 221924 152708
rect 201920 152668 201926 152680
rect 221918 152668 221924 152680
rect 221976 152668 221982 152720
rect 223942 152668 223948 152720
rect 224000 152708 224006 152720
rect 282914 152708 282920 152720
rect 224000 152680 282920 152708
rect 224000 152668 224006 152680
rect 282914 152668 282920 152680
rect 282972 152668 282978 152720
rect 284386 152668 284392 152720
rect 284444 152708 284450 152720
rect 295794 152708 295800 152720
rect 284444 152680 295800 152708
rect 284444 152668 284450 152680
rect 295794 152668 295800 152680
rect 295852 152668 295858 152720
rect 295886 152668 295892 152720
rect 295944 152708 295950 152720
rect 344554 152708 344560 152720
rect 295944 152680 344560 152708
rect 295944 152668 295950 152680
rect 344554 152668 344560 152680
rect 344612 152668 344618 152720
rect 362954 152668 362960 152720
rect 363012 152708 363018 152720
rect 395982 152708 395988 152720
rect 363012 152680 395988 152708
rect 363012 152668 363018 152680
rect 395982 152668 395988 152680
rect 396040 152668 396046 152720
rect 396626 152668 396632 152720
rect 396684 152708 396690 152720
rect 421650 152708 421656 152720
rect 396684 152680 421656 152708
rect 396684 152668 396690 152680
rect 421650 152668 421656 152680
rect 421708 152668 421714 152720
rect 445478 152668 445484 152720
rect 445536 152708 445542 152720
rect 455690 152708 455696 152720
rect 445536 152680 455696 152708
rect 445536 152668 445542 152680
rect 455690 152668 455696 152680
rect 455748 152668 455754 152720
rect 455800 152708 455828 152748
rect 464614 152736 464620 152748
rect 464672 152736 464678 152788
rect 467190 152736 467196 152788
rect 467248 152776 467254 152788
rect 475562 152776 475568 152788
rect 467248 152748 475568 152776
rect 467248 152736 467254 152748
rect 475562 152736 475568 152748
rect 475620 152736 475626 152788
rect 466546 152708 466552 152720
rect 455800 152680 466552 152708
rect 466546 152668 466552 152680
rect 466604 152668 466610 152720
rect 468018 152668 468024 152720
rect 468076 152708 468082 152720
rect 476206 152708 476212 152720
rect 468076 152680 476212 152708
rect 468076 152668 468082 152680
rect 476206 152668 476212 152680
rect 476264 152668 476270 152720
rect 73522 152600 73528 152652
rect 73580 152640 73586 152652
rect 175090 152640 175096 152652
rect 73580 152612 175096 152640
rect 73580 152600 73586 152612
rect 175090 152600 175096 152612
rect 175148 152600 175154 152652
rect 212350 152600 212356 152652
rect 212408 152640 212414 152652
rect 272702 152640 272708 152652
rect 212408 152612 272708 152640
rect 212408 152600 212414 152612
rect 272702 152600 272708 152612
rect 272760 152600 272766 152652
rect 278682 152600 278688 152652
rect 278740 152640 278746 152652
rect 329190 152640 329196 152652
rect 278740 152612 329196 152640
rect 278740 152600 278746 152612
rect 329190 152600 329196 152612
rect 329248 152600 329254 152652
rect 329282 152600 329288 152652
rect 329340 152640 329346 152652
rect 370222 152640 370228 152652
rect 329340 152612 370228 152640
rect 329340 152600 329346 152612
rect 370222 152600 370228 152612
rect 370280 152600 370286 152652
rect 376662 152600 376668 152652
rect 376720 152640 376726 152652
rect 406194 152640 406200 152652
rect 376720 152612 406200 152640
rect 376720 152600 376726 152612
rect 406194 152600 406200 152612
rect 406252 152600 406258 152652
rect 406930 152600 406936 152652
rect 406988 152640 406994 152652
rect 428642 152640 428648 152652
rect 406988 152612 428648 152640
rect 406988 152600 406994 152612
rect 428642 152600 428648 152612
rect 428700 152600 428706 152652
rect 450354 152600 450360 152652
rect 450412 152640 450418 152652
rect 462682 152640 462688 152652
rect 450412 152612 462688 152640
rect 450412 152600 450418 152612
rect 462682 152600 462688 152612
rect 462740 152600 462746 152652
rect 462958 152600 462964 152652
rect 463016 152640 463022 152652
rect 472342 152640 472348 152652
rect 463016 152612 472348 152640
rect 463016 152600 463022 152612
rect 472342 152600 472348 152612
rect 472400 152600 472406 152652
rect 518802 152600 518808 152652
rect 518860 152640 518866 152652
rect 523494 152640 523500 152652
rect 518860 152612 523500 152640
rect 518860 152600 518866 152612
rect 523494 152600 523500 152612
rect 523552 152600 523558 152652
rect 23382 152532 23388 152584
rect 23440 152572 23446 152584
rect 136542 152572 136548 152584
rect 23440 152544 136548 152572
rect 23440 152532 23446 152544
rect 136542 152532 136548 152544
rect 136600 152532 136606 152584
rect 147582 152532 147588 152584
rect 147640 152572 147646 152584
rect 231578 152572 231584 152584
rect 147640 152544 231584 152572
rect 147640 152532 147646 152544
rect 231578 152532 231584 152544
rect 231636 152532 231642 152584
rect 242434 152532 242440 152584
rect 242492 152572 242498 152584
rect 254670 152572 254676 152584
rect 242492 152544 254676 152572
rect 242492 152532 242498 152544
rect 254670 152532 254676 152544
rect 254728 152532 254734 152584
rect 255222 152532 255228 152584
rect 255280 152572 255286 152584
rect 313734 152572 313740 152584
rect 255280 152544 313740 152572
rect 255280 152532 255286 152544
rect 313734 152532 313740 152544
rect 313792 152532 313798 152584
rect 314930 152532 314936 152584
rect 314988 152572 314994 152584
rect 359366 152572 359372 152584
rect 314988 152544 359372 152572
rect 314988 152532 314994 152544
rect 359366 152532 359372 152544
rect 359424 152532 359430 152584
rect 365438 152532 365444 152584
rect 365496 152572 365502 152584
rect 397822 152572 397828 152584
rect 365496 152544 397828 152572
rect 365496 152532 365502 152544
rect 397822 152532 397828 152544
rect 397880 152532 397886 152584
rect 399018 152532 399024 152584
rect 399076 152572 399082 152584
rect 423582 152572 423588 152584
rect 399076 152544 423588 152572
rect 399076 152532 399082 152544
rect 423582 152532 423588 152544
rect 423640 152532 423646 152584
rect 446950 152532 446956 152584
rect 447008 152572 447014 152584
rect 460106 152572 460112 152584
rect 447008 152544 460112 152572
rect 447008 152532 447014 152544
rect 460106 152532 460112 152544
rect 460164 152532 460170 152584
rect 469766 152572 469772 152584
rect 460216 152544 469772 152572
rect 6270 152464 6276 152516
rect 6328 152504 6334 152516
rect 123662 152504 123668 152516
rect 6328 152476 123668 152504
rect 6328 152464 6334 152476
rect 123662 152464 123668 152476
rect 123720 152464 123726 152516
rect 125686 152464 125692 152516
rect 125744 152504 125750 152516
rect 127526 152504 127532 152516
rect 125744 152476 127532 152504
rect 125744 152464 125750 152476
rect 127526 152464 127532 152476
rect 127584 152464 127590 152516
rect 134058 152464 134064 152516
rect 134116 152504 134122 152516
rect 221274 152504 221280 152516
rect 134116 152476 221280 152504
rect 134116 152464 134122 152476
rect 221274 152464 221280 152476
rect 221332 152464 221338 152516
rect 222010 152464 222016 152516
rect 222068 152504 222074 152516
rect 224586 152504 224592 152516
rect 222068 152476 224592 152504
rect 222068 152464 222074 152476
rect 224586 152464 224592 152476
rect 224644 152464 224650 152516
rect 234982 152464 234988 152516
rect 235040 152504 235046 152516
rect 298370 152504 298376 152516
rect 235040 152476 298376 152504
rect 235040 152464 235046 152476
rect 298370 152464 298376 152476
rect 298428 152464 298434 152516
rect 302326 152464 302332 152516
rect 302384 152504 302390 152516
rect 349706 152504 349712 152516
rect 302384 152476 349712 152504
rect 302384 152464 302390 152476
rect 349706 152464 349712 152476
rect 349764 152464 349770 152516
rect 385586 152504 385592 152516
rect 354646 152476 385592 152504
rect 109126 152396 109132 152448
rect 109184 152436 109190 152448
rect 122374 152436 122380 152448
rect 109184 152408 122380 152436
rect 109184 152396 109190 152408
rect 122374 152396 122380 152408
rect 122432 152396 122438 152448
rect 124122 152396 124128 152448
rect 124180 152436 124186 152448
rect 128814 152436 128820 152448
rect 124180 152408 128820 152436
rect 124180 152396 124186 152408
rect 128814 152396 128820 152408
rect 128872 152396 128878 152448
rect 129826 152396 129832 152448
rect 129884 152436 129890 152448
rect 139118 152436 139124 152448
rect 129884 152408 139124 152436
rect 129884 152396 129890 152408
rect 139118 152396 139124 152408
rect 139176 152396 139182 152448
rect 143074 152396 143080 152448
rect 143132 152436 143138 152448
rect 216122 152436 216128 152448
rect 143132 152408 216128 152436
rect 143132 152396 143138 152408
rect 216122 152396 216128 152408
rect 216180 152396 216186 152448
rect 216214 152396 216220 152448
rect 216272 152436 216278 152448
rect 247586 152436 247592 152448
rect 216272 152408 247592 152436
rect 216272 152396 216278 152408
rect 247586 152396 247592 152408
rect 247644 152396 247650 152448
rect 256694 152396 256700 152448
rect 256752 152436 256758 152448
rect 301590 152436 301596 152448
rect 256752 152408 301596 152436
rect 256752 152396 256758 152408
rect 301590 152396 301596 152408
rect 301648 152396 301654 152448
rect 301682 152396 301688 152448
rect 301740 152436 301746 152448
rect 311158 152436 311164 152448
rect 301740 152408 311164 152436
rect 301740 152396 301746 152408
rect 311158 152396 311164 152408
rect 311216 152396 311222 152448
rect 321462 152436 321468 152448
rect 311866 152408 321468 152436
rect 144822 152328 144828 152380
rect 144880 152368 144886 152380
rect 209130 152368 209136 152380
rect 144880 152340 209136 152368
rect 144880 152328 144886 152340
rect 209130 152328 209136 152340
rect 209188 152328 209194 152380
rect 230750 152328 230756 152380
rect 230808 152368 230814 152380
rect 257246 152368 257252 152380
rect 230808 152340 257252 152368
rect 230808 152328 230814 152340
rect 257246 152328 257252 152340
rect 257304 152328 257310 152380
rect 260742 152328 260748 152380
rect 260800 152368 260806 152380
rect 270126 152368 270132 152380
rect 260800 152340 270132 152368
rect 260800 152328 260806 152340
rect 270126 152328 270132 152340
rect 270184 152328 270190 152380
rect 272518 152328 272524 152380
rect 272576 152368 272582 152380
rect 285490 152368 285496 152380
rect 272576 152340 285496 152368
rect 272576 152328 272582 152340
rect 285490 152328 285496 152340
rect 285548 152328 285554 152380
rect 109218 152260 109224 152312
rect 109276 152300 109282 152312
rect 157058 152300 157064 152312
rect 109276 152272 157064 152300
rect 109276 152260 109282 152272
rect 157058 152260 157064 152272
rect 157116 152260 157122 152312
rect 157334 152260 157340 152312
rect 157392 152300 157398 152312
rect 160922 152300 160928 152312
rect 157392 152272 160928 152300
rect 157392 152260 157398 152272
rect 160922 152260 160928 152272
rect 160980 152260 160986 152312
rect 174906 152260 174912 152312
rect 174964 152300 174970 152312
rect 226426 152300 226432 152312
rect 174964 152272 226432 152300
rect 174964 152260 174970 152272
rect 226426 152260 226432 152272
rect 226484 152260 226490 152312
rect 256786 152260 256792 152312
rect 256844 152300 256850 152312
rect 264974 152300 264980 152312
rect 256844 152272 264980 152300
rect 256844 152260 256850 152272
rect 264974 152260 264980 152272
rect 265032 152260 265038 152312
rect 265066 152260 265072 152312
rect 265124 152300 265130 152312
rect 275278 152300 275284 152312
rect 265124 152272 275284 152300
rect 265124 152260 265130 152272
rect 275278 152260 275284 152272
rect 275336 152260 275342 152312
rect 288250 152260 288256 152312
rect 288308 152300 288314 152312
rect 300946 152300 300952 152312
rect 288308 152272 300952 152300
rect 288308 152260 288314 152272
rect 300946 152260 300952 152272
rect 301004 152260 301010 152312
rect 311066 152260 311072 152312
rect 311124 152300 311130 152312
rect 311866 152300 311894 152408
rect 321462 152396 321468 152408
rect 321520 152396 321526 152448
rect 349430 152396 349436 152448
rect 349488 152436 349494 152448
rect 354646 152436 354674 152476
rect 385586 152464 385592 152476
rect 385644 152464 385650 152516
rect 392302 152464 392308 152516
rect 392360 152504 392366 152516
rect 418430 152504 418436 152516
rect 392360 152476 418436 152504
rect 392360 152464 392366 152476
rect 418430 152464 418436 152476
rect 418488 152464 418494 152516
rect 437382 152464 437388 152516
rect 437440 152504 437446 152516
rect 452470 152504 452476 152516
rect 437440 152476 452476 152504
rect 437440 152464 437446 152476
rect 452470 152464 452476 152476
rect 452528 152464 452534 152516
rect 459646 152464 459652 152516
rect 459704 152504 459710 152516
rect 460216 152504 460244 152544
rect 469766 152532 469772 152544
rect 469824 152532 469830 152584
rect 470502 152532 470508 152584
rect 470560 152572 470566 152584
rect 478138 152572 478144 152584
rect 470560 152544 478144 152572
rect 470560 152532 470566 152544
rect 478138 152532 478144 152544
rect 478196 152532 478202 152584
rect 463970 152504 463976 152516
rect 459704 152476 460244 152504
rect 460906 152476 463976 152504
rect 459704 152464 459710 152476
rect 349488 152408 354674 152436
rect 349488 152396 349494 152408
rect 414290 152396 414296 152448
rect 414348 152436 414354 152448
rect 415854 152436 415860 152448
rect 414348 152408 415860 152436
rect 414348 152396 414354 152408
rect 415854 152396 415860 152408
rect 415912 152396 415918 152448
rect 452010 152396 452016 152448
rect 452068 152436 452074 152448
rect 460906 152436 460934 152476
rect 463970 152464 463976 152476
rect 464028 152464 464034 152516
rect 464982 152464 464988 152516
rect 465040 152504 465046 152516
rect 473630 152504 473636 152516
rect 465040 152476 473636 152504
rect 465040 152464 465046 152476
rect 473630 152464 473636 152476
rect 473688 152464 473694 152516
rect 517422 152464 517428 152516
rect 517480 152504 517486 152516
rect 521838 152504 521844 152516
rect 517480 152476 521844 152504
rect 517480 152464 517486 152476
rect 521838 152464 521844 152476
rect 521896 152464 521902 152516
rect 452068 152408 460934 152436
rect 452068 152396 452074 152408
rect 507118 152328 507124 152380
rect 507176 152368 507182 152380
rect 507854 152368 507860 152380
rect 507176 152340 507860 152368
rect 507176 152328 507182 152340
rect 507854 152328 507860 152340
rect 507912 152328 507918 152380
rect 511626 152328 511632 152380
rect 511684 152368 511690 152380
rect 513558 152368 513564 152380
rect 511684 152340 513564 152368
rect 511684 152328 511690 152340
rect 513558 152328 513564 152340
rect 513616 152328 513622 152380
rect 311124 152272 311894 152300
rect 311124 152260 311130 152272
rect 54202 152192 54208 152244
rect 54260 152232 54266 152244
rect 89162 152232 89168 152244
rect 54260 152204 89168 152232
rect 54260 152192 54266 152204
rect 89162 152192 89168 152204
rect 89220 152192 89226 152244
rect 204162 152192 204168 152244
rect 204220 152232 204226 152244
rect 252094 152232 252100 152244
rect 204220 152204 252100 152232
rect 204220 152192 204226 152204
rect 252094 152192 252100 152204
rect 252152 152192 252158 152244
rect 513558 152192 513564 152244
rect 513616 152232 513622 152244
rect 516134 152232 516140 152244
rect 513616 152204 516140 152232
rect 513616 152192 513622 152204
rect 516134 152192 516140 152204
rect 516192 152192 516198 152244
rect 23290 152124 23296 152176
rect 23348 152164 23354 152176
rect 110046 152164 110052 152176
rect 23348 152136 110052 152164
rect 23348 152124 23354 152136
rect 110046 152124 110052 152136
rect 110104 152124 110110 152176
rect 71406 152056 71412 152108
rect 71464 152096 71470 152108
rect 82814 152096 82820 152108
rect 71464 152068 82820 152096
rect 71464 152056 71470 152068
rect 82814 152056 82820 152068
rect 82872 152056 82878 152108
rect 95510 152056 95516 152108
rect 95568 152096 95574 152108
rect 114370 152096 114376 152108
rect 95568 152068 114376 152096
rect 95568 152056 95574 152068
rect 114370 152056 114376 152068
rect 114428 152056 114434 152108
rect 88610 151988 88616 152040
rect 88668 152028 88674 152040
rect 110138 152028 110144 152040
rect 88668 152000 110144 152028
rect 88668 151988 88674 152000
rect 110138 151988 110144 152000
rect 110196 151988 110202 152040
rect 515490 151988 515496 152040
rect 515548 152028 515554 152040
rect 518986 152028 518992 152040
rect 515548 152000 518992 152028
rect 515548 151988 515554 152000
rect 518986 151988 518992 152000
rect 519044 151988 519050 152040
rect 33594 151920 33600 151972
rect 33652 151960 33658 151972
rect 110230 151960 110236 151972
rect 33652 151932 110236 151960
rect 33652 151920 33658 151932
rect 110230 151920 110236 151932
rect 110288 151920 110294 151972
rect 138014 151920 138020 151972
rect 138072 151960 138078 151972
rect 144270 151960 144276 151972
rect 138072 151932 144276 151960
rect 138072 151920 138078 151932
rect 144270 151920 144276 151932
rect 144328 151920 144334 151972
rect 507762 151920 507768 151972
rect 507820 151960 507826 151972
rect 509234 151960 509240 151972
rect 507820 151932 509240 151960
rect 507820 151920 507826 151932
rect 509234 151920 509240 151932
rect 509292 151920 509298 151972
rect 516778 151920 516784 151972
rect 516836 151960 516842 151972
rect 520274 151960 520280 151972
rect 516836 151932 520280 151960
rect 516836 151920 516842 151932
rect 520274 151920 520280 151932
rect 520332 151920 520338 151972
rect 26694 151852 26700 151904
rect 26752 151892 26758 151904
rect 109770 151892 109776 151904
rect 26752 151864 109776 151892
rect 26752 151852 26758 151864
rect 109770 151852 109776 151864
rect 109828 151852 109834 151904
rect 127618 151852 127624 151904
rect 127676 151892 127682 151904
rect 133966 151892 133972 151904
rect 127676 151864 133972 151892
rect 127676 151852 127682 151864
rect 133966 151852 133972 151864
rect 134024 151852 134030 151904
rect 139486 151852 139492 151904
rect 139544 151892 139550 151904
rect 142982 151892 142988 151904
rect 139544 151864 142988 151892
rect 139544 151852 139550 151864
rect 142982 151852 142988 151864
rect 143040 151852 143046 151904
rect 194318 151852 194324 151904
rect 194376 151892 194382 151904
rect 202690 151892 202696 151904
rect 194376 151864 202696 151892
rect 194376 151852 194382 151864
rect 202690 151852 202696 151864
rect 202748 151852 202754 151904
rect 320726 151852 320732 151904
rect 320784 151892 320790 151904
rect 326614 151892 326620 151904
rect 320784 151864 326620 151892
rect 320784 151852 320790 151864
rect 326614 151852 326620 151864
rect 326672 151852 326678 151904
rect 332594 151852 332600 151904
rect 332652 151892 332658 151904
rect 336826 151892 336832 151904
rect 332652 151864 336832 151892
rect 332652 151852 332658 151864
rect 336826 151852 336832 151864
rect 336884 151852 336890 151904
rect 343634 151852 343640 151904
rect 343692 151892 343698 151904
rect 347130 151892 347136 151904
rect 343692 151864 347136 151892
rect 343692 151852 343698 151864
rect 347130 151852 347136 151864
rect 347188 151852 347194 151904
rect 359458 151852 359464 151904
rect 359516 151892 359522 151904
rect 364518 151892 364524 151904
rect 359516 151864 364524 151892
rect 359516 151852 359522 151864
rect 364518 151852 364524 151864
rect 364576 151852 364582 151904
rect 508406 151852 508412 151904
rect 508464 151892 508470 151904
rect 510062 151892 510068 151904
rect 508464 151864 510068 151892
rect 508464 151852 508470 151864
rect 510062 151852 510068 151864
rect 510120 151852 510126 151904
rect 81710 151784 81716 151836
rect 81768 151824 81774 151836
rect 97718 151824 97724 151836
rect 81768 151796 97724 151824
rect 81768 151784 81774 151796
rect 97718 151784 97724 151796
rect 97776 151784 97782 151836
rect 102318 151784 102324 151836
rect 102376 151824 102382 151836
rect 110322 151824 110328 151836
rect 102376 151796 110328 151824
rect 102376 151784 102382 151796
rect 110322 151784 110328 151796
rect 110380 151784 110386 151836
rect 208394 151784 208400 151836
rect 208452 151824 208458 151836
rect 210418 151824 210424 151836
rect 208452 151796 210424 151824
rect 208452 151784 208458 151796
rect 210418 151784 210424 151796
rect 210476 151784 210482 151836
rect 509050 151784 509056 151836
rect 509108 151824 509114 151836
rect 510890 151824 510896 151836
rect 509108 151796 510896 151824
rect 509108 151784 509114 151796
rect 510890 151784 510896 151796
rect 510948 151784 510954 151836
rect 516042 151784 516048 151836
rect 516100 151824 516106 151836
rect 520182 151824 520188 151836
rect 516100 151796 520188 151824
rect 516100 151784 516106 151796
rect 520182 151784 520188 151796
rect 520240 151784 520246 151836
rect 132402 151716 132408 151768
rect 132460 151756 132466 151768
rect 219342 151756 219348 151768
rect 132460 151728 219348 151756
rect 132460 151716 132466 151728
rect 219342 151716 219348 151728
rect 219400 151716 219406 151768
rect 122742 151648 122748 151700
rect 122800 151688 122806 151700
rect 211614 151688 211620 151700
rect 122800 151660 211620 151688
rect 122800 151648 122806 151660
rect 211614 151648 211620 151660
rect 211672 151648 211678 151700
rect 111702 151580 111708 151632
rect 111760 151620 111766 151632
rect 203978 151620 203984 151632
rect 111760 151592 203984 151620
rect 111760 151580 111766 151592
rect 203978 151580 203984 151592
rect 204036 151580 204042 151632
rect 104802 151512 104808 151564
rect 104860 151552 104866 151564
rect 198826 151552 198832 151564
rect 104860 151524 198832 151552
rect 104860 151512 104866 151524
rect 198826 151512 198832 151524
rect 198884 151512 198890 151564
rect 212442 151512 212448 151564
rect 212500 151552 212506 151564
rect 280982 151552 280988 151564
rect 212500 151524 280988 151552
rect 212500 151512 212506 151524
rect 280982 151512 280988 151524
rect 281040 151512 281046 151564
rect 97902 151444 97908 151496
rect 97960 151484 97966 151496
rect 193674 151484 193680 151496
rect 97960 151456 193680 151484
rect 97960 151444 97966 151456
rect 193674 151444 193680 151456
rect 193732 151444 193738 151496
rect 202782 151444 202788 151496
rect 202840 151484 202846 151496
rect 273254 151484 273260 151496
rect 202840 151456 273260 151484
rect 202840 151444 202846 151456
rect 273254 151444 273260 151456
rect 273312 151444 273318 151496
rect 92382 151376 92388 151428
rect 92440 151416 92446 151428
rect 188522 151416 188528 151428
rect 92440 151388 188528 151416
rect 92440 151376 92446 151388
rect 188522 151376 188528 151388
rect 188580 151376 188586 151428
rect 195882 151376 195888 151428
rect 195940 151416 195946 151428
rect 268194 151416 268200 151428
rect 195940 151388 268200 151416
rect 195940 151376 195946 151388
rect 268194 151376 268200 151388
rect 268252 151376 268258 151428
rect 78582 151308 78588 151360
rect 78640 151348 78646 151360
rect 178310 151348 178316 151360
rect 78640 151320 178316 151348
rect 78640 151308 78646 151320
rect 178310 151308 178316 151320
rect 178368 151308 178374 151360
rect 180702 151308 180708 151360
rect 180760 151348 180766 151360
rect 256602 151348 256608 151360
rect 180760 151320 256608 151348
rect 180760 151308 180766 151320
rect 256602 151308 256608 151320
rect 256660 151308 256666 151360
rect 64782 151240 64788 151292
rect 64840 151280 64846 151292
rect 64840 151252 167592 151280
rect 64840 151240 64846 151252
rect 57882 151172 57888 151224
rect 57940 151212 57946 151224
rect 162854 151212 162860 151224
rect 57940 151184 162860 151212
rect 57940 151172 57946 151184
rect 162854 151172 162860 151184
rect 162912 151172 162918 151224
rect 167564 151212 167592 151252
rect 167638 151240 167644 151292
rect 167696 151280 167702 151292
rect 245010 151280 245016 151292
rect 167696 151252 245016 151280
rect 167696 151240 167702 151252
rect 245010 151240 245016 151252
rect 245068 151240 245074 151292
rect 168006 151212 168012 151224
rect 167564 151184 168012 151212
rect 168006 151172 168012 151184
rect 168064 151172 168070 151224
rect 168098 151172 168104 151224
rect 168156 151212 168162 151224
rect 246298 151212 246304 151224
rect 168156 151184 246304 151212
rect 168156 151172 168162 151184
rect 246298 151172 246304 151184
rect 246356 151172 246362 151224
rect 50982 151104 50988 151156
rect 51040 151144 51046 151156
rect 157702 151144 157708 151156
rect 51040 151116 157708 151144
rect 51040 151104 51046 151116
rect 157702 151104 157708 151116
rect 157760 151104 157766 151156
rect 158622 151104 158628 151156
rect 158680 151144 158686 151156
rect 239950 151144 239956 151156
rect 158680 151116 239956 151144
rect 158680 151104 158686 151116
rect 239950 151104 239956 151116
rect 240008 151104 240014 151156
rect 38562 151036 38568 151088
rect 38620 151076 38626 151088
rect 147490 151076 147496 151088
rect 38620 151048 147496 151076
rect 38620 151036 38626 151048
rect 147490 151036 147496 151048
rect 147548 151036 147554 151088
rect 151722 151036 151728 151088
rect 151780 151076 151786 151088
rect 234798 151076 234804 151088
rect 151780 151048 234804 151076
rect 151780 151036 151786 151048
rect 234798 151036 234804 151048
rect 234856 151036 234862 151088
rect 146202 150968 146208 151020
rect 146260 151008 146266 151020
rect 229646 151008 229652 151020
rect 146260 150980 229652 151008
rect 146260 150968 146266 150980
rect 229646 150968 229652 150980
rect 229704 150968 229710 151020
rect 153102 150900 153108 150952
rect 153160 150940 153166 150952
rect 235442 150940 235448 150952
rect 153160 150912 235448 150940
rect 153160 150900 153166 150912
rect 235442 150900 235448 150912
rect 235500 150900 235506 150952
rect 166902 150832 166908 150884
rect 166960 150872 166966 150884
rect 168098 150872 168104 150884
rect 166960 150844 168104 150872
rect 166960 150832 166966 150844
rect 168098 150832 168104 150844
rect 168156 150832 168162 150884
rect 105814 150628 105820 150680
rect 105872 150668 105878 150680
rect 116026 150668 116032 150680
rect 105872 150640 116032 150668
rect 105872 150628 105878 150640
rect 116026 150628 116032 150640
rect 116084 150628 116090 150680
rect 98914 150560 98920 150612
rect 98972 150600 98978 150612
rect 114462 150600 114468 150612
rect 98972 150572 114468 150600
rect 98972 150560 98978 150572
rect 114462 150560 114468 150572
rect 114520 150560 114526 150612
rect 92014 150492 92020 150544
rect 92072 150532 92078 150544
rect 114002 150532 114008 150544
rect 92072 150504 114008 150532
rect 92072 150492 92078 150504
rect 114002 150492 114008 150504
rect 114060 150492 114066 150544
rect 85206 150424 85212 150476
rect 85264 150464 85270 150476
rect 117038 150464 117044 150476
rect 85264 150436 117044 150464
rect 85264 150424 85270 150436
rect 117038 150424 117044 150436
rect 117096 150424 117102 150476
rect 127066 150152 127072 150204
rect 127124 150192 127130 150204
rect 128216 150192 128222 150204
rect 127124 150164 128222 150192
rect 127124 150152 127130 150164
rect 128216 150152 128222 150164
rect 128274 150152 128280 150204
rect 132494 150152 132500 150204
rect 132552 150192 132558 150204
rect 133368 150192 133374 150204
rect 132552 150164 133374 150192
rect 132552 150152 132558 150164
rect 133368 150152 133374 150164
rect 133426 150152 133432 150204
rect 139394 150152 139400 150204
rect 139452 150192 139458 150204
rect 140452 150192 140458 150204
rect 139452 150164 140458 150192
rect 139452 150152 139458 150164
rect 140452 150152 140458 150164
rect 140510 150152 140516 150204
rect 145098 150152 145104 150204
rect 145156 150192 145162 150204
rect 146248 150192 146254 150204
rect 145156 150164 146254 150192
rect 145156 150152 145162 150164
rect 146248 150152 146254 150164
rect 146306 150152 146312 150204
rect 147674 150152 147680 150204
rect 147732 150192 147738 150204
rect 148824 150192 148830 150204
rect 147732 150164 148830 150192
rect 147732 150152 147738 150164
rect 148824 150152 148830 150164
rect 148882 150152 148888 150204
rect 149146 150152 149152 150204
rect 149204 150192 149210 150204
rect 150020 150192 150026 150204
rect 149204 150164 150026 150192
rect 149204 150152 149210 150164
rect 150020 150152 150026 150164
rect 150078 150152 150084 150204
rect 150526 150152 150532 150204
rect 150584 150192 150590 150204
rect 151308 150192 151314 150204
rect 150584 150164 151314 150192
rect 150584 150152 150590 150164
rect 151308 150152 151314 150164
rect 151366 150152 151372 150204
rect 154666 150152 154672 150204
rect 154724 150192 154730 150204
rect 155816 150192 155822 150204
rect 154724 150164 155822 150192
rect 154724 150152 154730 150164
rect 155816 150152 155822 150164
rect 155874 150152 155880 150204
rect 161474 150152 161480 150204
rect 161532 150192 161538 150204
rect 162256 150192 162262 150204
rect 161532 150164 162262 150192
rect 161532 150152 161538 150164
rect 162256 150152 162262 150164
rect 162314 150152 162320 150204
rect 163038 150152 163044 150204
rect 163096 150192 163102 150204
rect 164188 150192 164194 150204
rect 163096 150164 164194 150192
rect 163096 150152 163102 150164
rect 164188 150152 164194 150164
rect 164246 150152 164252 150204
rect 168374 150152 168380 150204
rect 168432 150192 168438 150204
rect 169340 150192 169346 150204
rect 168432 150164 169346 150192
rect 168432 150152 168438 150164
rect 169340 150152 169346 150164
rect 169398 150152 169404 150204
rect 169846 150152 169852 150204
rect 169904 150192 169910 150204
rect 170628 150192 170634 150204
rect 169904 150164 170634 150192
rect 169904 150152 169910 150164
rect 170628 150152 170634 150164
rect 170686 150152 170692 150204
rect 171134 150152 171140 150204
rect 171192 150192 171198 150204
rect 171916 150192 171922 150204
rect 171192 150164 171922 150192
rect 171192 150152 171198 150164
rect 171916 150152 171922 150164
rect 171974 150152 171980 150204
rect 172698 150152 172704 150204
rect 172756 150192 172762 150204
rect 173848 150192 173854 150204
rect 172756 150164 173854 150192
rect 172756 150152 172762 150164
rect 173848 150152 173854 150164
rect 173906 150152 173912 150204
rect 179414 150152 179420 150204
rect 179472 150192 179478 150204
rect 180288 150192 180294 150204
rect 179472 150164 180294 150192
rect 179472 150152 179478 150164
rect 180288 150152 180294 150164
rect 180346 150152 180352 150204
rect 180978 150152 180984 150204
rect 181036 150192 181042 150204
rect 182128 150192 182134 150204
rect 181036 150164 182134 150192
rect 181036 150152 181042 150164
rect 182128 150152 182134 150164
rect 182186 150152 182192 150204
rect 183554 150152 183560 150204
rect 183612 150192 183618 150204
rect 184704 150192 184710 150204
rect 183612 150164 184710 150192
rect 183612 150152 183618 150164
rect 184704 150152 184710 150164
rect 184762 150152 184768 150204
rect 190730 150152 190736 150204
rect 190788 150192 190794 150204
rect 191788 150192 191794 150204
rect 190788 150164 191794 150192
rect 190788 150152 190794 150164
rect 191788 150152 191794 150164
rect 191846 150152 191852 150204
rect 194594 150152 194600 150204
rect 194652 150192 194658 150204
rect 195652 150192 195658 150204
rect 194652 150164 195658 150192
rect 194652 150152 194658 150164
rect 195652 150152 195658 150164
rect 195710 150152 195716 150204
rect 200298 150152 200304 150204
rect 200356 150192 200362 150204
rect 201448 150192 201454 150204
rect 200356 150164 201454 150192
rect 200356 150152 200362 150164
rect 201448 150152 201454 150164
rect 201506 150152 201512 150204
rect 209958 150152 209964 150204
rect 210016 150192 210022 150204
rect 211108 150192 211114 150204
rect 210016 150164 211114 150192
rect 210016 150152 210022 150164
rect 211108 150152 211114 150164
rect 211166 150152 211172 150204
rect 224954 150152 224960 150204
rect 225012 150192 225018 150204
rect 225828 150192 225834 150204
rect 225012 150164 225834 150192
rect 225012 150152 225018 150164
rect 225828 150152 225834 150164
rect 225886 150152 225892 150204
rect 229186 150152 229192 150204
rect 229244 150192 229250 150204
rect 230336 150192 230342 150204
rect 229244 150164 230342 150192
rect 229244 150152 229250 150164
rect 230336 150152 230342 150164
rect 230394 150152 230400 150204
rect 233234 150152 233240 150204
rect 233292 150192 233298 150204
rect 234200 150192 234206 150204
rect 233292 150164 234206 150192
rect 233292 150152 233298 150164
rect 234200 150152 234206 150164
rect 234258 150152 234264 150204
rect 240134 150152 240140 150204
rect 240192 150192 240198 150204
rect 241284 150192 241290 150204
rect 240192 150164 241290 150192
rect 240192 150152 240198 150164
rect 241284 150152 241290 150164
rect 241342 150152 241348 150204
rect 242894 150152 242900 150204
rect 242952 150192 242958 150204
rect 243768 150192 243774 150204
rect 242952 150164 243774 150192
rect 242952 150152 242958 150164
rect 243768 150152 243774 150164
rect 243826 150152 243832 150204
rect 247126 150152 247132 150204
rect 247184 150192 247190 150204
rect 248276 150192 248282 150204
rect 247184 150164 248282 150192
rect 247184 150152 247190 150164
rect 248276 150152 248282 150164
rect 248334 150152 248340 150204
rect 252554 150152 252560 150204
rect 252612 150192 252618 150204
rect 253428 150192 253434 150204
rect 252612 150164 253434 150192
rect 252612 150152 252618 150164
rect 253428 150152 253434 150164
rect 253486 150152 253492 150204
rect 258074 150152 258080 150204
rect 258132 150192 258138 150204
rect 259224 150192 259230 150204
rect 258132 150164 259230 150192
rect 258132 150152 258138 150164
rect 259224 150152 259230 150164
rect 259282 150152 259288 150204
rect 260834 150152 260840 150204
rect 260892 150192 260898 150204
rect 261800 150192 261806 150204
rect 260892 150164 261806 150192
rect 260892 150152 260898 150164
rect 261800 150152 261806 150164
rect 261858 150152 261864 150204
rect 263594 150152 263600 150204
rect 263652 150192 263658 150204
rect 264376 150192 264382 150204
rect 263652 150164 264382 150192
rect 263652 150152 263658 150164
rect 264376 150152 264382 150164
rect 264434 150152 264440 150204
rect 265158 150152 265164 150204
rect 265216 150192 265222 150204
rect 266308 150192 266314 150204
rect 265216 150164 266314 150192
rect 265216 150152 265222 150164
rect 266308 150152 266314 150164
rect 266366 150152 266372 150204
rect 273438 150152 273444 150204
rect 273496 150192 273502 150204
rect 274588 150192 274594 150204
rect 273496 150164 274594 150192
rect 273496 150152 273502 150164
rect 274588 150152 274594 150164
rect 274646 150152 274652 150204
rect 276014 150152 276020 150204
rect 276072 150192 276078 150204
rect 277164 150192 277170 150204
rect 276072 150164 277170 150192
rect 276072 150152 276078 150164
rect 277164 150152 277170 150164
rect 277222 150152 277228 150204
rect 283098 150152 283104 150204
rect 283156 150192 283162 150204
rect 284248 150192 284254 150204
rect 283156 150164 284254 150192
rect 283156 150152 283162 150164
rect 284248 150152 284254 150164
rect 284306 150152 284312 150204
rect 291194 150152 291200 150204
rect 291252 150192 291258 150204
rect 291976 150192 291982 150204
rect 291252 150164 291982 150192
rect 291252 150152 291258 150164
rect 291976 150152 291982 150164
rect 292034 150152 292040 150204
rect 292758 150152 292764 150204
rect 292816 150192 292822 150204
rect 293908 150192 293914 150204
rect 292816 150164 293914 150192
rect 292816 150152 292822 150164
rect 293908 150152 293914 150164
rect 293966 150152 293972 150204
rect 299474 150152 299480 150204
rect 299532 150192 299538 150204
rect 300348 150192 300354 150204
rect 299532 150164 300354 150192
rect 299532 150152 299538 150164
rect 300348 150152 300354 150164
rect 300406 150152 300412 150204
rect 310606 150152 310612 150204
rect 310664 150192 310670 150204
rect 311848 150192 311854 150204
rect 310664 150164 311854 150192
rect 310664 150152 310670 150164
rect 311848 150152 311854 150164
rect 311906 150152 311912 150204
rect 311986 150152 311992 150204
rect 312044 150192 312050 150204
rect 313136 150192 313142 150204
rect 312044 150164 313142 150192
rect 312044 150152 312050 150164
rect 313136 150152 313142 150164
rect 313194 150152 313200 150204
rect 330018 150152 330024 150204
rect 330076 150192 330082 150204
rect 331168 150192 331174 150204
rect 330076 150164 331174 150192
rect 330076 150152 330082 150164
rect 331168 150152 331174 150164
rect 331226 150152 331232 150204
rect 331306 150152 331312 150204
rect 331364 150192 331370 150204
rect 332456 150192 332462 150204
rect 331364 150164 332462 150192
rect 331364 150152 331370 150164
rect 332456 150152 332462 150164
rect 332514 150152 332520 150204
rect 339586 150152 339592 150204
rect 339644 150192 339650 150204
rect 340736 150192 340742 150204
rect 339644 150164 340742 150192
rect 339644 150152 339650 150164
rect 340736 150152 340742 150164
rect 340794 150152 340800 150204
rect 349246 150152 349252 150204
rect 349304 150192 349310 150204
rect 350396 150192 350402 150204
rect 349304 150164 350402 150192
rect 349304 150152 349310 150164
rect 350396 150152 350402 150164
rect 350454 150152 350460 150204
rect 350534 150152 350540 150204
rect 350592 150192 350598 150204
rect 351684 150192 351690 150204
rect 350592 150164 351690 150192
rect 350592 150152 350598 150164
rect 351684 150152 351690 150164
rect 351742 150152 351748 150204
rect 351914 150152 351920 150204
rect 351972 150192 351978 150204
rect 352972 150192 352978 150204
rect 351972 150164 352978 150192
rect 351972 150152 351978 150164
rect 352972 150152 352978 150164
rect 353030 150152 353036 150204
rect 357618 150152 357624 150204
rect 357676 150192 357682 150204
rect 358768 150192 358774 150204
rect 357676 150164 358774 150192
rect 357676 150152 357682 150164
rect 358768 150152 358774 150164
rect 358826 150152 358832 150204
rect 360194 150152 360200 150204
rect 360252 150192 360258 150204
rect 361344 150192 361350 150204
rect 360252 150164 361350 150192
rect 360252 150152 360258 150164
rect 361344 150152 361350 150164
rect 361402 150152 361408 150204
rect 361574 150152 361580 150204
rect 361632 150192 361638 150204
rect 362632 150192 362638 150204
rect 361632 150164 362638 150192
rect 361632 150152 361638 150164
rect 362632 150152 362638 150164
rect 362690 150152 362696 150204
rect 365898 150152 365904 150204
rect 365956 150192 365962 150204
rect 367048 150192 367054 150204
rect 365956 150164 367054 150192
rect 365956 150152 365962 150164
rect 367048 150152 367054 150164
rect 367106 150152 367112 150204
rect 383654 150152 383660 150204
rect 383712 150192 383718 150204
rect 384436 150192 384442 150204
rect 383712 150164 384442 150192
rect 383712 150152 383718 150164
rect 384436 150152 384442 150164
rect 384494 150152 384500 150204
rect 385218 150152 385224 150204
rect 385276 150192 385282 150204
rect 386368 150192 386374 150204
rect 385276 150164 386374 150192
rect 385276 150152 385282 150164
rect 386368 150152 386374 150164
rect 386426 150152 386432 150204
rect 386506 150152 386512 150204
rect 386564 150192 386570 150204
rect 387656 150192 387662 150204
rect 386564 150164 387662 150192
rect 386564 150152 386570 150164
rect 387656 150152 387662 150164
rect 387714 150152 387720 150204
rect 391934 150152 391940 150204
rect 391992 150192 391998 150204
rect 392808 150192 392814 150204
rect 391992 150164 392814 150192
rect 391992 150152 391998 150164
rect 392808 150152 392814 150164
rect 392866 150152 392872 150204
rect 396166 150152 396172 150204
rect 396224 150192 396230 150204
rect 397224 150192 397230 150204
rect 396224 150164 397230 150192
rect 396224 150152 396230 150164
rect 397224 150152 397230 150164
rect 397282 150152 397288 150204
rect 400214 150152 400220 150204
rect 400272 150192 400278 150204
rect 401088 150192 401094 150204
rect 400272 150164 401094 150192
rect 400272 150152 400278 150164
rect 401088 150152 401094 150164
rect 401146 150152 401152 150204
rect 412818 150152 412824 150204
rect 412876 150192 412882 150204
rect 413968 150192 413974 150204
rect 412876 150164 413974 150192
rect 412876 150152 412882 150164
rect 413968 150152 413974 150164
rect 414026 150152 414032 150204
rect 423766 150152 423772 150204
rect 423824 150192 423830 150204
rect 424916 150192 424922 150204
rect 423824 150164 424922 150192
rect 423824 150152 423830 150164
rect 424916 150152 424922 150164
rect 424974 150152 424980 150204
rect 434714 150152 434720 150204
rect 434772 150192 434778 150204
rect 435772 150192 435778 150204
rect 434772 150164 435778 150192
rect 434772 150152 434778 150164
rect 435772 150152 435778 150164
rect 435830 150152 435836 150204
rect 441706 150152 441712 150204
rect 441764 150192 441770 150204
rect 442856 150192 442862 150204
rect 441764 150164 442862 150192
rect 441764 150152 441770 150164
rect 442856 150152 442862 150164
rect 442914 150152 442920 150204
rect 442994 150152 443000 150204
rect 443052 150192 443058 150204
rect 444144 150192 444150 150204
rect 443052 150164 444150 150192
rect 443052 150152 443058 150164
rect 444144 150152 444150 150164
rect 444202 150152 444208 150204
rect 444374 150152 444380 150204
rect 444432 150192 444438 150204
rect 445432 150192 445438 150204
rect 444432 150164 445438 150192
rect 444432 150152 444438 150164
rect 445432 150152 445438 150164
rect 445490 150152 445496 150204
rect 456794 150152 456800 150204
rect 456852 150192 456858 150204
rect 457668 150192 457674 150204
rect 456852 150164 457674 150192
rect 456852 150152 456858 150164
rect 457668 150152 457674 150164
rect 457726 150152 457732 150204
rect 477678 150152 477684 150204
rect 477736 150192 477742 150204
rect 478828 150192 478834 150204
rect 477736 150164 478834 150192
rect 477736 150152 477742 150164
rect 478828 150152 478834 150164
rect 478886 150152 478892 150204
rect 478966 150152 478972 150204
rect 479024 150192 479030 150204
rect 480116 150192 480122 150204
rect 479024 150164 480122 150192
rect 479024 150152 479030 150164
rect 480116 150152 480122 150164
rect 480174 150152 480180 150204
rect 483014 150152 483020 150204
rect 483072 150192 483078 150204
rect 483980 150192 483986 150204
rect 483072 150164 483986 150192
rect 483072 150152 483078 150164
rect 483980 150152 483986 150164
rect 484038 150152 484044 150204
rect 485774 150152 485780 150204
rect 485832 150192 485838 150204
rect 486556 150192 486562 150204
rect 485832 150164 486562 150192
rect 485832 150152 485838 150164
rect 486556 150152 486562 150164
rect 486614 150152 486620 150204
rect 488626 150152 488632 150204
rect 488684 150192 488690 150204
rect 489684 150192 489690 150204
rect 488684 150164 489690 150192
rect 488684 150152 488690 150164
rect 489684 150152 489690 150164
rect 489742 150152 489748 150204
rect 489914 150152 489920 150204
rect 489972 150192 489978 150204
rect 490972 150192 490978 150204
rect 489972 150164 490978 150192
rect 489972 150152 489978 150164
rect 490972 150152 490978 150164
rect 491030 150152 491036 150204
rect 491294 150152 491300 150204
rect 491352 150192 491358 150204
rect 492260 150192 492266 150204
rect 491352 150164 492266 150192
rect 491352 150152 491358 150164
rect 492260 150152 492266 150164
rect 492318 150152 492324 150204
rect 97718 149880 97724 149932
rect 97776 149920 97782 149932
rect 116486 149920 116492 149932
rect 97776 149892 116492 149920
rect 97776 149880 97782 149892
rect 116486 149880 116492 149892
rect 116544 149880 116550 149932
rect 89162 149812 89168 149864
rect 89220 149852 89226 149864
rect 116210 149852 116216 149864
rect 89220 149824 116216 149852
rect 89220 149812 89226 149824
rect 116210 149812 116216 149824
rect 116268 149812 116274 149864
rect 82814 149744 82820 149796
rect 82872 149784 82878 149796
rect 117130 149784 117136 149796
rect 82872 149756 117136 149784
rect 82872 149744 82878 149756
rect 117130 149744 117136 149756
rect 117188 149744 117194 149796
rect 78582 149676 78588 149728
rect 78640 149716 78646 149728
rect 112806 149716 112812 149728
rect 78640 149688 112812 149716
rect 78640 149676 78646 149688
rect 112806 149676 112812 149688
rect 112864 149676 112870 149728
rect 75178 149608 75184 149660
rect 75236 149648 75242 149660
rect 114186 149648 114192 149660
rect 75236 149620 114192 149648
rect 75236 149608 75242 149620
rect 114186 149608 114192 149620
rect 114244 149608 114250 149660
rect 68370 149540 68376 149592
rect 68428 149580 68434 149592
rect 112714 149580 112720 149592
rect 68428 149552 112720 149580
rect 68428 149540 68434 149552
rect 112714 149540 112720 149552
rect 112772 149540 112778 149592
rect 64690 149472 64696 149524
rect 64748 149512 64754 149524
rect 111242 149512 111248 149524
rect 64748 149484 111248 149512
rect 64748 149472 64754 149484
rect 111242 149472 111248 149484
rect 111300 149472 111306 149524
rect 61378 149404 61384 149456
rect 61436 149444 61442 149456
rect 112622 149444 112628 149456
rect 61436 149416 112628 149444
rect 61436 149404 61442 149416
rect 112622 149404 112628 149416
rect 112680 149404 112686 149456
rect 57882 149336 57888 149388
rect 57940 149376 57946 149388
rect 112530 149376 112536 149388
rect 57940 149348 112536 149376
rect 57940 149336 57946 149348
rect 112530 149336 112536 149348
rect 112588 149336 112594 149388
rect 40770 149268 40776 149320
rect 40828 149268 40834 149320
rect 44082 149268 44088 149320
rect 44140 149308 44146 149320
rect 44140 149280 45554 149308
rect 44140 149268 44146 149280
rect 40788 149104 40816 149268
rect 45526 149172 45554 149280
rect 47578 149268 47584 149320
rect 47636 149268 47642 149320
rect 50982 149268 50988 149320
rect 51040 149308 51046 149320
rect 112438 149308 112444 149320
rect 51040 149280 112444 149308
rect 51040 149268 51046 149280
rect 112438 149268 112444 149280
rect 112496 149268 112502 149320
rect 47596 149240 47624 149268
rect 111150 149240 111156 149252
rect 47596 149212 111156 149240
rect 111150 149200 111156 149212
rect 111208 149200 111214 149252
rect 111058 149172 111064 149184
rect 45526 149144 111064 149172
rect 111058 149132 111064 149144
rect 111116 149132 111122 149184
rect 109678 149104 109684 149116
rect 40788 149076 109684 149104
rect 109678 149064 109684 149076
rect 109736 149064 109742 149116
rect 109586 148996 109592 149048
rect 109644 149036 109650 149048
rect 116118 149036 116124 149048
rect 109644 149008 116124 149036
rect 109644 148996 109650 149008
rect 116118 148996 116124 149008
rect 116176 148996 116182 149048
rect 110322 147024 110328 147076
rect 110380 147064 110386 147076
rect 116118 147064 116124 147076
rect 110380 147036 116124 147064
rect 110380 147024 110386 147036
rect 116118 147024 116124 147036
rect 116176 147024 116182 147076
rect 110046 146956 110052 147008
rect 110104 146996 110110 147008
rect 116854 146996 116860 147008
rect 110104 146968 116860 146996
rect 110104 146956 110110 146968
rect 116854 146956 116860 146968
rect 116912 146956 116918 147008
rect 110230 146888 110236 146940
rect 110288 146928 110294 146940
rect 116946 146928 116952 146940
rect 110288 146900 116952 146928
rect 110288 146888 110294 146900
rect 116946 146888 116952 146900
rect 117004 146888 117010 146940
rect 110138 145528 110144 145580
rect 110196 145568 110202 145580
rect 116394 145568 116400 145580
rect 110196 145540 116400 145568
rect 110196 145528 110202 145540
rect 116394 145528 116400 145540
rect 116452 145528 116458 145580
rect 113726 143556 113732 143608
rect 113784 143596 113790 143608
rect 115198 143596 115204 143608
rect 113784 143568 115204 143596
rect 113784 143556 113790 143568
rect 115198 143556 115204 143568
rect 115256 143556 115262 143608
rect 114462 143488 114468 143540
rect 114520 143528 114526 143540
rect 115934 143528 115940 143540
rect 114520 143500 115940 143528
rect 114520 143488 114526 143500
rect 115934 143488 115940 143500
rect 115992 143488 115998 143540
rect 114370 141720 114376 141772
rect 114428 141760 114434 141772
rect 115934 141760 115940 141772
rect 114428 141732 115940 141760
rect 114428 141720 114434 141732
rect 115934 141720 115940 141732
rect 115992 141720 115998 141772
rect 114002 140700 114008 140752
rect 114060 140740 114066 140752
rect 115934 140740 115940 140752
rect 114060 140712 115940 140740
rect 114060 140700 114066 140712
rect 115934 140700 115940 140712
rect 115992 140700 115998 140752
rect 109770 134512 109776 134564
rect 109828 134552 109834 134564
rect 117038 134552 117044 134564
rect 109828 134524 117044 134552
rect 109828 134512 109834 134524
rect 117038 134512 117044 134524
rect 117096 134512 117102 134564
rect 112806 132404 112812 132456
rect 112864 132444 112870 132456
rect 116118 132444 116124 132456
rect 112864 132416 116124 132444
rect 112864 132404 112870 132416
rect 116118 132404 116124 132416
rect 116176 132404 116182 132456
rect 114186 131044 114192 131096
rect 114244 131084 114250 131096
rect 115934 131084 115940 131096
rect 114244 131056 115940 131084
rect 114244 131044 114250 131056
rect 115934 131044 115940 131056
rect 115992 131044 115998 131096
rect 112714 126896 112720 126948
rect 112772 126936 112778 126948
rect 116118 126936 116124 126948
rect 112772 126908 116124 126936
rect 112772 126896 112778 126908
rect 116118 126896 116124 126908
rect 116176 126896 116182 126948
rect 111242 124108 111248 124160
rect 111300 124148 111306 124160
rect 116118 124148 116124 124160
rect 111300 124120 116124 124148
rect 111300 124108 111306 124120
rect 116118 124108 116124 124120
rect 116176 124108 116182 124160
rect 112622 122748 112628 122800
rect 112680 122788 112686 122800
rect 115934 122788 115940 122800
rect 112680 122760 115940 122788
rect 112680 122748 112686 122760
rect 115934 122748 115940 122760
rect 115992 122748 115998 122800
rect 112530 121388 112536 121440
rect 112588 121428 112594 121440
rect 115934 121428 115940 121440
rect 112588 121400 115940 121428
rect 112588 121388 112594 121400
rect 115934 121388 115940 121400
rect 115992 121388 115998 121440
rect 114186 118804 114192 118856
rect 114244 118844 114250 118856
rect 115290 118844 115296 118856
rect 114244 118816 115296 118844
rect 114244 118804 114250 118816
rect 115290 118804 115296 118816
rect 115348 118804 115354 118856
rect 112438 117240 112444 117292
rect 112496 117280 112502 117292
rect 116026 117280 116032 117292
rect 112496 117252 116032 117280
rect 112496 117240 112502 117252
rect 116026 117240 116032 117252
rect 116084 117240 116090 117292
rect 111150 114452 111156 114504
rect 111208 114492 111214 114504
rect 116118 114492 116124 114504
rect 111208 114464 116124 114492
rect 111208 114452 111214 114464
rect 116118 114452 116124 114464
rect 116176 114452 116182 114504
rect 111058 113092 111064 113144
rect 111116 113132 111122 113144
rect 116118 113132 116124 113144
rect 111116 113104 116124 113132
rect 111116 113092 111122 113104
rect 116118 113092 116124 113104
rect 116176 113092 116182 113144
rect 109678 111732 109684 111784
rect 109736 111772 109742 111784
rect 116118 111772 116124 111784
rect 109736 111744 116124 111772
rect 109736 111732 109742 111744
rect 116118 111732 116124 111744
rect 116176 111732 116182 111784
rect 113542 109556 113548 109608
rect 113600 109596 113606 109608
rect 115382 109596 115388 109608
rect 113600 109568 115388 109596
rect 113600 109556 113606 109568
rect 115382 109556 115388 109568
rect 115440 109556 115446 109608
rect 114278 108944 114284 108996
rect 114336 108984 114342 108996
rect 116394 108984 116400 108996
rect 114336 108956 116400 108984
rect 114336 108944 114342 108956
rect 116394 108944 116400 108956
rect 116452 108944 116458 108996
rect 114094 104796 114100 104848
rect 114152 104836 114158 104848
rect 115934 104836 115940 104848
rect 114152 104808 115940 104836
rect 114152 104796 114158 104808
rect 115934 104796 115940 104808
rect 115992 104796 115998 104848
rect 114462 96840 114468 96892
rect 114520 96880 114526 96892
rect 116762 96880 116768 96892
rect 114520 96852 116768 96880
rect 114520 96840 114526 96852
rect 116762 96840 116768 96852
rect 116820 96840 116826 96892
rect 113818 93576 113824 93628
rect 113876 93616 113882 93628
rect 116486 93616 116492 93628
rect 113876 93588 116492 93616
rect 113876 93576 113882 93588
rect 116486 93576 116492 93588
rect 116544 93576 116550 93628
rect 113910 92420 113916 92472
rect 113968 92460 113974 92472
rect 116118 92460 116124 92472
rect 113968 92432 116124 92460
rect 113968 92420 113974 92432
rect 116118 92420 116124 92432
rect 116176 92420 116182 92472
rect 115198 91604 115204 91656
rect 115256 91644 115262 91656
rect 116854 91644 116860 91656
rect 115256 91616 116860 91644
rect 115256 91604 115262 91616
rect 116854 91604 116860 91616
rect 116912 91604 116918 91656
rect 114462 87184 114468 87236
rect 114520 87224 114526 87236
rect 116670 87224 116676 87236
rect 114520 87196 116676 87224
rect 114520 87184 114526 87196
rect 116670 87184 116676 87196
rect 116728 87184 116734 87236
rect 114002 86912 114008 86964
rect 114060 86952 114066 86964
rect 116210 86952 116216 86964
rect 114060 86924 116216 86952
rect 114060 86912 114066 86924
rect 116210 86912 116216 86924
rect 116268 86912 116274 86964
rect 113818 71748 113824 71800
rect 113876 71788 113882 71800
rect 116394 71788 116400 71800
rect 113876 71760 116400 71788
rect 113876 71748 113882 71760
rect 116394 71748 116400 71760
rect 116452 71748 116458 71800
rect 114094 69028 114100 69080
rect 114152 69068 114158 69080
rect 116302 69068 116308 69080
rect 114152 69040 116308 69068
rect 114152 69028 114158 69040
rect 116302 69028 116308 69040
rect 116360 69028 116366 69080
rect 114186 67600 114192 67652
rect 114244 67640 114250 67652
rect 116210 67640 116216 67652
rect 114244 67612 116216 67640
rect 114244 67600 114250 67612
rect 116210 67600 116216 67612
rect 116268 67600 116274 67652
rect 114462 64676 114468 64728
rect 114520 64716 114526 64728
rect 116578 64716 116584 64728
rect 114520 64688 116584 64716
rect 114520 64676 114526 64688
rect 116578 64676 116584 64688
rect 116636 64676 116642 64728
rect 112438 62092 112444 62144
rect 112496 62132 112502 62144
rect 116118 62132 116124 62144
rect 112496 62104 116124 62132
rect 112496 62092 112502 62104
rect 116118 62092 116124 62104
rect 116176 62092 116182 62144
rect 111058 59372 111064 59424
rect 111116 59412 111122 59424
rect 116118 59412 116124 59424
rect 111116 59384 116124 59412
rect 111116 59372 111122 59384
rect 116118 59372 116124 59384
rect 116176 59372 116182 59424
rect 113818 51076 113824 51128
rect 113876 51116 113882 51128
rect 115934 51116 115940 51128
rect 113876 51088 115940 51116
rect 113876 51076 113882 51088
rect 115934 51076 115940 51088
rect 115992 51076 115998 51128
rect 114278 48220 114284 48272
rect 114336 48260 114342 48272
rect 116854 48260 116860 48272
rect 114336 48232 116860 48260
rect 114336 48220 114342 48232
rect 116854 48220 116860 48232
rect 116912 48220 116918 48272
rect 113910 46928 113916 46980
rect 113968 46968 113974 46980
rect 116026 46968 116032 46980
rect 113968 46940 116032 46968
rect 113968 46928 113974 46940
rect 116026 46928 116032 46940
rect 116084 46928 116090 46980
rect 114002 42780 114008 42832
rect 114060 42820 114066 42832
rect 116394 42820 116400 42832
rect 114060 42792 116400 42820
rect 114060 42780 114066 42792
rect 116394 42780 116400 42792
rect 116452 42780 116458 42832
rect 114094 38632 114100 38684
rect 114152 38672 114158 38684
rect 115934 38672 115940 38684
rect 114152 38644 115940 38672
rect 114152 38632 114158 38644
rect 115934 38632 115940 38644
rect 115992 38632 115998 38684
rect 109678 37272 109684 37324
rect 109736 37312 109742 37324
rect 116118 37312 116124 37324
rect 109736 37284 116124 37312
rect 109736 37272 109742 37284
rect 116118 37272 116124 37284
rect 116176 37272 116182 37324
rect 109770 33124 109776 33176
rect 109828 33164 109834 33176
rect 116118 33164 116124 33176
rect 109828 33136 116124 33164
rect 109828 33124 109834 33136
rect 116118 33124 116124 33136
rect 116176 33124 116182 33176
rect 116302 31016 116308 31068
rect 116360 31056 116366 31068
rect 117222 31056 117228 31068
rect 116360 31028 117228 31056
rect 116360 31016 116366 31028
rect 117222 31016 117228 31028
rect 117280 31016 117286 31068
rect 112530 27616 112536 27668
rect 112588 27656 112594 27668
rect 116118 27656 116124 27668
rect 112588 27628 116124 27656
rect 112588 27616 112594 27628
rect 116118 27616 116124 27628
rect 116176 27616 116182 27668
rect 112622 23468 112628 23520
rect 112680 23508 112686 23520
rect 116118 23508 116124 23520
rect 112680 23480 116124 23508
rect 112680 23468 112686 23480
rect 116118 23468 116124 23480
rect 116176 23468 116182 23520
rect 111242 22788 111248 22840
rect 111300 22828 111306 22840
rect 117038 22828 117044 22840
rect 111300 22800 117044 22828
rect 111300 22788 111306 22800
rect 117038 22788 117044 22800
rect 117096 22788 117102 22840
rect 111150 22720 111156 22772
rect 111208 22760 111214 22772
rect 116302 22760 116308 22772
rect 111208 22732 116308 22760
rect 111208 22720 111214 22732
rect 116302 22720 116308 22732
rect 116360 22720 116366 22772
rect 112714 22108 112720 22160
rect 112772 22148 112778 22160
rect 116118 22148 116124 22160
rect 112772 22120 116124 22148
rect 112772 22108 112778 22120
rect 116118 22108 116124 22120
rect 116176 22108 116182 22160
rect 111334 19320 111340 19372
rect 111392 19360 111398 19372
rect 116118 19360 116124 19372
rect 111392 19332 116124 19360
rect 111392 19320 111398 19332
rect 116118 19320 116124 19332
rect 116176 19320 116182 19372
rect 111426 17960 111432 18012
rect 111484 18000 111490 18012
rect 116118 18000 116124 18012
rect 111484 17972 116124 18000
rect 111484 17960 111490 17972
rect 116118 17960 116124 17972
rect 116176 17960 116182 18012
rect 111610 15172 111616 15224
rect 111668 15212 111674 15224
rect 116118 15212 116124 15224
rect 111668 15184 116124 15212
rect 111668 15172 111674 15184
rect 116118 15172 116124 15184
rect 116176 15172 116182 15224
rect 114278 13812 114284 13864
rect 114336 13852 114342 13864
rect 115934 13852 115940 13864
rect 114336 13824 115940 13852
rect 114336 13812 114342 13824
rect 115934 13812 115940 13824
rect 115992 13812 115998 13864
rect 114186 7964 114192 8016
rect 114244 8004 114250 8016
rect 115198 8004 115204 8016
rect 114244 7976 115204 8004
rect 114244 7964 114250 7976
rect 115198 7964 115204 7976
rect 115256 7964 115262 8016
rect 109862 4836 109868 4888
rect 109920 4876 109926 4888
rect 116946 4876 116952 4888
rect 109920 4848 116952 4876
rect 109920 4836 109926 4848
rect 116946 4836 116952 4848
rect 117004 4836 117010 4888
rect 109954 4768 109960 4820
rect 110012 4808 110018 4820
rect 117222 4808 117228 4820
rect 110012 4780 117228 4808
rect 110012 4768 110018 4780
rect 117222 4768 117228 4780
rect 117280 4768 117286 4820
rect 109586 4496 109592 4548
rect 109644 4536 109650 4548
rect 112438 4536 112444 4548
rect 109644 4508 112444 4536
rect 109644 4496 109650 4508
rect 112438 4496 112444 4508
rect 112496 4496 112502 4548
rect 111518 3040 111524 3052
rect 38626 3012 41414 3040
rect 38626 2972 38654 3012
rect 26206 2944 28994 2972
rect 2498 2796 2504 2848
rect 2556 2836 2562 2848
rect 26206 2836 26234 2944
rect 2556 2808 26234 2836
rect 2556 2796 2562 2808
rect 28966 2564 28994 2944
rect 33244 2944 38654 2972
rect 32766 2592 32772 2644
rect 32824 2632 32830 2644
rect 33244 2632 33272 2944
rect 41386 2904 41414 3012
rect 84166 3012 111524 3040
rect 84166 2904 84194 3012
rect 111518 3000 111524 3012
rect 111576 3000 111582 3052
rect 118694 2972 118700 2984
rect 41386 2876 84194 2904
rect 106108 2944 118700 2972
rect 32824 2604 33272 2632
rect 33796 2808 96614 2836
rect 32824 2592 32830 2604
rect 33796 2564 33824 2808
rect 28966 2536 33824 2564
rect 96586 2564 96614 2808
rect 106108 2768 106136 2944
rect 118694 2932 118700 2944
rect 118752 2932 118758 2984
rect 116118 2836 116124 2848
rect 98288 2740 106136 2768
rect 106246 2808 116124 2836
rect 98288 2644 98316 2740
rect 106246 2700 106274 2808
rect 116118 2796 116124 2808
rect 116176 2796 116182 2848
rect 101600 2672 106274 2700
rect 98270 2592 98276 2644
rect 98328 2592 98334 2644
rect 101600 2564 101628 2672
rect 106182 2592 106188 2644
rect 106240 2632 106246 2644
rect 111058 2632 111064 2644
rect 106240 2604 111064 2632
rect 106240 2592 106246 2604
rect 111058 2592 111064 2604
rect 111116 2592 111122 2644
rect 96586 2536 101628 2564
rect 93026 2116 93032 2168
rect 93084 2156 93090 2168
rect 116670 2156 116676 2168
rect 93084 2128 116676 2156
rect 93084 2116 93090 2128
rect 116670 2116 116676 2128
rect 116728 2116 116734 2168
rect 86402 2048 86408 2100
rect 86460 2088 86466 2100
rect 116762 2088 116768 2100
rect 86460 2060 116768 2088
rect 86460 2048 86466 2060
rect 116762 2048 116768 2060
rect 116820 2048 116826 2100
rect 79594 1980 79600 2032
rect 79652 2020 79658 2032
rect 116854 2020 116860 2032
rect 79652 1992 116860 2020
rect 79652 1980 79658 1992
rect 116854 1980 116860 1992
rect 116912 1980 116918 2032
rect 72694 1912 72700 1964
rect 72752 1952 72758 1964
rect 109862 1952 109868 1964
rect 72752 1924 109868 1952
rect 72752 1912 72758 1924
rect 109862 1912 109868 1924
rect 109920 1912 109926 1964
rect 65978 1844 65984 1896
rect 66036 1884 66042 1896
rect 109678 1884 109684 1896
rect 66036 1856 109684 1884
rect 66036 1844 66042 1856
rect 109678 1844 109684 1856
rect 109736 1844 109742 1896
rect 59354 1776 59360 1828
rect 59412 1816 59418 1828
rect 109770 1816 109776 1828
rect 59412 1788 109776 1816
rect 59412 1776 59418 1788
rect 109770 1776 109776 1788
rect 109828 1776 109834 1828
rect 52638 1708 52644 1760
rect 52696 1748 52702 1760
rect 116486 1748 116492 1760
rect 52696 1720 116492 1748
rect 52696 1708 52702 1720
rect 116486 1708 116492 1720
rect 116544 1708 116550 1760
rect 46014 1640 46020 1692
rect 46072 1680 46078 1692
rect 112530 1680 112536 1692
rect 46072 1652 112536 1680
rect 46072 1640 46078 1652
rect 112530 1640 112536 1652
rect 112588 1640 112594 1692
rect 49326 1572 49332 1624
rect 49384 1612 49390 1624
rect 116394 1612 116400 1624
rect 49384 1584 116400 1612
rect 49384 1572 49390 1584
rect 116394 1572 116400 1584
rect 116452 1572 116458 1624
rect 32674 1504 32680 1556
rect 32732 1544 32738 1556
rect 111334 1544 111340 1556
rect 32732 1516 111340 1544
rect 32732 1504 32738 1516
rect 111334 1504 111340 1516
rect 111392 1504 111398 1556
rect 12618 1436 12624 1488
rect 12676 1476 12682 1488
rect 97994 1476 98000 1488
rect 12676 1448 98000 1476
rect 12676 1436 12682 1448
rect 97994 1436 98000 1448
rect 98052 1436 98058 1488
rect 99374 1436 99380 1488
rect 99432 1476 99438 1488
rect 111150 1476 111156 1488
rect 99432 1448 111156 1476
rect 99432 1436 99438 1448
rect 111150 1436 111156 1448
rect 111208 1436 111214 1488
rect 118694 1436 118700 1488
rect 118752 1476 118758 1488
rect 143626 1476 143632 1488
rect 118752 1448 143632 1476
rect 118752 1436 118758 1448
rect 143626 1436 143632 1448
rect 143684 1436 143690 1488
rect 394234 1436 394240 1488
rect 394292 1476 394298 1488
rect 425790 1476 425796 1488
rect 394292 1448 425796 1476
rect 394292 1436 394298 1448
rect 425790 1436 425796 1448
rect 425848 1436 425854 1488
rect 444282 1436 444288 1488
rect 444340 1476 444346 1488
rect 491294 1476 491300 1488
rect 444340 1448 491300 1476
rect 444340 1436 444346 1448
rect 491294 1436 491300 1448
rect 491352 1436 491358 1488
rect 9306 1368 9312 1420
rect 9364 1408 9370 1420
rect 100754 1408 100760 1420
rect 9364 1380 100760 1408
rect 9364 1368 9370 1380
rect 100754 1368 100760 1380
rect 100812 1368 100818 1420
rect 102686 1368 102692 1420
rect 102744 1408 102750 1420
rect 111242 1408 111248 1420
rect 102744 1380 111248 1408
rect 102744 1368 102750 1380
rect 111242 1368 111248 1380
rect 111300 1368 111306 1420
rect 111518 1368 111524 1420
rect 111576 1408 111582 1420
rect 193582 1408 193588 1420
rect 111576 1380 193588 1408
rect 111576 1368 111582 1380
rect 193582 1368 193588 1380
rect 193640 1368 193646 1420
rect 193674 1368 193680 1420
rect 193732 1408 193738 1420
rect 243630 1408 243636 1420
rect 193732 1380 243636 1408
rect 193732 1368 193738 1380
rect 243630 1368 243636 1380
rect 243688 1368 243694 1420
rect 243722 1368 243728 1420
rect 243780 1408 243786 1420
rect 293586 1408 293592 1420
rect 243780 1380 293592 1408
rect 243780 1368 243786 1380
rect 293586 1368 293592 1380
rect 293644 1368 293650 1420
rect 295334 1368 295340 1420
rect 295392 1408 295398 1420
rect 493594 1408 493600 1420
rect 295392 1380 493600 1408
rect 295392 1368 295398 1380
rect 493594 1368 493600 1380
rect 493652 1368 493658 1420
rect 95970 1300 95976 1352
rect 96028 1340 96034 1352
rect 116578 1340 116584 1352
rect 96028 1312 116584 1340
rect 96028 1300 96034 1312
rect 116578 1300 116584 1312
rect 116636 1300 116642 1352
rect 35986 1232 35992 1284
rect 36044 1272 36050 1284
rect 112714 1272 112720 1284
rect 36044 1244 112720 1272
rect 36044 1232 36050 1244
rect 112714 1232 112720 1244
rect 112772 1232 112778 1284
rect 39298 1164 39304 1216
rect 39356 1204 39362 1216
rect 112622 1204 112628 1216
rect 39356 1176 112628 1204
rect 39356 1164 39362 1176
rect 112622 1164 112628 1176
rect 112680 1164 112686 1216
rect 62666 1096 62672 1148
rect 62724 1136 62730 1148
rect 117130 1136 117136 1148
rect 62724 1108 117136 1136
rect 62724 1096 62730 1108
rect 117130 1096 117136 1108
rect 117188 1096 117194 1148
rect 69290 1028 69296 1080
rect 69348 1068 69354 1080
rect 114094 1068 114100 1080
rect 69348 1040 114100 1068
rect 69348 1028 69354 1040
rect 114094 1028 114100 1040
rect 114152 1028 114158 1080
rect 76006 960 76012 1012
rect 76064 1000 76070 1012
rect 114002 1000 114008 1012
rect 76064 972 114008 1000
rect 76064 960 76070 972
rect 114002 960 114008 972
rect 114060 960 114066 1012
rect 82630 892 82636 944
rect 82688 932 82694 944
rect 113910 932 113916 944
rect 82688 904 113916 932
rect 82688 892 82694 904
rect 113910 892 113916 904
rect 113968 892 113974 944
rect 89346 824 89352 876
rect 89404 864 89410 876
rect 113818 864 113824 876
rect 89404 836 113824 864
rect 89404 824 89410 836
rect 113818 824 113824 836
rect 113876 824 113882 876
rect 22646 756 22652 808
rect 22704 796 22710 808
rect 114186 796 114192 808
rect 22704 768 114192 796
rect 22704 756 22710 768
rect 114186 756 114192 768
rect 114244 756 114250 808
<< via1 >>
rect 43260 162596 43312 162648
rect 151912 162596 151964 162648
rect 39856 162528 39908 162580
rect 149428 162528 149480 162580
rect 108856 162460 108908 162512
rect 202052 162460 202104 162512
rect 102140 162392 102192 162444
rect 196900 162392 196952 162444
rect 95424 162324 95476 162376
rect 190736 162324 190788 162376
rect 98736 162256 98788 162308
rect 193404 162256 193456 162308
rect 92020 162188 92072 162240
rect 189172 162188 189224 162240
rect 88708 162120 88760 162172
rect 186320 162120 186372 162172
rect 81900 162052 81952 162104
rect 181076 162052 181128 162104
rect 71872 161984 71924 162036
rect 172704 161984 172756 162036
rect 78588 161916 78640 161968
rect 178224 161916 178276 161968
rect 75184 161848 75236 161900
rect 175556 161848 175608 161900
rect 68468 161780 68520 161832
rect 171324 161780 171376 161832
rect 65156 161712 65208 161764
rect 168472 161712 168524 161764
rect 56692 161644 56744 161696
rect 161480 161644 161532 161696
rect 61752 161576 61804 161628
rect 165620 161576 165672 161628
rect 115572 161508 115624 161560
rect 207020 161508 207072 161560
rect 112260 161440 112312 161492
rect 204260 161440 204312 161492
rect 114744 161372 114796 161424
rect 206560 161372 206612 161424
rect 108028 161304 108080 161356
rect 200304 161304 200356 161356
rect 101312 161236 101364 161288
rect 196256 161236 196308 161288
rect 94596 161168 94648 161220
rect 191104 161168 191156 161220
rect 205548 161168 205600 161220
rect 275836 161168 275888 161220
rect 81072 161100 81124 161152
rect 180892 161100 180944 161152
rect 198832 161100 198884 161152
rect 270500 161100 270552 161152
rect 67640 161032 67692 161084
rect 169852 161032 169904 161084
rect 183744 161032 183796 161084
rect 258080 161032 258132 161084
rect 60924 160964 60976 161016
rect 165436 160964 165488 161016
rect 175280 160964 175332 161016
rect 252744 160964 252796 161016
rect 54208 160896 54260 160948
rect 160284 160896 160336 160948
rect 161848 160896 161900 160948
rect 242072 160896 242124 160948
rect 47492 160828 47544 160880
rect 155040 160828 155092 160880
rect 166080 160828 166132 160880
rect 245752 160828 245804 160880
rect 40684 160760 40736 160812
rect 149152 160760 149204 160812
rect 155132 160760 155184 160812
rect 237380 160760 237432 160812
rect 36544 160692 36596 160744
rect 146852 160692 146904 160744
rect 148416 160692 148468 160744
rect 231952 160692 232004 160744
rect 124864 160624 124916 160676
rect 213920 160624 213972 160676
rect 141700 160556 141752 160608
rect 227076 160556 227128 160608
rect 149244 160488 149296 160540
rect 232872 160488 232924 160540
rect 93676 160012 93728 160064
rect 165528 160012 165580 160064
rect 181168 160012 181220 160064
rect 230756 160012 230808 160064
rect 240876 160012 240928 160064
rect 263876 160012 263928 160064
rect 265348 160012 265400 160064
rect 311072 160012 311124 160064
rect 318340 160012 318392 160064
rect 336648 160012 336700 160064
rect 342720 160012 342772 160064
rect 372620 160012 372672 160064
rect 409144 160012 409196 160064
rect 86960 159944 87012 159996
rect 158720 159944 158772 159996
rect 164332 159944 164384 159996
rect 222016 159944 222068 159996
rect 234160 159944 234212 159996
rect 255504 159944 255556 159996
rect 258540 159944 258592 159996
rect 305000 159944 305052 159996
rect 311532 159944 311584 159996
rect 330208 159944 330260 159996
rect 332600 159944 332652 159996
rect 368572 159944 368624 159996
rect 386420 159944 386472 159996
rect 412824 159944 412876 159996
rect 425980 160012 426032 160064
rect 426440 160012 426492 160064
rect 431224 159944 431276 159996
rect 484860 159944 484912 159996
rect 489000 159944 489052 159996
rect 76932 159876 76984 159928
rect 147772 159876 147824 159928
rect 150900 159876 150952 159928
rect 207112 159876 207164 159928
rect 208952 159876 209004 159928
rect 220176 159876 220228 159928
rect 222384 159876 222436 159928
rect 225696 159876 225748 159928
rect 70124 159808 70176 159860
rect 140872 159808 140924 159860
rect 171140 159808 171192 159860
rect 230388 159876 230440 159928
rect 238392 159876 238444 159928
rect 288256 159876 288308 159928
rect 291384 159876 291436 159928
rect 311900 159876 311952 159928
rect 325884 159876 325936 159928
rect 362132 159876 362184 159928
rect 393136 159876 393188 159928
rect 419080 159876 419132 159928
rect 231676 159808 231728 159860
rect 284392 159808 284444 159860
rect 305644 159808 305696 159860
rect 345940 159808 345992 159860
rect 375472 159808 375524 159860
rect 405556 159808 405608 159860
rect 406660 159808 406712 159860
rect 429384 159808 429436 159860
rect 472256 159808 472308 159860
rect 479432 159808 479484 159860
rect 46572 159740 46624 159792
rect 120172 159740 120224 159792
rect 124036 159740 124088 159792
rect 187700 159740 187752 159792
rect 194692 159740 194744 159792
rect 212632 159740 212684 159792
rect 218244 159740 218296 159792
rect 272524 159740 272576 159792
rect 277952 159740 278004 159792
rect 287060 159740 287112 159792
rect 287980 159740 288032 159792
rect 288624 159740 288676 159792
rect 298928 159740 298980 159792
rect 343640 159740 343692 159792
rect 368756 159740 368808 159792
rect 400404 159740 400456 159792
rect 402428 159740 402480 159792
rect 426164 159740 426216 159792
rect 481456 159740 481508 159792
rect 485780 159740 485832 159792
rect 492404 159740 492456 159792
rect 494796 159740 494848 159792
rect 53380 159672 53432 159724
rect 128360 159672 128412 159724
rect 130752 159672 130804 159724
rect 195244 159672 195296 159724
rect 211436 159672 211488 159724
rect 268936 159672 268988 159724
rect 282092 159672 282144 159724
rect 291108 159672 291160 159724
rect 292212 159672 292264 159724
rect 338396 159672 338448 159724
rect 346032 159672 346084 159724
rect 378324 159672 378376 159724
rect 382188 159672 382240 159724
rect 408500 159672 408552 159724
rect 413376 159672 413428 159724
rect 434444 159672 434496 159724
rect 478972 159672 479024 159724
rect 484400 159672 484452 159724
rect 3700 159604 3752 159656
rect 77208 159604 77260 159656
rect 80244 159604 80296 159656
rect 156052 159604 156104 159656
rect 157616 159604 157668 159656
rect 216864 159604 216916 159656
rect 224960 159604 225012 159656
rect 281172 159604 281224 159656
rect 285496 159604 285548 159656
rect 332600 159604 332652 159656
rect 352748 159604 352800 159656
rect 385960 159604 386012 159656
rect 388996 159604 389048 159656
rect 414296 159604 414348 159656
rect 420092 159604 420144 159656
rect 435824 159604 435876 159656
rect 441068 159604 441120 159656
rect 445484 159604 445536 159656
rect 478144 159604 478196 159656
rect 483020 159604 483072 159656
rect 33968 159536 34020 159588
rect 63500 159536 63552 159588
rect 66812 159536 66864 159588
rect 144828 159536 144880 159588
rect 170220 159536 170272 159588
rect 176660 159536 176712 159588
rect 198004 159536 198056 159588
rect 260748 159536 260800 159588
rect 272064 159536 272116 159588
rect 320732 159536 320784 159588
rect 339316 159536 339368 159588
rect 377956 159536 378008 159588
rect 379704 159536 379756 159588
rect 408776 159536 408828 159588
rect 431868 159536 431920 159588
rect 436560 159536 436612 159588
rect 2872 159468 2924 159520
rect 92480 159468 92532 159520
rect 100484 159468 100536 159520
rect 169760 159468 169812 159520
rect 184572 159468 184624 159520
rect 247224 159468 247276 159520
rect 251824 159468 251876 159520
rect 301688 159468 301740 159520
rect 308220 159468 308272 159520
rect 317788 159468 317840 159520
rect 319168 159468 319220 159520
rect 361580 159468 361632 159520
rect 366272 159468 366324 159520
rect 398472 159468 398524 159520
rect 399852 159468 399904 159520
rect 424232 159468 424284 159520
rect 433524 159468 433576 159520
rect 449808 159468 449860 159520
rect 451188 159468 451240 159520
rect 455328 159468 455380 159520
rect 26424 159400 26476 159452
rect 129832 159400 129884 159452
rect 139124 159400 139176 159452
rect 157432 159400 157484 159452
rect 177856 159400 177908 159452
rect 242440 159400 242492 159452
rect 245108 159400 245160 159452
rect 299388 159400 299440 159452
rect 312452 159400 312504 159452
rect 355692 159400 355744 159452
rect 359556 159400 359608 159452
rect 393412 159400 393464 159452
rect 395712 159400 395764 159452
rect 421104 159400 421156 159452
rect 432696 159400 432748 159452
rect 447140 159400 447192 159452
rect 479800 159400 479852 159452
rect 485228 159400 485280 159452
rect 496636 159400 496688 159452
rect 498016 159400 498068 159452
rect 12992 159332 13044 159384
rect 124128 159332 124180 159384
rect 132408 159332 132460 159384
rect 135812 159332 135864 159384
rect 140780 159332 140832 159384
rect 174912 159332 174964 159384
rect 191288 159332 191340 159384
rect 256792 159332 256844 159384
rect 261944 159332 261996 159384
rect 263508 159332 263560 159384
rect 287060 159332 287112 159384
rect 291476 159332 291528 159384
rect 331772 159332 331824 159384
rect 372068 159332 372120 159384
rect 372988 159332 373040 159384
rect 403164 159332 403216 159384
rect 434352 159332 434404 159384
rect 450084 159332 450136 159384
rect 461308 159332 461360 159384
rect 464896 159332 464948 159384
rect 477316 159332 477368 159384
rect 483296 159332 483348 159384
rect 497464 159332 497516 159384
rect 498660 159332 498712 159384
rect 49976 159264 50028 159316
rect 109224 159264 109276 159316
rect 110512 159264 110564 159316
rect 179420 159264 179472 159316
rect 187884 159264 187936 159316
rect 210884 159264 210936 159316
rect 214840 159264 214892 159316
rect 223948 159264 224000 159316
rect 227444 159264 227496 159316
rect 247040 159264 247092 159316
rect 261116 159264 261168 159316
rect 269028 159264 269080 159316
rect 271236 159264 271288 159316
rect 296812 159264 296864 159316
rect 298100 159264 298152 159316
rect 311992 159264 312044 159316
rect 325056 159264 325108 159316
rect 352012 159264 352064 159316
rect 480628 159264 480680 159316
rect 485872 159264 485924 159316
rect 494980 159264 495032 159316
rect 496728 159264 496780 159316
rect 76012 159196 76064 159248
rect 79968 159196 80020 159248
rect 120632 159196 120684 159248
rect 184848 159196 184900 159248
rect 208124 159196 208176 159248
rect 222108 159196 222160 159248
rect 228272 159196 228324 159248
rect 239956 159196 240008 159248
rect 250996 159196 251048 159248
rect 274640 159196 274692 159248
rect 284668 159196 284720 159248
rect 305460 159196 305512 159248
rect 489920 159196 489972 159248
rect 492680 159196 492732 159248
rect 37372 159128 37424 159180
rect 38568 159128 38620 159180
rect 127348 159128 127400 159180
rect 143080 159128 143132 159180
rect 144184 159128 144236 159180
rect 193128 159128 193180 159180
rect 201408 159128 201460 159180
rect 212356 159128 212408 159180
rect 237564 159128 237616 159180
rect 251732 159128 251784 159180
rect 257712 159128 257764 159180
rect 279884 159128 279936 159180
rect 304816 159128 304868 159180
rect 324320 159128 324372 159180
rect 493232 159128 493284 159180
rect 495440 159128 495492 159180
rect 91192 159060 91244 159112
rect 92388 159060 92440 159112
rect 155960 159060 156012 159112
rect 197360 159060 197412 159112
rect 214012 159060 214064 159112
rect 216680 159060 216732 159112
rect 217324 159060 217376 159112
rect 223488 159060 223540 159112
rect 247684 159060 247736 159112
rect 262128 159060 262180 159112
rect 264428 159060 264480 159112
rect 284300 159060 284352 159112
rect 426808 159060 426860 159112
rect 433064 159060 433116 159112
rect 471428 159060 471480 159112
rect 477684 159060 477736 159112
rect 484032 159060 484084 159112
rect 488448 159060 488500 159112
rect 174452 158992 174504 159044
rect 204168 158992 204220 159044
rect 210608 158992 210660 159044
rect 215024 158992 215076 159044
rect 267832 158992 267884 159044
rect 279516 158992 279568 159044
rect 390652 158992 390704 159044
rect 391848 158992 391900 159044
rect 453764 158992 453816 159044
rect 458180 158992 458232 159044
rect 473084 158992 473136 159044
rect 478972 158992 479024 159044
rect 486516 158992 486568 159044
rect 490288 158992 490340 159044
rect 118976 158924 119028 158976
rect 125508 158924 125560 158976
rect 224132 158924 224184 158976
rect 227720 158924 227772 158976
rect 278780 158924 278832 158976
rect 275376 158856 275428 158908
rect 278688 158856 278740 158908
rect 327540 158924 327592 158976
rect 328368 158924 328420 158976
rect 362040 158924 362092 158976
rect 366824 158924 366876 158976
rect 372160 158924 372212 158976
rect 374276 158924 374328 158976
rect 437756 158924 437808 158976
rect 444288 158924 444340 158976
rect 447876 158924 447928 158976
rect 452476 158924 452528 158976
rect 463792 158924 463844 158976
rect 471796 158924 471848 158976
rect 475568 158924 475620 158976
rect 481640 158924 481692 158976
rect 487344 158924 487396 158976
rect 489920 158924 489972 158976
rect 491576 158924 491628 158976
rect 494152 158924 494204 158976
rect 331772 158856 331824 158908
rect 473912 158856 473964 158908
rect 480260 158856 480312 158908
rect 482284 158856 482336 158908
rect 487160 158856 487212 158908
rect 489092 158856 489144 158908
rect 491300 158856 491352 158908
rect 121460 158788 121512 158840
rect 122748 158788 122800 158840
rect 129004 158788 129056 158840
rect 132132 158788 132184 158840
rect 145840 158788 145892 158840
rect 150440 158788 150492 158840
rect 241796 158788 241848 158840
rect 244556 158788 244608 158840
rect 315764 158788 315816 158840
rect 318708 158788 318760 158840
rect 378876 158788 378928 158840
rect 380992 158788 381044 158840
rect 389824 158788 389876 158840
rect 391572 158788 391624 158840
rect 405740 158788 405792 158840
rect 406936 158788 406988 158840
rect 436100 158788 436152 158840
rect 438860 158788 438912 158840
rect 449532 158788 449584 158840
rect 453948 158788 454000 158840
rect 474740 158788 474792 158840
rect 481364 158788 481416 158840
rect 483204 158788 483256 158840
rect 487528 158788 487580 158840
rect 488172 158788 488224 158840
rect 491576 158788 491628 158840
rect 388 158720 440 158772
rect 2044 158720 2096 158772
rect 64236 158720 64288 158772
rect 64788 158720 64840 158772
rect 65984 158720 66036 158772
rect 71044 158720 71096 158772
rect 71688 158720 71740 158772
rect 77760 158720 77812 158772
rect 78588 158720 78640 158772
rect 84476 158720 84528 158772
rect 85488 158720 85540 158772
rect 103796 158720 103848 158772
rect 109040 158720 109092 158772
rect 116400 158720 116452 158772
rect 119528 158720 119580 158772
rect 131580 158720 131632 158772
rect 132408 158720 132460 158772
rect 145012 158720 145064 158772
rect 146208 158720 146260 158772
rect 152556 158720 152608 158772
rect 153108 158720 153160 158772
rect 165252 158720 165304 158772
rect 167644 158720 167696 158772
rect 196348 158720 196400 158772
rect 198740 158720 198792 158772
rect 202236 158720 202288 158772
rect 202788 158720 202840 158772
rect 203064 158720 203116 158772
rect 208492 158720 208544 158772
rect 220728 158720 220780 158772
rect 227904 158720 227956 158772
rect 230848 158720 230900 158772
rect 238024 158720 238076 158772
rect 248512 158720 248564 158772
rect 249616 158720 249668 158772
rect 256884 158720 256936 158772
rect 257988 158720 258040 158772
rect 268660 158720 268712 158772
rect 271696 158720 271748 158772
rect 286324 158720 286376 158772
rect 286876 158720 286928 158772
rect 288900 158720 288952 158772
rect 292304 158720 292356 158772
rect 301504 158720 301556 158772
rect 304816 158720 304868 158772
rect 336004 158720 336056 158772
rect 337752 158720 337804 158772
rect 385592 158720 385644 158772
rect 389088 158720 389140 158772
rect 430212 158720 430264 158772
rect 433248 158720 433300 158772
rect 458732 158720 458784 158772
rect 463332 158720 463384 158772
rect 476396 158720 476448 158772
rect 482652 158720 482704 158772
rect 485688 158720 485740 158772
rect 488632 158720 488684 158772
rect 490748 158720 490800 158772
rect 493508 158720 493560 158772
rect 494060 158720 494112 158772
rect 495716 158720 495768 158772
rect 495808 158720 495860 158772
rect 497004 158720 497056 158772
rect 499672 158720 499724 158772
rect 500592 158720 500644 158772
rect 504456 158720 504508 158772
rect 505008 158720 505060 158772
rect 86132 158652 86184 158704
rect 183560 158652 183612 158704
rect 195244 158652 195296 158704
rect 218704 158652 218756 158704
rect 220176 158652 220228 158704
rect 277952 158652 278004 158704
rect 321652 158652 321704 158704
rect 359464 158652 359516 158704
rect 168380 158584 168432 158636
rect 169760 158584 169812 158636
rect 194600 158584 194652 158636
rect 200580 158584 200632 158636
rect 272064 158584 272116 158636
rect 279608 158584 279660 158636
rect 331312 158584 331364 158636
rect 351920 158584 351972 158636
rect 386512 158584 386564 158636
rect 62580 158516 62632 158568
rect 166724 158516 166776 158568
rect 190460 158516 190512 158568
rect 263784 158516 263836 158568
rect 274548 158516 274600 158568
rect 328552 158516 328604 158568
rect 351092 158516 351144 158568
rect 386972 158516 387024 158568
rect 29828 158448 29880 158500
rect 55772 158448 55824 158500
rect 59268 158448 59320 158500
rect 163044 158448 163096 158500
rect 165528 158448 165580 158500
rect 190552 158448 190604 158500
rect 197176 158448 197228 158500
rect 269396 158448 269448 158500
rect 272892 158448 272944 158500
rect 327080 158448 327132 158500
rect 338488 158448 338540 158500
rect 376852 158448 376904 158500
rect 377220 158448 377272 158500
rect 406844 158448 406896 158500
rect 52460 158380 52512 158432
rect 45744 158312 45796 158364
rect 153384 158312 153436 158364
rect 158720 158380 158772 158432
rect 185032 158380 185084 158432
rect 187056 158380 187108 158432
rect 260840 158380 260892 158432
rect 266176 158380 266228 158432
rect 322112 158380 322164 158432
rect 330116 158380 330168 158432
rect 370872 158380 370924 158432
rect 158996 158312 159048 158364
rect 177028 158312 177080 158364
rect 254032 158312 254084 158364
rect 256056 158312 256108 158364
rect 314384 158312 314436 158364
rect 320824 158312 320876 158364
rect 363512 158312 363564 158364
rect 378048 158312 378100 158364
rect 407396 158312 407448 158364
rect 42432 158244 42484 158296
rect 150532 158244 150584 158296
rect 173624 158244 173676 158296
rect 251456 158244 251508 158296
rect 252652 158244 252704 158296
rect 310612 158244 310664 158296
rect 317420 158244 317472 158296
rect 360200 158244 360252 158296
rect 367100 158244 367152 158296
rect 399116 158244 399168 158296
rect 426440 158244 426492 158296
rect 443000 158244 443052 158296
rect 31484 158176 31536 158228
rect 139492 158176 139544 158228
rect 163504 158176 163556 158228
rect 242900 158176 242952 158228
rect 245936 158176 245988 158228
rect 306380 158176 306432 158228
rect 314108 158176 314160 158228
rect 357624 158176 357676 158228
rect 361212 158176 361264 158228
rect 394700 158176 394752 158228
rect 404912 158176 404964 158228
rect 428004 158176 428056 158228
rect 439412 158176 439464 158228
rect 454408 158176 454460 158228
rect 32312 158108 32364 158160
rect 143632 158108 143684 158160
rect 153476 158108 153528 158160
rect 236092 158108 236144 158160
rect 242624 158108 242676 158160
rect 304080 158108 304132 158160
rect 307392 158108 307444 158160
rect 353300 158108 353352 158160
rect 358636 158108 358688 158160
rect 391940 158108 391992 158160
rect 404084 158108 404136 158160
rect 427360 158108 427412 158160
rect 428464 158108 428516 158160
rect 445760 158108 445812 158160
rect 448704 158108 448756 158160
rect 461400 158108 461452 158160
rect 18880 158040 18932 158092
rect 132500 158040 132552 158092
rect 139952 158040 140004 158092
rect 224960 158040 225012 158092
rect 229100 158040 229152 158092
rect 292764 158040 292816 158092
rect 293040 158040 293092 158092
rect 342260 158040 342312 158092
rect 350264 158040 350316 158092
rect 385224 158040 385276 158092
rect 393964 158040 394016 158092
rect 419540 158040 419592 158092
rect 420920 158040 420972 158092
rect 440332 158040 440384 158092
rect 443644 158040 443696 158092
rect 456800 158040 456852 158092
rect 466368 158040 466420 158092
rect 474924 158040 474976 158092
rect 2136 157972 2188 158024
rect 120080 157972 120132 158024
rect 133236 157972 133288 158024
rect 220636 157972 220688 158024
rect 225696 157972 225748 158024
rect 288440 157972 288492 158024
rect 289728 157972 289780 158024
rect 340052 157972 340104 158024
rect 340144 157972 340196 158024
rect 378600 157972 378652 158024
rect 388076 157972 388128 158024
rect 414572 157972 414624 158024
rect 415032 157972 415084 158024
rect 434720 157972 434772 158024
rect 435180 157972 435232 158024
rect 451096 157972 451148 158024
rect 457904 157972 457956 158024
rect 468484 157972 468536 158024
rect 99564 157904 99616 157956
rect 194968 157904 195020 157956
rect 207112 157904 207164 157956
rect 233240 157904 233292 157956
rect 239220 157904 239272 157956
rect 256700 157904 256752 157956
rect 262772 157904 262824 157956
rect 319536 157904 319588 157956
rect 324320 157904 324372 157956
rect 350540 157904 350592 157956
rect 106372 157836 106424 157888
rect 200120 157836 200172 157888
rect 221556 157836 221608 157888
rect 245660 157836 245712 157888
rect 259460 157836 259512 157888
rect 316960 157836 317012 157888
rect 123116 157768 123168 157820
rect 207112 157768 207164 157820
rect 269488 157768 269540 157820
rect 324688 157768 324740 157820
rect 144828 157700 144880 157752
rect 169944 157700 169996 157752
rect 201316 157700 201368 157752
rect 223856 157700 223908 157752
rect 311900 157700 311952 157752
rect 341340 157700 341392 157752
rect 79968 157292 80020 157344
rect 177028 157292 177080 157344
rect 193772 157292 193824 157344
rect 266912 157292 266964 157344
rect 296444 157292 296496 157344
rect 345020 157292 345072 157344
rect 356152 157292 356204 157344
rect 358912 157292 358964 157344
rect 69296 157224 69348 157276
rect 171140 157224 171192 157276
rect 179512 157224 179564 157276
rect 255872 157224 255924 157276
rect 276204 157224 276256 157276
rect 329840 157224 329892 157276
rect 352012 157224 352064 157276
rect 365904 157224 365956 157276
rect 4528 157156 4580 157208
rect 109132 157156 109184 157208
rect 113088 157156 113140 157208
rect 205272 157156 205324 157208
rect 209780 157156 209832 157208
rect 278780 157156 278832 157208
rect 288624 157156 288676 157208
rect 338672 157156 338724 157208
rect 347780 157156 347832 157208
rect 383660 157156 383712 157208
rect 55864 157088 55916 157140
rect 161572 157088 161624 157140
rect 172796 157088 172848 157140
rect 250812 157088 250864 157140
rect 260288 157088 260340 157140
rect 317420 157088 317472 157140
rect 346860 157088 346912 157140
rect 383752 157088 383804 157140
rect 49148 157020 49200 157072
rect 156420 157020 156472 157072
rect 176108 157020 176160 157072
rect 252560 157020 252612 157072
rect 254400 157020 254452 157072
rect 311900 157020 311952 157072
rect 336832 157020 336884 157072
rect 376024 157020 376076 157072
rect 383108 157020 383160 157072
rect 411352 157020 411404 157072
rect 39028 156952 39080 157004
rect 147680 156952 147732 157004
rect 169392 156952 169444 157004
rect 247132 156952 247184 157004
rect 253572 156952 253624 157004
rect 307024 156952 307076 157004
rect 330944 156952 330996 157004
rect 371240 156952 371292 157004
rect 374644 156952 374696 157004
rect 404452 156952 404504 157004
rect 423404 156952 423456 157004
rect 442172 156952 442224 157004
rect 464896 156952 464948 157004
rect 471060 156952 471112 157004
rect 28080 156884 28132 156936
rect 139400 156884 139452 156936
rect 160192 156884 160244 156936
rect 240140 156884 240192 156936
rect 249340 156884 249392 156936
rect 306380 156884 306432 156936
rect 24768 156816 24820 156868
rect 137836 156816 137888 156868
rect 150072 156816 150124 156868
rect 233516 156816 233568 156868
rect 246764 156816 246816 156868
rect 307300 156884 307352 156936
rect 310704 156884 310756 156936
rect 356152 156884 356204 156936
rect 373816 156884 373868 156936
rect 404084 156884 404136 156936
rect 411628 156884 411680 156936
rect 433156 156884 433208 156936
rect 436560 156884 436612 156936
rect 448612 156884 448664 156936
rect 306656 156816 306708 156868
rect 351920 156816 351972 156868
rect 363696 156816 363748 156868
rect 396540 156816 396592 156868
rect 400772 156816 400824 156868
rect 423772 156816 423824 156868
rect 433248 156816 433300 156868
rect 447324 156816 447376 156868
rect 18052 156748 18104 156800
rect 132684 156748 132736 156800
rect 136640 156748 136692 156800
rect 222752 156748 222804 156800
rect 240048 156748 240100 156800
rect 302240 156748 302292 156800
rect 303160 156748 303212 156800
rect 349252 156748 349304 156800
rect 357808 156748 357860 156800
rect 392124 156748 392176 156800
rect 401600 156748 401652 156800
rect 425152 156748 425204 156800
rect 427636 156748 427688 156800
rect 444380 156748 444432 156800
rect 11244 156680 11296 156732
rect 125692 156680 125744 156732
rect 126520 156680 126572 156732
rect 215484 156680 215536 156732
rect 216680 156680 216732 156732
rect 282092 156680 282144 156732
rect 283012 156680 283064 156732
rect 334900 156680 334952 156732
rect 341892 156680 341944 156732
rect 379888 156680 379940 156732
rect 384764 156680 384816 156732
rect 412640 156680 412692 156732
rect 419264 156680 419316 156732
rect 438952 156680 439004 156732
rect 446128 156680 446180 156732
rect 459468 156680 459520 156732
rect 14648 156612 14700 156664
rect 129740 156612 129792 156664
rect 129924 156612 129976 156664
rect 218060 156612 218112 156664
rect 236736 156612 236788 156664
rect 299664 156612 299716 156664
rect 299756 156612 299808 156664
rect 347780 156612 347832 156664
rect 348608 156612 348660 156664
rect 385040 156612 385092 156664
rect 387248 156612 387300 156664
rect 414112 156612 414164 156664
rect 414204 156612 414256 156664
rect 435088 156612 435140 156664
rect 445300 156612 445352 156664
rect 96252 156544 96304 156596
rect 192392 156544 192444 156596
rect 215024 156544 215076 156596
rect 279332 156544 279384 156596
rect 303988 156544 304040 156596
rect 351000 156544 351052 156596
rect 458180 156612 458232 156664
rect 465264 156612 465316 156664
rect 458364 156544 458416 156596
rect 109684 156476 109736 156528
rect 194324 156476 194376 156528
rect 227720 156476 227772 156528
rect 290004 156476 290056 156528
rect 307024 156476 307076 156528
rect 312452 156476 312504 156528
rect 317788 156476 317840 156528
rect 354220 156476 354272 156528
rect 133420 156408 133472 156460
rect 164424 156408 164476 156460
rect 176660 156408 176712 156460
rect 248880 156408 248932 156460
rect 251732 156408 251784 156460
rect 299480 156408 299532 156460
rect 306380 156408 306432 156460
rect 309232 156408 309284 156460
rect 311992 156408 312044 156460
rect 346492 156408 346544 156460
rect 140872 156340 140924 156392
rect 172520 156340 172572 156392
rect 279516 156340 279568 156392
rect 323400 156340 323452 156392
rect 89536 155864 89588 155916
rect 187240 155864 187292 155916
rect 203892 155864 203944 155916
rect 273444 155864 273496 155916
rect 324228 155864 324280 155916
rect 366272 155864 366324 155916
rect 85304 155796 85356 155848
rect 184020 155796 184072 155848
rect 206468 155796 206520 155848
rect 276480 155796 276532 155848
rect 287152 155796 287204 155848
rect 296628 155796 296680 155848
rect 297272 155796 297324 155848
rect 345848 155796 345900 155848
rect 345940 155796 345992 155848
rect 352288 155796 352340 155848
rect 72700 155728 72752 155780
rect 174452 155728 174504 155780
rect 199660 155728 199712 155780
rect 271052 155728 271104 155780
rect 280436 155728 280488 155780
rect 333060 155728 333112 155780
rect 336648 155728 336700 155780
rect 361948 155728 362000 155780
rect 362132 155728 362184 155780
rect 367652 155728 367704 155780
rect 370412 155728 370464 155780
rect 401692 155728 401744 155780
rect 55036 155660 55088 155712
rect 157340 155660 157392 155712
rect 192944 155660 192996 155712
rect 265164 155660 265216 155712
rect 273720 155660 273772 155712
rect 327908 155660 327960 155712
rect 328368 155660 328420 155712
rect 368940 155660 368992 155712
rect 369584 155660 369636 155712
rect 400220 155660 400272 155712
rect 48320 155592 48372 155644
rect 154672 155592 154724 155644
rect 186228 155592 186280 155644
rect 261116 155592 261168 155644
rect 277124 155592 277176 155644
rect 330484 155592 330536 155644
rect 334256 155592 334308 155644
rect 374092 155592 374144 155644
rect 378324 155592 378376 155644
rect 383108 155592 383160 155644
rect 41604 155524 41656 155576
rect 150624 155524 150676 155576
rect 156788 155524 156840 155576
rect 237932 155524 237984 155576
rect 238024 155524 238076 155576
rect 23940 155456 23992 155508
rect 136732 155456 136784 155508
rect 138296 155456 138348 155508
rect 221740 155456 221792 155508
rect 225788 155456 225840 155508
rect 291292 155456 291344 155508
rect 22192 155388 22244 155440
rect 135904 155388 135956 155440
rect 146668 155388 146720 155440
rect 230940 155388 230992 155440
rect 232504 155388 232556 155440
rect 294788 155524 294840 155576
rect 343916 155524 343968 155576
rect 364524 155524 364576 155576
rect 396172 155524 396224 155576
rect 293868 155456 293920 155508
rect 343272 155456 343324 155508
rect 353668 155456 353720 155508
rect 388352 155456 388404 155508
rect 408316 155456 408368 155508
rect 430580 155456 430632 155508
rect 433064 155456 433116 155508
rect 444748 155456 444800 155508
rect 15476 155320 15528 155372
rect 130292 155320 130344 155372
rect 135812 155320 135864 155372
rect 219532 155320 219584 155372
rect 223212 155320 223264 155372
rect 289360 155320 289412 155372
rect 295156 155388 295208 155440
rect 300676 155388 300728 155440
rect 348424 155388 348476 155440
rect 354496 155388 354548 155440
rect 389548 155388 389600 155440
rect 394884 155388 394936 155440
rect 420368 155388 420420 155440
rect 429292 155388 429344 155440
rect 446680 155388 446732 155440
rect 296444 155320 296496 155372
rect 8760 155252 8812 155304
rect 125600 155252 125652 155304
rect 125784 155252 125836 155304
rect 214840 155252 214892 155304
rect 219072 155252 219124 155304
rect 286140 155252 286192 155304
rect 290556 155252 290608 155304
rect 339592 155320 339644 155372
rect 345204 155320 345256 155372
rect 382280 155320 382332 155372
rect 397368 155320 397420 155372
rect 422300 155320 422352 155372
rect 424324 155320 424376 155372
rect 441712 155320 441764 155372
rect 444472 155320 444524 155372
rect 458180 155320 458232 155372
rect 296628 155252 296680 155304
rect 338120 155252 338172 155304
rect 344376 155252 344428 155304
rect 381452 155252 381504 155304
rect 383936 155252 383988 155304
rect 411996 155252 412048 155304
rect 421748 155252 421800 155304
rect 440884 155252 440936 155304
rect 441988 155252 442040 155304
rect 1216 155184 1268 155236
rect 118792 155184 118844 155236
rect 119528 155184 119580 155236
rect 207572 155184 207624 155236
rect 216496 155184 216548 155236
rect 283104 155184 283156 155236
rect 283840 155184 283892 155236
rect 335544 155184 335596 155236
rect 343548 155184 343600 155236
rect 380900 155184 380952 155236
rect 381360 155184 381412 155236
rect 410064 155184 410116 155236
rect 410800 155184 410852 155236
rect 432052 155184 432104 155236
rect 442816 155184 442868 155236
rect 456248 155252 456300 155304
rect 467104 155252 467156 155304
rect 92480 155116 92532 155168
rect 121092 155116 121144 155168
rect 150440 155116 150492 155168
rect 229192 155116 229244 155168
rect 230020 155116 230072 155168
rect 294052 155116 294104 155168
rect 330208 155116 330260 155168
rect 356796 155116 356848 155168
rect 456340 155184 456392 155236
rect 456984 155116 457036 155168
rect 128176 155048 128228 155100
rect 198096 155048 198148 155100
rect 226616 155048 226668 155100
rect 291200 155048 291252 155100
rect 291476 155048 291528 155100
rect 330024 155048 330076 155100
rect 134892 154980 134944 155032
rect 201868 154980 201920 155032
rect 269028 154980 269080 155032
rect 317972 154980 318024 155032
rect 118148 154912 118200 154964
rect 144828 154912 144880 154964
rect 157432 154912 157484 154964
rect 225144 154912 225196 154964
rect 262128 154912 262180 154964
rect 307944 154912 307996 154964
rect 105452 154504 105504 154556
rect 199476 154504 199528 154556
rect 215668 154504 215720 154556
rect 283564 154504 283616 154556
rect 284300 154504 284352 154556
rect 320916 154504 320968 154556
rect 338396 154504 338448 154556
rect 341984 154504 342036 154556
rect 463332 154504 463384 154556
rect 468944 154504 468996 154556
rect 471796 154504 471848 154556
rect 472992 154504 473044 154556
rect 103428 154436 103480 154488
rect 197544 154436 197596 154488
rect 213184 154436 213236 154488
rect 281632 154436 281684 154488
rect 313280 154436 313332 154488
rect 358084 154436 358136 154488
rect 366824 154436 366876 154488
rect 395344 154436 395396 154488
rect 92848 154368 92900 154420
rect 189816 154368 189868 154420
rect 198740 154368 198792 154420
rect 268844 154368 268896 154420
rect 281540 154368 281592 154420
rect 333704 154368 333756 154420
rect 335084 154368 335136 154420
rect 338948 154368 339000 154420
rect 340972 154368 341024 154420
rect 379244 154368 379296 154420
rect 58348 154300 58400 154352
rect 163504 154300 163556 154352
rect 192116 154300 192168 154352
rect 265716 154300 265768 154352
rect 270316 154300 270368 154352
rect 325332 154300 325384 154352
rect 333428 154300 333480 154352
rect 373448 154300 373500 154352
rect 51632 154232 51684 154284
rect 155960 154232 156012 154284
rect 188804 154232 188856 154284
rect 263048 154232 263100 154284
rect 267004 154232 267056 154284
rect 322848 154232 322900 154284
rect 326988 154232 327040 154284
rect 368296 154232 368348 154284
rect 44916 154164 44968 154216
rect 153200 154164 153252 154216
rect 154304 154164 154356 154216
rect 182364 154164 182416 154216
rect 185400 154164 185452 154216
rect 260472 154164 260524 154216
rect 263600 154164 263652 154216
rect 320180 154164 320232 154216
rect 323308 154164 323360 154216
rect 365720 154164 365772 154216
rect 371332 154164 371384 154216
rect 402336 154164 402388 154216
rect 422576 154164 422628 154216
rect 34796 154096 34848 154148
rect 145564 154096 145616 154148
rect 147772 154096 147824 154148
rect 177672 154096 177724 154148
rect 181996 154096 182048 154148
rect 257896 154096 257948 154148
rect 257988 154096 258040 154148
rect 315028 154096 315080 154148
rect 319996 154096 320048 154148
rect 363236 154096 363288 154148
rect 368388 154096 368440 154148
rect 399760 154096 399812 154148
rect 407488 154096 407540 154148
rect 429936 154096 429988 154148
rect 25596 154028 25648 154080
rect 138480 154028 138532 154080
rect 172428 154028 172480 154080
rect 250168 154028 250220 154080
rect 250260 154028 250312 154080
rect 309876 154028 309928 154080
rect 316592 154028 316644 154080
rect 360660 154028 360712 154080
rect 20536 153960 20588 154012
rect 134616 153960 134668 154012
rect 143356 153960 143408 154012
rect 228364 153960 228416 154012
rect 243452 153960 243504 154012
rect 304724 153960 304776 154012
rect 304816 153960 304868 154012
rect 349068 153960 349120 154012
rect 360384 153960 360436 154012
rect 394056 154028 394108 154080
rect 398196 154028 398248 154080
rect 422944 154028 422996 154080
rect 438860 154164 438912 154216
rect 451832 154164 451884 154216
rect 431040 154096 431092 154148
rect 447968 154096 448020 154148
rect 441436 154028 441488 154080
rect 17132 153892 17184 153944
rect 132040 153892 132092 153944
rect 132132 153892 132184 153944
rect 217416 153892 217468 153944
rect 219900 153892 219952 153944
rect 286784 153892 286836 153944
rect 286876 153892 286928 153944
rect 337476 153892 337528 153944
rect 338028 153892 338080 153944
rect 360844 153892 360896 153944
rect 13820 153824 13872 153876
rect 129464 153824 129516 153876
rect 135720 153824 135772 153876
rect 222568 153824 222620 153876
rect 233332 153824 233384 153876
rect 297088 153824 297140 153876
rect 309968 153824 310020 153876
rect 355508 153824 355560 153876
rect 357348 153824 357400 153876
rect 391480 153960 391532 154012
rect 391848 153960 391900 154012
rect 417148 153960 417200 154012
rect 425244 153960 425296 154012
rect 443460 153960 443512 154012
rect 361028 153892 361080 153944
rect 376576 153892 376628 153944
rect 380808 153892 380860 153944
rect 409420 153892 409472 153944
rect 417516 153892 417568 153944
rect 63408 153756 63460 153808
rect 118700 153756 118752 153808
rect 119804 153756 119856 153808
rect 208400 153756 208452 153808
rect 244280 153756 244332 153808
rect 305368 153756 305420 153808
rect 305460 153756 305512 153808
rect 336188 153756 336240 153808
rect 355324 153756 355376 153808
rect 390192 153824 390244 153876
rect 391756 153824 391808 153876
rect 417792 153824 417844 153876
rect 418436 153892 418488 153944
rect 438308 153892 438360 153944
rect 440240 153892 440292 153944
rect 455052 153892 455104 153944
rect 437664 153824 437716 153876
rect 453948 153824 454000 153876
rect 462044 153824 462096 153876
rect 438584 153756 438636 153808
rect 453764 153756 453816 153808
rect 77208 153688 77260 153740
rect 121736 153688 121788 153740
rect 122656 153688 122708 153740
rect 212264 153688 212316 153740
rect 263600 153688 263652 153740
rect 263784 153688 263836 153740
rect 274640 153688 274692 153740
rect 310520 153688 310572 153740
rect 128360 153620 128412 153672
rect 159640 153620 159692 153672
rect 208492 153620 208544 153672
rect 273904 153620 273956 153672
rect 279884 153620 279936 153672
rect 315672 153620 315724 153672
rect 168564 153552 168616 153604
rect 216220 153552 216272 153604
rect 296812 153552 296864 153604
rect 325976 153552 326028 153604
rect 197360 153484 197412 153536
rect 237840 153484 237892 153536
rect 237472 153212 237524 153264
rect 240600 153212 240652 153264
rect 455328 153212 455380 153264
rect 463332 153212 463384 153264
rect 118700 153144 118752 153196
rect 167368 153144 167420 153196
rect 167736 153144 167788 153196
rect 246948 153144 247000 153196
rect 247224 153144 247276 153196
rect 259828 153144 259880 153196
rect 268936 153144 268988 153196
rect 280344 153144 280396 153196
rect 281172 153144 281224 153196
rect 290648 153144 290700 153196
rect 291108 153144 291160 153196
rect 334348 153144 334400 153196
rect 338948 153144 339000 153196
rect 63500 153076 63552 153128
rect 144920 153076 144972 153128
rect 155960 153076 156012 153128
rect 158352 153076 158404 153128
rect 161388 153076 161440 153128
rect 241888 153076 241940 153128
rect 245660 153076 245712 153128
rect 288072 153076 288124 153128
rect 292304 153076 292356 153128
rect 339408 153076 339460 153128
rect 355692 153144 355744 153196
rect 357440 153144 357492 153196
rect 368572 153144 368624 153196
rect 372804 153144 372856 153196
rect 385960 153144 386012 153196
rect 388260 153144 388312 153196
rect 408500 153144 408552 153196
rect 410708 153144 410760 153196
rect 435824 153144 435876 153196
rect 439596 153144 439648 153196
rect 447140 153144 447192 153196
rect 449256 153144 449308 153196
rect 452476 153144 452528 153196
rect 460664 153144 460716 153196
rect 498292 153144 498344 153196
rect 499304 153144 499356 153196
rect 505836 153144 505888 153196
rect 506756 153144 506808 153196
rect 509700 153144 509752 153196
rect 511724 153144 511776 153196
rect 512276 153144 512328 153196
rect 514852 153144 514904 153196
rect 374736 153076 374788 153128
rect 465540 153076 465592 153128
rect 474280 153076 474332 153128
rect 506388 153076 506440 153128
rect 507584 153076 507636 153128
rect 510988 153076 511040 153128
rect 513472 153076 513524 153128
rect 514208 153076 514260 153128
rect 517612 153076 517664 153128
rect 109040 153008 109092 153060
rect 198004 153008 198056 153060
rect 198096 153008 198148 153060
rect 216772 153008 216824 153060
rect 216864 153008 216916 153060
rect 239312 153008 239364 153060
rect 239956 153008 240008 153060
rect 293224 153008 293276 153060
rect 299388 153008 299440 153060
rect 306012 153008 306064 153060
rect 318708 153008 318760 153060
rect 360016 153008 360068 153060
rect 409972 153008 410024 153060
rect 431868 153008 431920 153060
rect 462136 153008 462188 153060
rect 471704 153008 471756 153060
rect 512920 153008 512972 153060
rect 515956 153008 516008 153060
rect 117228 152940 117280 152992
rect 208492 152940 208544 152992
rect 212632 152940 212684 152992
rect 267556 152940 267608 152992
rect 271696 152940 271748 152992
rect 324044 152940 324096 152992
rect 337752 152940 337804 152992
rect 375380 152940 375432 152992
rect 389088 152940 389140 152992
rect 413284 152940 413336 152992
rect 415860 152940 415912 152992
rect 436376 152940 436428 152992
rect 454592 152940 454644 152992
rect 113916 152872 113968 152924
rect 205916 152872 205968 152924
rect 210884 152872 210936 152924
rect 262404 152872 262456 152924
rect 263508 152872 263560 152924
rect 318892 152872 318944 152924
rect 328276 152872 328328 152924
rect 369584 152872 369636 152924
rect 372620 152872 372672 152924
rect 380532 152872 380584 152924
rect 380992 152872 381044 152924
rect 408132 152872 408184 152924
rect 412548 152872 412600 152924
rect 433800 152872 433852 152924
rect 452844 152872 452896 152924
rect 107476 152804 107528 152856
rect 200764 152804 200816 152856
rect 207112 152804 207164 152856
rect 212908 152804 212960 152856
rect 221740 152804 221792 152856
rect 224500 152804 224552 152856
rect 224592 152804 224644 152856
rect 244372 152804 244424 152856
rect 244556 152804 244608 152856
rect 303528 152804 303580 152856
rect 305000 152804 305052 152856
rect 316316 152804 316368 152856
rect 322756 152804 322808 152856
rect 365168 152804 365220 152856
rect 374276 152804 374328 152856
rect 402980 152804 403032 152856
rect 403256 152804 403308 152856
rect 426808 152804 426860 152856
rect 97080 152736 97132 152788
rect 193036 152736 193088 152788
rect 193128 152736 193180 152788
rect 229008 152736 229060 152788
rect 230388 152736 230440 152788
rect 249524 152736 249576 152788
rect 249616 152736 249668 152788
rect 308588 152736 308640 152788
rect 309048 152736 309100 152788
rect 354864 152736 354916 152788
rect 358912 152736 358964 152788
rect 390836 152736 390888 152788
rect 391572 152736 391624 152788
rect 416504 152736 416556 152788
rect 416688 152736 416740 152788
rect 437020 152736 437072 152788
rect 444288 152736 444340 152788
rect 453120 152736 453172 152788
rect 455420 152736 455472 152788
rect 460848 152940 460900 152992
rect 470324 152940 470376 152992
rect 514852 152940 514904 152992
rect 518532 152940 518584 152992
rect 457076 152872 457128 152924
rect 467840 152872 467892 152924
rect 469128 152872 469180 152924
rect 476856 152872 476908 152924
rect 465908 152804 465960 152856
rect 469680 152804 469732 152856
rect 477500 152804 477552 152856
rect 510344 152804 510396 152856
rect 512000 152804 512052 152856
rect 518072 152804 518124 152856
rect 522672 152804 522724 152856
rect 90364 152668 90416 152720
rect 187884 152668 187936 152720
rect 201868 152668 201920 152720
rect 221924 152668 221976 152720
rect 223948 152668 224000 152720
rect 282920 152668 282972 152720
rect 284392 152668 284444 152720
rect 295800 152668 295852 152720
rect 295892 152668 295944 152720
rect 344560 152668 344612 152720
rect 362960 152668 363012 152720
rect 395988 152668 396040 152720
rect 396632 152668 396684 152720
rect 421656 152668 421708 152720
rect 445484 152668 445536 152720
rect 455696 152668 455748 152720
rect 464620 152736 464672 152788
rect 467196 152736 467248 152788
rect 475568 152736 475620 152788
rect 466552 152668 466604 152720
rect 468024 152668 468076 152720
rect 476212 152668 476264 152720
rect 73528 152600 73580 152652
rect 175096 152600 175148 152652
rect 212356 152600 212408 152652
rect 272708 152600 272760 152652
rect 278688 152600 278740 152652
rect 329196 152600 329248 152652
rect 329288 152600 329340 152652
rect 370228 152600 370280 152652
rect 376668 152600 376720 152652
rect 406200 152600 406252 152652
rect 406936 152600 406988 152652
rect 428648 152600 428700 152652
rect 450360 152600 450412 152652
rect 462688 152600 462740 152652
rect 462964 152600 463016 152652
rect 472348 152600 472400 152652
rect 518808 152600 518860 152652
rect 523500 152600 523552 152652
rect 23388 152532 23440 152584
rect 136548 152532 136600 152584
rect 147588 152532 147640 152584
rect 231584 152532 231636 152584
rect 242440 152532 242492 152584
rect 254676 152532 254728 152584
rect 255228 152532 255280 152584
rect 313740 152532 313792 152584
rect 314936 152532 314988 152584
rect 359372 152532 359424 152584
rect 365444 152532 365496 152584
rect 397828 152532 397880 152584
rect 399024 152532 399076 152584
rect 423588 152532 423640 152584
rect 446956 152532 447008 152584
rect 460112 152532 460164 152584
rect 6276 152464 6328 152516
rect 123668 152464 123720 152516
rect 125692 152464 125744 152516
rect 127532 152464 127584 152516
rect 134064 152464 134116 152516
rect 221280 152464 221332 152516
rect 222016 152464 222068 152516
rect 224592 152464 224644 152516
rect 234988 152464 235040 152516
rect 298376 152464 298428 152516
rect 302332 152464 302384 152516
rect 349712 152464 349764 152516
rect 109132 152396 109184 152448
rect 122380 152396 122432 152448
rect 124128 152396 124180 152448
rect 128820 152396 128872 152448
rect 129832 152396 129884 152448
rect 139124 152396 139176 152448
rect 143080 152396 143132 152448
rect 216128 152396 216180 152448
rect 216220 152396 216272 152448
rect 247592 152396 247644 152448
rect 256700 152396 256752 152448
rect 301596 152396 301648 152448
rect 301688 152396 301740 152448
rect 311164 152396 311216 152448
rect 144828 152328 144880 152380
rect 209136 152328 209188 152380
rect 230756 152328 230808 152380
rect 257252 152328 257304 152380
rect 260748 152328 260800 152380
rect 270132 152328 270184 152380
rect 272524 152328 272576 152380
rect 285496 152328 285548 152380
rect 109224 152260 109276 152312
rect 157064 152260 157116 152312
rect 157340 152260 157392 152312
rect 160928 152260 160980 152312
rect 174912 152260 174964 152312
rect 226432 152260 226484 152312
rect 256792 152260 256844 152312
rect 264980 152260 265032 152312
rect 265072 152260 265124 152312
rect 275284 152260 275336 152312
rect 288256 152260 288308 152312
rect 300952 152260 301004 152312
rect 311072 152260 311124 152312
rect 321468 152396 321520 152448
rect 349436 152396 349488 152448
rect 385592 152464 385644 152516
rect 392308 152464 392360 152516
rect 418436 152464 418488 152516
rect 437388 152464 437440 152516
rect 452476 152464 452528 152516
rect 459652 152464 459704 152516
rect 469772 152532 469824 152584
rect 470508 152532 470560 152584
rect 478144 152532 478196 152584
rect 414296 152396 414348 152448
rect 415860 152396 415912 152448
rect 452016 152396 452068 152448
rect 463976 152464 464028 152516
rect 464988 152464 465040 152516
rect 473636 152464 473688 152516
rect 517428 152464 517480 152516
rect 521844 152464 521896 152516
rect 507124 152328 507176 152380
rect 507860 152328 507912 152380
rect 511632 152328 511684 152380
rect 513564 152328 513616 152380
rect 54208 152192 54260 152244
rect 89168 152192 89220 152244
rect 204168 152192 204220 152244
rect 252100 152192 252152 152244
rect 513564 152192 513616 152244
rect 516140 152192 516192 152244
rect 23296 152124 23348 152176
rect 110052 152124 110104 152176
rect 71412 152056 71464 152108
rect 82820 152056 82872 152108
rect 95516 152056 95568 152108
rect 114376 152056 114428 152108
rect 88616 151988 88668 152040
rect 110144 151988 110196 152040
rect 515496 151988 515548 152040
rect 518992 151988 519044 152040
rect 33600 151920 33652 151972
rect 110236 151920 110288 151972
rect 138020 151920 138072 151972
rect 144276 151920 144328 151972
rect 507768 151920 507820 151972
rect 509240 151920 509292 151972
rect 516784 151920 516836 151972
rect 520280 151920 520332 151972
rect 26700 151852 26752 151904
rect 109776 151852 109828 151904
rect 127624 151852 127676 151904
rect 133972 151852 134024 151904
rect 139492 151852 139544 151904
rect 142988 151852 143040 151904
rect 194324 151852 194376 151904
rect 202696 151852 202748 151904
rect 320732 151852 320784 151904
rect 326620 151852 326672 151904
rect 332600 151852 332652 151904
rect 336832 151852 336884 151904
rect 343640 151852 343692 151904
rect 347136 151852 347188 151904
rect 359464 151852 359516 151904
rect 364524 151852 364576 151904
rect 508412 151852 508464 151904
rect 510068 151852 510120 151904
rect 81716 151784 81768 151836
rect 97724 151784 97776 151836
rect 102324 151784 102376 151836
rect 110328 151784 110380 151836
rect 208400 151784 208452 151836
rect 210424 151784 210476 151836
rect 509056 151784 509108 151836
rect 510896 151784 510948 151836
rect 516048 151784 516100 151836
rect 520188 151784 520240 151836
rect 132408 151716 132460 151768
rect 219348 151716 219400 151768
rect 122748 151648 122800 151700
rect 211620 151648 211672 151700
rect 111708 151580 111760 151632
rect 203984 151580 204036 151632
rect 104808 151512 104860 151564
rect 198832 151512 198884 151564
rect 212448 151512 212500 151564
rect 280988 151512 281040 151564
rect 97908 151444 97960 151496
rect 193680 151444 193732 151496
rect 202788 151444 202840 151496
rect 273260 151444 273312 151496
rect 92388 151376 92440 151428
rect 188528 151376 188580 151428
rect 195888 151376 195940 151428
rect 268200 151376 268252 151428
rect 78588 151308 78640 151360
rect 178316 151308 178368 151360
rect 180708 151308 180760 151360
rect 256608 151308 256660 151360
rect 64788 151240 64840 151292
rect 57888 151172 57940 151224
rect 162860 151172 162912 151224
rect 167644 151240 167696 151292
rect 245016 151240 245068 151292
rect 168012 151172 168064 151224
rect 168104 151172 168156 151224
rect 246304 151172 246356 151224
rect 50988 151104 51040 151156
rect 157708 151104 157760 151156
rect 158628 151104 158680 151156
rect 239956 151104 240008 151156
rect 38568 151036 38620 151088
rect 147496 151036 147548 151088
rect 151728 151036 151780 151088
rect 234804 151036 234856 151088
rect 146208 150968 146260 151020
rect 229652 150968 229704 151020
rect 153108 150900 153160 150952
rect 235448 150900 235500 150952
rect 166908 150832 166960 150884
rect 168104 150832 168156 150884
rect 105820 150628 105872 150680
rect 116032 150628 116084 150680
rect 98920 150560 98972 150612
rect 114468 150560 114520 150612
rect 92020 150492 92072 150544
rect 114008 150492 114060 150544
rect 85212 150424 85264 150476
rect 117044 150424 117096 150476
rect 127072 150152 127124 150204
rect 128222 150152 128274 150204
rect 132500 150152 132552 150204
rect 133374 150152 133426 150204
rect 139400 150152 139452 150204
rect 140458 150152 140510 150204
rect 145104 150152 145156 150204
rect 146254 150152 146306 150204
rect 147680 150152 147732 150204
rect 148830 150152 148882 150204
rect 149152 150152 149204 150204
rect 150026 150152 150078 150204
rect 150532 150152 150584 150204
rect 151314 150152 151366 150204
rect 154672 150152 154724 150204
rect 155822 150152 155874 150204
rect 161480 150152 161532 150204
rect 162262 150152 162314 150204
rect 163044 150152 163096 150204
rect 164194 150152 164246 150204
rect 168380 150152 168432 150204
rect 169346 150152 169398 150204
rect 169852 150152 169904 150204
rect 170634 150152 170686 150204
rect 171140 150152 171192 150204
rect 171922 150152 171974 150204
rect 172704 150152 172756 150204
rect 173854 150152 173906 150204
rect 179420 150152 179472 150204
rect 180294 150152 180346 150204
rect 180984 150152 181036 150204
rect 182134 150152 182186 150204
rect 183560 150152 183612 150204
rect 184710 150152 184762 150204
rect 190736 150152 190788 150204
rect 191794 150152 191846 150204
rect 194600 150152 194652 150204
rect 195658 150152 195710 150204
rect 200304 150152 200356 150204
rect 201454 150152 201506 150204
rect 209964 150152 210016 150204
rect 211114 150152 211166 150204
rect 224960 150152 225012 150204
rect 225834 150152 225886 150204
rect 229192 150152 229244 150204
rect 230342 150152 230394 150204
rect 233240 150152 233292 150204
rect 234206 150152 234258 150204
rect 240140 150152 240192 150204
rect 241290 150152 241342 150204
rect 242900 150152 242952 150204
rect 243774 150152 243826 150204
rect 247132 150152 247184 150204
rect 248282 150152 248334 150204
rect 252560 150152 252612 150204
rect 253434 150152 253486 150204
rect 258080 150152 258132 150204
rect 259230 150152 259282 150204
rect 260840 150152 260892 150204
rect 261806 150152 261858 150204
rect 263600 150152 263652 150204
rect 264382 150152 264434 150204
rect 265164 150152 265216 150204
rect 266314 150152 266366 150204
rect 273444 150152 273496 150204
rect 274594 150152 274646 150204
rect 276020 150152 276072 150204
rect 277170 150152 277222 150204
rect 283104 150152 283156 150204
rect 284254 150152 284306 150204
rect 291200 150152 291252 150204
rect 291982 150152 292034 150204
rect 292764 150152 292816 150204
rect 293914 150152 293966 150204
rect 299480 150152 299532 150204
rect 300354 150152 300406 150204
rect 310612 150152 310664 150204
rect 311854 150152 311906 150204
rect 311992 150152 312044 150204
rect 313142 150152 313194 150204
rect 330024 150152 330076 150204
rect 331174 150152 331226 150204
rect 331312 150152 331364 150204
rect 332462 150152 332514 150204
rect 339592 150152 339644 150204
rect 340742 150152 340794 150204
rect 349252 150152 349304 150204
rect 350402 150152 350454 150204
rect 350540 150152 350592 150204
rect 351690 150152 351742 150204
rect 351920 150152 351972 150204
rect 352978 150152 353030 150204
rect 357624 150152 357676 150204
rect 358774 150152 358826 150204
rect 360200 150152 360252 150204
rect 361350 150152 361402 150204
rect 361580 150152 361632 150204
rect 362638 150152 362690 150204
rect 365904 150152 365956 150204
rect 367054 150152 367106 150204
rect 383660 150152 383712 150204
rect 384442 150152 384494 150204
rect 385224 150152 385276 150204
rect 386374 150152 386426 150204
rect 386512 150152 386564 150204
rect 387662 150152 387714 150204
rect 391940 150152 391992 150204
rect 392814 150152 392866 150204
rect 396172 150152 396224 150204
rect 397230 150152 397282 150204
rect 400220 150152 400272 150204
rect 401094 150152 401146 150204
rect 412824 150152 412876 150204
rect 413974 150152 414026 150204
rect 423772 150152 423824 150204
rect 424922 150152 424974 150204
rect 434720 150152 434772 150204
rect 435778 150152 435830 150204
rect 441712 150152 441764 150204
rect 442862 150152 442914 150204
rect 443000 150152 443052 150204
rect 444150 150152 444202 150204
rect 444380 150152 444432 150204
rect 445438 150152 445490 150204
rect 456800 150152 456852 150204
rect 457674 150152 457726 150204
rect 477684 150152 477736 150204
rect 478834 150152 478886 150204
rect 478972 150152 479024 150204
rect 480122 150152 480174 150204
rect 483020 150152 483072 150204
rect 483986 150152 484038 150204
rect 485780 150152 485832 150204
rect 486562 150152 486614 150204
rect 488632 150152 488684 150204
rect 489690 150152 489742 150204
rect 489920 150152 489972 150204
rect 490978 150152 491030 150204
rect 491300 150152 491352 150204
rect 492266 150152 492318 150204
rect 97724 149880 97776 149932
rect 116492 149880 116544 149932
rect 89168 149812 89220 149864
rect 116216 149812 116268 149864
rect 82820 149744 82872 149796
rect 117136 149744 117188 149796
rect 78588 149676 78640 149728
rect 112812 149676 112864 149728
rect 75184 149608 75236 149660
rect 114192 149608 114244 149660
rect 68376 149540 68428 149592
rect 112720 149540 112772 149592
rect 64696 149472 64748 149524
rect 111248 149472 111300 149524
rect 61384 149404 61436 149456
rect 112628 149404 112680 149456
rect 57888 149336 57940 149388
rect 112536 149336 112588 149388
rect 40776 149268 40828 149320
rect 44088 149268 44140 149320
rect 47584 149268 47636 149320
rect 50988 149268 51040 149320
rect 112444 149268 112496 149320
rect 111156 149200 111208 149252
rect 111064 149132 111116 149184
rect 109684 149064 109736 149116
rect 109592 148996 109644 149048
rect 116124 148996 116176 149048
rect 110328 147024 110380 147076
rect 116124 147024 116176 147076
rect 110052 146956 110104 147008
rect 116860 146956 116912 147008
rect 110236 146888 110288 146940
rect 116952 146888 117004 146940
rect 110144 145528 110196 145580
rect 116400 145528 116452 145580
rect 113732 143556 113784 143608
rect 115204 143556 115256 143608
rect 114468 143488 114520 143540
rect 115940 143488 115992 143540
rect 114376 141720 114428 141772
rect 115940 141720 115992 141772
rect 114008 140700 114060 140752
rect 115940 140700 115992 140752
rect 109776 134512 109828 134564
rect 117044 134512 117096 134564
rect 112812 132404 112864 132456
rect 116124 132404 116176 132456
rect 114192 131044 114244 131096
rect 115940 131044 115992 131096
rect 112720 126896 112772 126948
rect 116124 126896 116176 126948
rect 111248 124108 111300 124160
rect 116124 124108 116176 124160
rect 112628 122748 112680 122800
rect 115940 122748 115992 122800
rect 112536 121388 112588 121440
rect 115940 121388 115992 121440
rect 114192 118804 114244 118856
rect 115296 118804 115348 118856
rect 112444 117240 112496 117292
rect 116032 117240 116084 117292
rect 111156 114452 111208 114504
rect 116124 114452 116176 114504
rect 111064 113092 111116 113144
rect 116124 113092 116176 113144
rect 109684 111732 109736 111784
rect 116124 111732 116176 111784
rect 113548 109556 113600 109608
rect 115388 109556 115440 109608
rect 114284 108944 114336 108996
rect 116400 108944 116452 108996
rect 114100 104796 114152 104848
rect 115940 104796 115992 104848
rect 114468 96840 114520 96892
rect 116768 96840 116820 96892
rect 113824 93576 113876 93628
rect 116492 93576 116544 93628
rect 113916 92420 113968 92472
rect 116124 92420 116176 92472
rect 115204 91604 115256 91656
rect 116860 91604 116912 91656
rect 114468 87184 114520 87236
rect 116676 87184 116728 87236
rect 114008 86912 114060 86964
rect 116216 86912 116268 86964
rect 113824 71748 113876 71800
rect 116400 71748 116452 71800
rect 114100 69028 114152 69080
rect 116308 69028 116360 69080
rect 114192 67600 114244 67652
rect 116216 67600 116268 67652
rect 114468 64676 114520 64728
rect 116584 64676 116636 64728
rect 112444 62092 112496 62144
rect 116124 62092 116176 62144
rect 111064 59372 111116 59424
rect 116124 59372 116176 59424
rect 113824 51076 113876 51128
rect 115940 51076 115992 51128
rect 114284 48220 114336 48272
rect 116860 48220 116912 48272
rect 113916 46928 113968 46980
rect 116032 46928 116084 46980
rect 114008 42780 114060 42832
rect 116400 42780 116452 42832
rect 114100 38632 114152 38684
rect 115940 38632 115992 38684
rect 109684 37272 109736 37324
rect 116124 37272 116176 37324
rect 109776 33124 109828 33176
rect 116124 33124 116176 33176
rect 116308 31016 116360 31068
rect 117228 31016 117280 31068
rect 112536 27616 112588 27668
rect 116124 27616 116176 27668
rect 112628 23468 112680 23520
rect 116124 23468 116176 23520
rect 111248 22788 111300 22840
rect 117044 22788 117096 22840
rect 111156 22720 111208 22772
rect 116308 22720 116360 22772
rect 112720 22108 112772 22160
rect 116124 22108 116176 22160
rect 111340 19320 111392 19372
rect 116124 19320 116176 19372
rect 111432 17960 111484 18012
rect 116124 17960 116176 18012
rect 111616 15172 111668 15224
rect 116124 15172 116176 15224
rect 114284 13812 114336 13864
rect 115940 13812 115992 13864
rect 114192 7964 114244 8016
rect 115204 7964 115256 8016
rect 109868 4836 109920 4888
rect 116952 4836 117004 4888
rect 109960 4768 110012 4820
rect 117228 4768 117280 4820
rect 109592 4496 109644 4548
rect 112444 4496 112496 4548
rect 2504 2796 2556 2848
rect 32772 2592 32824 2644
rect 111524 3000 111576 3052
rect 118700 2932 118752 2984
rect 116124 2796 116176 2848
rect 98276 2592 98328 2644
rect 106188 2592 106240 2644
rect 111064 2592 111116 2644
rect 93032 2116 93084 2168
rect 116676 2116 116728 2168
rect 86408 2048 86460 2100
rect 116768 2048 116820 2100
rect 79600 1980 79652 2032
rect 116860 1980 116912 2032
rect 72700 1912 72752 1964
rect 109868 1912 109920 1964
rect 65984 1844 66036 1896
rect 109684 1844 109736 1896
rect 59360 1776 59412 1828
rect 109776 1776 109828 1828
rect 52644 1708 52696 1760
rect 116492 1708 116544 1760
rect 46020 1640 46072 1692
rect 112536 1640 112588 1692
rect 49332 1572 49384 1624
rect 116400 1572 116452 1624
rect 32680 1504 32732 1556
rect 111340 1504 111392 1556
rect 12624 1436 12676 1488
rect 98000 1436 98052 1488
rect 99380 1436 99432 1488
rect 111156 1436 111208 1488
rect 118700 1436 118752 1488
rect 143632 1436 143684 1488
rect 394240 1436 394292 1488
rect 425796 1436 425848 1488
rect 444288 1436 444340 1488
rect 491300 1436 491352 1488
rect 9312 1368 9364 1420
rect 100760 1368 100812 1420
rect 102692 1368 102744 1420
rect 111248 1368 111300 1420
rect 111524 1368 111576 1420
rect 193588 1368 193640 1420
rect 193680 1368 193732 1420
rect 243636 1368 243688 1420
rect 243728 1368 243780 1420
rect 293592 1368 293644 1420
rect 295340 1368 295392 1420
rect 493600 1368 493652 1420
rect 95976 1300 96028 1352
rect 116584 1300 116636 1352
rect 35992 1232 36044 1284
rect 112720 1232 112772 1284
rect 39304 1164 39356 1216
rect 112628 1164 112680 1216
rect 62672 1096 62724 1148
rect 117136 1096 117188 1148
rect 69296 1028 69348 1080
rect 114100 1028 114152 1080
rect 76012 960 76064 1012
rect 114008 960 114060 1012
rect 82636 892 82688 944
rect 113916 892 113968 944
rect 89352 824 89404 876
rect 113824 824 113876 876
rect 22652 756 22704 808
rect 114192 756 114244 808
<< metal2 >>
rect 386 163200 442 164400
rect 1214 163200 1270 164400
rect 2042 163200 2098 164400
rect 2870 163200 2926 164400
rect 3698 163200 3754 164400
rect 4526 163200 4582 164400
rect 5354 163200 5410 164400
rect 6274 163200 6330 164400
rect 7102 163200 7158 164400
rect 7930 163200 7986 164400
rect 8758 163200 8814 164400
rect 9586 163200 9642 164400
rect 10414 163200 10470 164400
rect 11242 163200 11298 164400
rect 12162 163200 12218 164400
rect 12990 163200 13046 164400
rect 13818 163200 13874 164400
rect 14646 163200 14702 164400
rect 15474 163200 15530 164400
rect 16302 163200 16358 164400
rect 17130 163200 17186 164400
rect 18050 163200 18106 164400
rect 18878 163200 18934 164400
rect 19706 163200 19762 164400
rect 20534 163200 20590 164400
rect 21362 163200 21418 164400
rect 22190 163200 22246 164400
rect 23018 163200 23074 164400
rect 23124 163254 23428 163282
rect 400 158778 428 163200
rect 388 158772 440 158778
rect 388 158714 440 158720
rect 1228 155242 1256 163200
rect 2056 161474 2084 163200
rect 2056 161446 2176 161474
rect 2044 158772 2096 158778
rect 2044 158714 2096 158720
rect 1216 155236 1268 155242
rect 1216 155178 1268 155184
rect 2056 151065 2084 158714
rect 2148 158030 2176 161446
rect 2884 159526 2912 163200
rect 3712 159662 3740 163200
rect 3700 159656 3752 159662
rect 3700 159598 3752 159604
rect 2872 159520 2924 159526
rect 2872 159462 2924 159468
rect 2136 158024 2188 158030
rect 2136 157966 2188 157972
rect 4540 157214 4568 163200
rect 4528 157208 4580 157214
rect 4528 157150 4580 157156
rect 5368 155281 5396 163200
rect 5354 155272 5410 155281
rect 5354 155207 5410 155216
rect 6288 152522 6316 163200
rect 7116 153785 7144 163200
rect 7944 156641 7972 163200
rect 7930 156632 7986 156641
rect 7930 156567 7986 156576
rect 8772 155310 8800 163200
rect 8760 155304 8812 155310
rect 8760 155246 8812 155252
rect 7102 153776 7158 153785
rect 7102 153711 7158 153720
rect 6276 152516 6328 152522
rect 6276 152458 6328 152464
rect 9600 152425 9628 163200
rect 10428 153921 10456 163200
rect 11256 156738 11284 163200
rect 12176 158001 12204 163200
rect 13004 159390 13032 163200
rect 12992 159384 13044 159390
rect 12992 159326 13044 159332
rect 12162 157992 12218 158001
rect 12162 157927 12218 157936
rect 11244 156732 11296 156738
rect 11244 156674 11296 156680
rect 10414 153912 10470 153921
rect 13832 153882 13860 163200
rect 14660 156670 14688 163200
rect 14648 156664 14700 156670
rect 14648 156606 14700 156612
rect 15488 155378 15516 163200
rect 15476 155372 15528 155378
rect 15476 155314 15528 155320
rect 10414 153847 10470 153856
rect 13820 153876 13872 153882
rect 13820 153818 13872 153824
rect 16316 152561 16344 163200
rect 17144 153950 17172 163200
rect 18064 156806 18092 163200
rect 18892 158098 18920 163200
rect 19720 159361 19748 163200
rect 19706 159352 19762 159361
rect 19706 159287 19762 159296
rect 18880 158092 18932 158098
rect 18880 158034 18932 158040
rect 18052 156800 18104 156806
rect 18052 156742 18104 156748
rect 20548 154018 20576 163200
rect 21376 156777 21404 163200
rect 21362 156768 21418 156777
rect 21362 156703 21418 156712
rect 22204 155446 22232 163200
rect 23032 163146 23060 163200
rect 23124 163146 23152 163254
rect 23032 163118 23152 163146
rect 22192 155440 22244 155446
rect 22192 155382 22244 155388
rect 20536 154012 20588 154018
rect 20536 153954 20588 153960
rect 17132 153944 17184 153950
rect 17132 153886 17184 153892
rect 23400 152590 23428 163254
rect 23938 163200 23994 164400
rect 24766 163200 24822 164400
rect 25594 163200 25650 164400
rect 26422 163200 26478 164400
rect 27250 163200 27306 164400
rect 28078 163200 28134 164400
rect 28906 163200 28962 164400
rect 29826 163200 29882 164400
rect 30654 163200 30710 164400
rect 31482 163200 31538 164400
rect 32310 163200 32366 164400
rect 33138 163200 33194 164400
rect 33966 163200 34022 164400
rect 34794 163200 34850 164400
rect 35714 163200 35770 164400
rect 36542 163200 36598 164400
rect 37370 163200 37426 164400
rect 38198 163200 38254 164400
rect 38304 163254 38516 163282
rect 23952 155514 23980 163200
rect 24780 156874 24808 163200
rect 24768 156868 24820 156874
rect 24768 156810 24820 156816
rect 23940 155508 23992 155514
rect 23940 155450 23992 155456
rect 25608 154086 25636 163200
rect 26436 159458 26464 163200
rect 26424 159452 26476 159458
rect 26424 159394 26476 159400
rect 27264 155417 27292 163200
rect 28092 156942 28120 163200
rect 28080 156936 28132 156942
rect 28080 156878 28132 156884
rect 27250 155408 27306 155417
rect 27250 155343 27306 155352
rect 25596 154080 25648 154086
rect 25596 154022 25648 154028
rect 23388 152584 23440 152590
rect 16302 152552 16358 152561
rect 23388 152526 23440 152532
rect 16302 152487 16358 152496
rect 9586 152416 9642 152425
rect 9586 152351 9642 152360
rect 23296 152176 23348 152182
rect 12990 152144 13046 152153
rect 23296 152118 23348 152124
rect 12990 152079 13046 152088
rect 9494 152008 9550 152017
rect 9494 151943 9550 151952
rect 2686 151872 2742 151881
rect 2686 151807 2742 151816
rect 2042 151056 2098 151065
rect 2042 150991 2098 151000
rect 2700 149940 2728 151807
rect 9508 149940 9536 151943
rect 13004 149940 13032 152079
rect 23308 149940 23336 152118
rect 26700 151904 26752 151910
rect 26700 151846 26752 151852
rect 26712 149940 26740 151846
rect 28920 151201 28948 163200
rect 29840 158506 29868 163200
rect 29828 158500 29880 158506
rect 29828 158442 29880 158448
rect 30668 155553 30696 163200
rect 31496 158234 31524 163200
rect 31484 158228 31536 158234
rect 31484 158170 31536 158176
rect 32324 158166 32352 163200
rect 33152 159497 33180 163200
rect 33980 159594 34008 163200
rect 33968 159588 34020 159594
rect 33968 159530 34020 159536
rect 33138 159488 33194 159497
rect 33138 159423 33194 159432
rect 32312 158160 32364 158166
rect 32312 158102 32364 158108
rect 30654 155544 30710 155553
rect 30654 155479 30710 155488
rect 34808 154154 34836 163200
rect 35728 158137 35756 163200
rect 36556 160750 36584 163200
rect 36544 160744 36596 160750
rect 36544 160686 36596 160692
rect 37384 159186 37412 163200
rect 38212 163146 38240 163200
rect 38304 163146 38332 163254
rect 38212 163118 38332 163146
rect 37372 159180 37424 159186
rect 37372 159122 37424 159128
rect 35714 158128 35770 158137
rect 35714 158063 35770 158072
rect 34796 154148 34848 154154
rect 34796 154090 34848 154096
rect 38488 154057 38516 163254
rect 39026 163200 39082 164400
rect 39854 163200 39910 164400
rect 40682 163200 40738 164400
rect 41602 163200 41658 164400
rect 42430 163200 42486 164400
rect 43258 163200 43314 164400
rect 44086 163200 44142 164400
rect 44914 163200 44970 164400
rect 45742 163200 45798 164400
rect 46570 163200 46626 164400
rect 47490 163200 47546 164400
rect 48318 163200 48374 164400
rect 49146 163200 49202 164400
rect 49974 163200 50030 164400
rect 50802 163200 50858 164400
rect 51630 163200 51686 164400
rect 52458 163200 52514 164400
rect 53378 163200 53434 164400
rect 54206 163200 54262 164400
rect 55034 163200 55090 164400
rect 55862 163200 55918 164400
rect 56690 163200 56746 164400
rect 57518 163200 57574 164400
rect 57624 163254 57928 163282
rect 38568 159180 38620 159186
rect 38568 159122 38620 159128
rect 38474 154048 38530 154057
rect 38474 153983 38530 153992
rect 33600 151972 33652 151978
rect 33600 151914 33652 151920
rect 28906 151192 28962 151201
rect 28906 151127 28962 151136
rect 30194 150512 30250 150521
rect 30194 150447 30250 150456
rect 30208 149940 30236 150447
rect 33612 149940 33640 151914
rect 38580 151094 38608 159122
rect 39040 157010 39068 163200
rect 39868 162586 39896 163200
rect 39856 162580 39908 162586
rect 39856 162522 39908 162528
rect 40696 160818 40724 163200
rect 40684 160812 40736 160818
rect 40684 160754 40736 160760
rect 39028 157004 39080 157010
rect 39028 156946 39080 156952
rect 41616 155582 41644 163200
rect 42444 158302 42472 163200
rect 43272 162654 43300 163200
rect 43260 162648 43312 162654
rect 43260 162590 43312 162596
rect 42432 158296 42484 158302
rect 42432 158238 42484 158244
rect 41604 155576 41656 155582
rect 41604 155518 41656 155524
rect 44100 151337 44128 163200
rect 44928 154222 44956 163200
rect 45756 158370 45784 163200
rect 46584 159798 46612 163200
rect 47504 160886 47532 163200
rect 47492 160880 47544 160886
rect 47492 160822 47544 160828
rect 46572 159792 46624 159798
rect 46572 159734 46624 159740
rect 45744 158364 45796 158370
rect 45744 158306 45796 158312
rect 48332 155650 48360 163200
rect 49160 157078 49188 163200
rect 49988 159322 50016 163200
rect 50816 161474 50844 163200
rect 50816 161446 51028 161474
rect 49976 159316 50028 159322
rect 49976 159258 50028 159264
rect 49148 157072 49200 157078
rect 49148 157014 49200 157020
rect 48320 155644 48372 155650
rect 48320 155586 48372 155592
rect 44916 154216 44968 154222
rect 44916 154158 44968 154164
rect 44086 151328 44142 151337
rect 44086 151263 44142 151272
rect 51000 151162 51028 161446
rect 51644 154290 51672 163200
rect 52472 158438 52500 163200
rect 53392 159730 53420 163200
rect 54220 160954 54248 163200
rect 54208 160948 54260 160954
rect 54208 160890 54260 160896
rect 53380 159724 53432 159730
rect 53380 159666 53432 159672
rect 52460 158432 52512 158438
rect 52460 158374 52512 158380
rect 55048 155718 55076 163200
rect 55772 158500 55824 158506
rect 55772 158442 55824 158448
rect 55036 155712 55088 155718
rect 55036 155654 55088 155660
rect 51632 154284 51684 154290
rect 51632 154226 51684 154232
rect 55784 152833 55812 158442
rect 55876 157146 55904 163200
rect 56704 161702 56732 163200
rect 57532 163146 57560 163200
rect 57624 163146 57652 163254
rect 57532 163118 57652 163146
rect 56692 161696 56744 161702
rect 56692 161638 56744 161644
rect 55864 157140 55916 157146
rect 55864 157082 55916 157088
rect 55770 152824 55826 152833
rect 55770 152759 55826 152768
rect 54208 152244 54260 152250
rect 54208 152186 54260 152192
rect 50988 151156 51040 151162
rect 50988 151098 51040 151104
rect 38568 151088 38620 151094
rect 38568 151030 38620 151036
rect 37002 150648 37058 150657
rect 37002 150583 37058 150592
rect 37016 149940 37044 150583
rect 54220 149940 54248 152186
rect 57900 151230 57928 163254
rect 58346 163200 58402 164400
rect 59266 163200 59322 164400
rect 60094 163200 60150 164400
rect 60922 163200 60978 164400
rect 61750 163200 61806 164400
rect 62578 163200 62634 164400
rect 63406 163200 63462 164400
rect 64234 163200 64290 164400
rect 65154 163200 65210 164400
rect 65982 163200 66038 164400
rect 66810 163200 66866 164400
rect 67638 163200 67694 164400
rect 68466 163200 68522 164400
rect 69294 163200 69350 164400
rect 70122 163200 70178 164400
rect 71042 163200 71098 164400
rect 71870 163200 71926 164400
rect 72698 163200 72754 164400
rect 73526 163200 73582 164400
rect 74354 163200 74410 164400
rect 75182 163200 75238 164400
rect 76010 163200 76066 164400
rect 76930 163200 76986 164400
rect 77758 163200 77814 164400
rect 78586 163200 78642 164400
rect 79414 163200 79470 164400
rect 80242 163200 80298 164400
rect 81070 163200 81126 164400
rect 81898 163200 81954 164400
rect 82818 163200 82874 164400
rect 83646 163200 83702 164400
rect 83752 163254 84148 163282
rect 58360 154358 58388 163200
rect 59280 158506 59308 163200
rect 60108 159633 60136 163200
rect 60936 161022 60964 163200
rect 61764 161634 61792 163200
rect 61752 161628 61804 161634
rect 61752 161570 61804 161576
rect 60924 161016 60976 161022
rect 60924 160958 60976 160964
rect 60094 159624 60150 159633
rect 60094 159559 60150 159568
rect 62592 158574 62620 163200
rect 62580 158568 62632 158574
rect 62580 158510 62632 158516
rect 59268 158500 59320 158506
rect 59268 158442 59320 158448
rect 58348 154352 58400 154358
rect 58348 154294 58400 154300
rect 63420 153814 63448 163200
rect 63500 159588 63552 159594
rect 63500 159530 63552 159536
rect 63408 153808 63460 153814
rect 63408 153750 63460 153756
rect 63512 153134 63540 159530
rect 64248 158778 64276 163200
rect 65168 161770 65196 163200
rect 65156 161764 65208 161770
rect 65156 161706 65208 161712
rect 65996 158778 66024 163200
rect 66824 159594 66852 163200
rect 67652 161090 67680 163200
rect 68480 161838 68508 163200
rect 68468 161832 68520 161838
rect 68468 161774 68520 161780
rect 67640 161084 67692 161090
rect 67640 161026 67692 161032
rect 66812 159588 66864 159594
rect 66812 159530 66864 159536
rect 64236 158772 64288 158778
rect 64236 158714 64288 158720
rect 64788 158772 64840 158778
rect 64788 158714 64840 158720
rect 65984 158772 66036 158778
rect 65984 158714 66036 158720
rect 63500 153128 63552 153134
rect 63500 153070 63552 153076
rect 64800 151298 64828 158714
rect 69308 157282 69336 163200
rect 70136 159866 70164 163200
rect 70124 159860 70176 159866
rect 70124 159802 70176 159808
rect 71056 158778 71084 163200
rect 71884 162042 71912 163200
rect 71872 162036 71924 162042
rect 71872 161978 71924 161984
rect 71044 158772 71096 158778
rect 71044 158714 71096 158720
rect 71688 158772 71740 158778
rect 71688 158714 71740 158720
rect 69296 157276 69348 157282
rect 69296 157218 69348 157224
rect 71412 152108 71464 152114
rect 71412 152050 71464 152056
rect 64788 151292 64840 151298
rect 64788 151234 64840 151240
rect 57888 151224 57940 151230
rect 57888 151166 57940 151172
rect 71424 149940 71452 152050
rect 71700 151473 71728 158714
rect 72712 155786 72740 163200
rect 72700 155780 72752 155786
rect 72700 155722 72752 155728
rect 73540 152658 73568 163200
rect 74368 160721 74396 163200
rect 75196 161906 75224 163200
rect 75184 161900 75236 161906
rect 75184 161842 75236 161848
rect 74354 160712 74410 160721
rect 74354 160647 74410 160656
rect 76024 159254 76052 163200
rect 76944 159934 76972 163200
rect 76932 159928 76984 159934
rect 76932 159870 76984 159876
rect 77208 159656 77260 159662
rect 77208 159598 77260 159604
rect 76012 159248 76064 159254
rect 76012 159190 76064 159196
rect 77220 153746 77248 159598
rect 77772 158778 77800 163200
rect 78600 161974 78628 163200
rect 78588 161968 78640 161974
rect 78588 161910 78640 161916
rect 77760 158772 77812 158778
rect 77760 158714 77812 158720
rect 78588 158772 78640 158778
rect 78588 158714 78640 158720
rect 77208 153740 77260 153746
rect 77208 153682 77260 153688
rect 73528 152652 73580 152658
rect 73528 152594 73580 152600
rect 71686 151464 71742 151473
rect 71686 151399 71742 151408
rect 78600 151366 78628 158714
rect 79428 158273 79456 163200
rect 80256 159662 80284 163200
rect 81084 161158 81112 163200
rect 81912 162110 81940 163200
rect 81900 162104 81952 162110
rect 81900 162046 81952 162052
rect 81072 161152 81124 161158
rect 81072 161094 81124 161100
rect 80244 159656 80296 159662
rect 80244 159598 80296 159604
rect 79968 159248 80020 159254
rect 79968 159190 80020 159196
rect 79414 158264 79470 158273
rect 79414 158199 79470 158208
rect 79980 157350 80008 159190
rect 79968 157344 80020 157350
rect 79968 157286 80020 157292
rect 82832 156913 82860 163200
rect 83660 163146 83688 163200
rect 83752 163146 83780 163254
rect 83660 163118 83780 163146
rect 82818 156904 82874 156913
rect 82818 156839 82874 156848
rect 84120 152697 84148 163254
rect 84474 163200 84530 164400
rect 85302 163200 85358 164400
rect 86130 163200 86186 164400
rect 86958 163200 87014 164400
rect 87786 163200 87842 164400
rect 88706 163200 88762 164400
rect 89534 163200 89590 164400
rect 90362 163200 90418 164400
rect 91190 163200 91246 164400
rect 92018 163200 92074 164400
rect 92846 163200 92902 164400
rect 93674 163200 93730 164400
rect 94594 163200 94650 164400
rect 95422 163200 95478 164400
rect 96250 163200 96306 164400
rect 97078 163200 97134 164400
rect 97906 163200 97962 164400
rect 98734 163200 98790 164400
rect 99562 163200 99618 164400
rect 100482 163200 100538 164400
rect 101310 163200 101366 164400
rect 102138 163200 102194 164400
rect 102966 163200 103022 164400
rect 103072 163254 103468 163282
rect 84488 158778 84516 163200
rect 84476 158772 84528 158778
rect 84476 158714 84528 158720
rect 85316 155854 85344 163200
rect 85488 158772 85540 158778
rect 85488 158714 85540 158720
rect 85304 155848 85356 155854
rect 85304 155790 85356 155796
rect 84106 152688 84162 152697
rect 84106 152623 84162 152632
rect 82820 152108 82872 152114
rect 82820 152050 82872 152056
rect 81716 151836 81768 151842
rect 81716 151778 81768 151784
rect 78588 151360 78640 151366
rect 78588 151302 78640 151308
rect 81728 149940 81756 151778
rect 82832 149802 82860 152050
rect 85500 151609 85528 158714
rect 86144 158710 86172 163200
rect 86972 160002 87000 163200
rect 87800 160857 87828 163200
rect 88720 162178 88748 163200
rect 88708 162172 88760 162178
rect 88708 162114 88760 162120
rect 87786 160848 87842 160857
rect 87786 160783 87842 160792
rect 86960 159996 87012 160002
rect 86960 159938 87012 159944
rect 86132 158704 86184 158710
rect 86132 158646 86184 158652
rect 89548 155922 89576 163200
rect 89536 155916 89588 155922
rect 89536 155858 89588 155864
rect 90376 152726 90404 163200
rect 91204 159118 91232 163200
rect 92032 162246 92060 163200
rect 92020 162240 92072 162246
rect 92020 162182 92072 162188
rect 92480 159520 92532 159526
rect 92480 159462 92532 159468
rect 91192 159112 91244 159118
rect 91192 159054 91244 159060
rect 92388 159112 92440 159118
rect 92388 159054 92440 159060
rect 90364 152720 90416 152726
rect 90364 152662 90416 152668
rect 89168 152244 89220 152250
rect 89168 152186 89220 152192
rect 88616 152040 88668 152046
rect 88616 151982 88668 151988
rect 85486 151600 85542 151609
rect 85486 151535 85542 151544
rect 85212 150476 85264 150482
rect 85212 150418 85264 150424
rect 85224 149940 85252 150418
rect 88628 149940 88656 151982
rect 89180 149870 89208 152186
rect 92400 151434 92428 159054
rect 92492 155174 92520 159462
rect 92480 155168 92532 155174
rect 92480 155110 92532 155116
rect 92860 154426 92888 163200
rect 93688 160070 93716 163200
rect 94608 161226 94636 163200
rect 95436 162382 95464 163200
rect 95424 162376 95476 162382
rect 95424 162318 95476 162324
rect 94596 161220 94648 161226
rect 94596 161162 94648 161168
rect 93676 160064 93728 160070
rect 93676 160006 93728 160012
rect 96264 156602 96292 163200
rect 96252 156596 96304 156602
rect 96252 156538 96304 156544
rect 92848 154420 92900 154426
rect 92848 154362 92900 154368
rect 97092 152794 97120 163200
rect 97080 152788 97132 152794
rect 97080 152730 97132 152736
rect 95516 152108 95568 152114
rect 95516 152050 95568 152056
rect 92388 151428 92440 151434
rect 92388 151370 92440 151376
rect 92020 150544 92072 150550
rect 92020 150486 92072 150492
rect 92032 149940 92060 150486
rect 95528 149940 95556 152050
rect 97724 151836 97776 151842
rect 97724 151778 97776 151784
rect 97736 149938 97764 151778
rect 97920 151502 97948 163200
rect 98748 162314 98776 163200
rect 98736 162308 98788 162314
rect 98736 162250 98788 162256
rect 99576 157962 99604 163200
rect 100496 159526 100524 163200
rect 101324 161294 101352 163200
rect 102152 162450 102180 163200
rect 102980 163146 103008 163200
rect 103072 163146 103100 163254
rect 102980 163118 103100 163146
rect 102140 162444 102192 162450
rect 102140 162386 102192 162392
rect 101312 161288 101364 161294
rect 101312 161230 101364 161236
rect 100484 159520 100536 159526
rect 100484 159462 100536 159468
rect 99564 157956 99616 157962
rect 99564 157898 99616 157904
rect 103440 154494 103468 163254
rect 103794 163200 103850 164400
rect 104622 163200 104678 164400
rect 105450 163200 105506 164400
rect 106370 163200 106426 164400
rect 107198 163200 107254 164400
rect 107304 163254 107516 163282
rect 103808 158778 103836 163200
rect 104636 161474 104664 163200
rect 104636 161446 104848 161474
rect 103796 158772 103848 158778
rect 103796 158714 103848 158720
rect 103428 154488 103480 154494
rect 103428 154430 103480 154436
rect 102324 151836 102376 151842
rect 102324 151778 102376 151784
rect 97908 151496 97960 151502
rect 97908 151438 97960 151444
rect 98920 150612 98972 150618
rect 98920 150554 98972 150560
rect 98932 149940 98960 150554
rect 102336 149940 102364 151778
rect 104820 151570 104848 161446
rect 105464 154562 105492 163200
rect 106384 157894 106412 163200
rect 107212 163146 107240 163200
rect 107304 163146 107332 163254
rect 107212 163118 107332 163146
rect 106372 157888 106424 157894
rect 106372 157830 106424 157836
rect 105452 154556 105504 154562
rect 105452 154498 105504 154504
rect 107488 152862 107516 163254
rect 108026 163200 108082 164400
rect 108854 163200 108910 164400
rect 109682 163200 109738 164400
rect 110510 163200 110566 164400
rect 111338 163200 111394 164400
rect 111444 163254 111748 163282
rect 108040 161362 108068 163200
rect 108868 162518 108896 163200
rect 108856 162512 108908 162518
rect 108856 162454 108908 162460
rect 108028 161356 108080 161362
rect 108028 161298 108080 161304
rect 109224 159316 109276 159322
rect 109224 159258 109276 159264
rect 109040 158772 109092 158778
rect 109040 158714 109092 158720
rect 109052 153066 109080 158714
rect 109132 157208 109184 157214
rect 109132 157150 109184 157156
rect 109040 153060 109092 153066
rect 109040 153002 109092 153008
rect 107476 152856 107528 152862
rect 107476 152798 107528 152804
rect 109144 152454 109172 157150
rect 109132 152448 109184 152454
rect 109132 152390 109184 152396
rect 109236 152318 109264 159258
rect 109696 156534 109724 163200
rect 110524 159322 110552 163200
rect 111352 163146 111380 163200
rect 111444 163146 111472 163254
rect 111352 163118 111472 163146
rect 110512 159316 110564 159322
rect 110512 159258 110564 159264
rect 109684 156528 109736 156534
rect 109684 156470 109736 156476
rect 109224 152312 109276 152318
rect 109224 152254 109276 152260
rect 110052 152176 110104 152182
rect 110052 152118 110104 152124
rect 109776 151904 109828 151910
rect 109776 151846 109828 151852
rect 104808 151564 104860 151570
rect 104808 151506 104860 151512
rect 105820 150680 105872 150686
rect 105820 150622 105872 150628
rect 105832 149940 105860 150622
rect 97724 149932 97776 149938
rect 97724 149874 97776 149880
rect 89168 149864 89220 149870
rect 89168 149806 89220 149812
rect 82820 149796 82872 149802
rect 82820 149738 82872 149744
rect 78588 149728 78640 149734
rect 74842 149666 75224 149682
rect 78338 149676 78588 149682
rect 78338 149670 78640 149676
rect 74842 149660 75236 149666
rect 74842 149654 75184 149660
rect 78338 149654 78628 149670
rect 75184 149602 75236 149608
rect 68376 149592 68428 149598
rect 64538 149530 64736 149546
rect 68034 149540 68376 149546
rect 68034 149534 68428 149540
rect 64538 149524 64748 149530
rect 64538 149518 64696 149524
rect 68034 149518 68416 149534
rect 64696 149466 64748 149472
rect 61384 149456 61436 149462
rect 6366 149424 6422 149433
rect 6118 149382 6366 149410
rect 16486 149424 16542 149433
rect 16422 149382 16486 149410
rect 6366 149359 6422 149368
rect 20166 149424 20222 149433
rect 19826 149382 20166 149410
rect 16486 149359 16542 149368
rect 40526 149382 40816 149410
rect 43930 149382 44128 149410
rect 47334 149382 47624 149410
rect 50830 149382 51028 149410
rect 57730 149394 57928 149410
rect 61134 149404 61384 149410
rect 61134 149398 61436 149404
rect 57730 149388 57940 149394
rect 57730 149382 57888 149388
rect 20166 149359 20222 149368
rect 40788 149326 40816 149382
rect 44100 149326 44128 149382
rect 47596 149326 47624 149382
rect 51000 149326 51028 149382
rect 61134 149382 61424 149398
rect 109250 149382 109632 149410
rect 57888 149330 57940 149336
rect 40776 149320 40828 149326
rect 40776 149262 40828 149268
rect 44088 149320 44140 149326
rect 44088 149262 44140 149268
rect 47584 149320 47636 149326
rect 47584 149262 47636 149268
rect 50988 149320 51040 149326
rect 50988 149262 51040 149268
rect 109604 149054 109632 149382
rect 109684 149116 109736 149122
rect 109684 149058 109736 149064
rect 109592 149048 109644 149054
rect 109592 148990 109644 148996
rect 109696 111790 109724 149058
rect 109788 134570 109816 151846
rect 110064 147014 110092 152118
rect 110144 152040 110196 152046
rect 110144 151982 110196 151988
rect 110052 147008 110104 147014
rect 110052 146950 110104 146956
rect 110156 145586 110184 151982
rect 110236 151972 110288 151978
rect 110236 151914 110288 151920
rect 110248 146946 110276 151914
rect 110328 151836 110380 151842
rect 110328 151778 110380 151784
rect 110340 147082 110368 151778
rect 111720 151638 111748 163254
rect 112258 163200 112314 164400
rect 113086 163200 113142 164400
rect 113914 163200 113970 164400
rect 114742 163200 114798 164400
rect 115570 163200 115626 164400
rect 116398 163200 116454 164400
rect 117226 163200 117282 164400
rect 118146 163200 118202 164400
rect 118974 163200 119030 164400
rect 119802 163200 119858 164400
rect 120630 163200 120686 164400
rect 121458 163200 121514 164400
rect 122286 163200 122342 164400
rect 122392 163254 122696 163282
rect 112272 161498 112300 163200
rect 112260 161492 112312 161498
rect 112260 161434 112312 161440
rect 113100 157214 113128 163200
rect 113088 157208 113140 157214
rect 113088 157150 113140 157156
rect 113928 152930 113956 163200
rect 114756 161430 114784 163200
rect 115584 161566 115612 163200
rect 115572 161560 115624 161566
rect 115572 161502 115624 161508
rect 114744 161424 114796 161430
rect 114744 161366 114796 161372
rect 116412 158778 116440 163200
rect 116400 158772 116452 158778
rect 116400 158714 116452 158720
rect 117240 152998 117268 163200
rect 118160 154970 118188 163200
rect 118988 158982 119016 163200
rect 118976 158976 119028 158982
rect 118976 158918 119028 158924
rect 119528 158772 119580 158778
rect 119528 158714 119580 158720
rect 119540 155242 119568 158714
rect 118792 155236 118844 155242
rect 118792 155178 118844 155184
rect 119528 155236 119580 155242
rect 119528 155178 119580 155184
rect 118148 154964 118200 154970
rect 118148 154906 118200 154912
rect 118700 153808 118752 153814
rect 118700 153750 118752 153756
rect 118712 153202 118740 153750
rect 118700 153196 118752 153202
rect 118700 153138 118752 153144
rect 117228 152992 117280 152998
rect 117228 152934 117280 152940
rect 113916 152924 113968 152930
rect 113916 152866 113968 152872
rect 116306 152144 116362 152153
rect 114376 152108 114428 152114
rect 116306 152079 116362 152088
rect 114376 152050 114428 152056
rect 113822 152008 113878 152017
rect 113822 151943 113878 151952
rect 111708 151632 111760 151638
rect 111708 151574 111760 151580
rect 112812 149728 112864 149734
rect 112812 149670 112864 149676
rect 112720 149592 112772 149598
rect 112720 149534 112772 149540
rect 111248 149524 111300 149530
rect 111248 149466 111300 149472
rect 111156 149252 111208 149258
rect 111156 149194 111208 149200
rect 111064 149184 111116 149190
rect 111064 149126 111116 149132
rect 110328 147076 110380 147082
rect 110328 147018 110380 147024
rect 110236 146940 110288 146946
rect 110236 146882 110288 146888
rect 110144 145580 110196 145586
rect 110144 145522 110196 145528
rect 109776 134564 109828 134570
rect 109776 134506 109828 134512
rect 111076 113150 111104 149126
rect 111168 114510 111196 149194
rect 111260 124166 111288 149466
rect 112628 149456 112680 149462
rect 112628 149398 112680 149404
rect 112536 149388 112588 149394
rect 112536 149330 112588 149336
rect 112444 149320 112496 149326
rect 112444 149262 112496 149268
rect 111248 124160 111300 124166
rect 111248 124102 111300 124108
rect 112456 117298 112484 149262
rect 112548 121446 112576 149330
rect 112640 122806 112668 149398
rect 112732 126954 112760 149534
rect 112824 132462 112852 149670
rect 113730 144256 113786 144265
rect 113730 144191 113786 144200
rect 113744 143614 113772 144191
rect 113732 143608 113784 143614
rect 113732 143550 113784 143556
rect 112812 132456 112864 132462
rect 112812 132398 112864 132404
rect 112720 126948 112772 126954
rect 112720 126890 112772 126896
rect 112628 122800 112680 122806
rect 112628 122742 112680 122748
rect 112536 121440 112588 121446
rect 112536 121382 112588 121388
rect 112444 117292 112496 117298
rect 112444 117234 112496 117240
rect 111156 114504 111208 114510
rect 111156 114446 111208 114452
rect 111064 113144 111116 113150
rect 111064 113086 111116 113092
rect 109684 111784 109736 111790
rect 109684 111726 109736 111732
rect 113546 110120 113602 110129
rect 113546 110055 113602 110064
rect 113560 109614 113588 110055
rect 113548 109608 113600 109614
rect 113548 109550 113600 109556
rect 113836 93634 113864 151943
rect 114282 150648 114338 150657
rect 114282 150583 114338 150592
rect 114008 150544 114060 150550
rect 114008 150486 114060 150492
rect 114098 150512 114154 150521
rect 113914 149152 113970 149161
rect 113914 149087 113970 149096
rect 113824 93628 113876 93634
rect 113824 93570 113876 93576
rect 113928 92478 113956 149087
rect 114020 140758 114048 150486
rect 114098 150447 114154 150456
rect 114008 140752 114060 140758
rect 114008 140694 114060 140700
rect 114006 132832 114062 132841
rect 114006 132767 114062 132776
rect 113916 92472 113968 92478
rect 113916 92414 113968 92420
rect 114020 86970 114048 132767
rect 114112 104854 114140 150447
rect 114192 149660 114244 149666
rect 114192 149602 114244 149608
rect 114204 131102 114232 149602
rect 114192 131096 114244 131102
rect 114192 131038 114244 131044
rect 114190 121408 114246 121417
rect 114190 121343 114246 121352
rect 114204 118862 114232 121343
rect 114192 118856 114244 118862
rect 114192 118798 114244 118804
rect 114296 109002 114324 150583
rect 114388 141778 114416 152050
rect 116320 151814 116348 152079
rect 118804 151814 118832 155178
rect 119816 153814 119844 163200
rect 120172 159792 120224 159798
rect 120172 159734 120224 159740
rect 120080 158024 120132 158030
rect 120080 157966 120132 157972
rect 119804 153808 119856 153814
rect 119804 153750 119856 153756
rect 120092 151814 120120 157966
rect 120184 155689 120212 159734
rect 120644 159254 120672 163200
rect 120632 159248 120684 159254
rect 120632 159190 120684 159196
rect 121472 158846 121500 163200
rect 122300 163146 122328 163200
rect 122392 163146 122420 163254
rect 122300 163118 122420 163146
rect 121460 158840 121512 158846
rect 121460 158782 121512 158788
rect 120170 155680 120226 155689
rect 120170 155615 120226 155624
rect 121092 155168 121144 155174
rect 121092 155110 121144 155116
rect 116320 151786 116716 151814
rect 118804 151786 119844 151814
rect 120092 151786 120488 151814
rect 116032 150680 116084 150686
rect 116032 150622 116084 150628
rect 114468 150612 114520 150618
rect 114468 150554 114520 150560
rect 114480 143546 114508 150554
rect 116044 147121 116072 150622
rect 116492 149932 116544 149938
rect 116492 149874 116544 149880
rect 116216 149864 116268 149870
rect 116216 149806 116268 149812
rect 116124 149048 116176 149054
rect 116122 149016 116124 149025
rect 116176 149016 116178 149025
rect 116122 148951 116178 148960
rect 116030 147112 116086 147121
rect 116030 147047 116086 147056
rect 116124 147076 116176 147082
rect 116124 147018 116176 147024
rect 116136 145217 116164 147018
rect 116122 145208 116178 145217
rect 116122 145143 116178 145152
rect 115204 143608 115256 143614
rect 115204 143550 115256 143556
rect 114468 143540 114520 143546
rect 114468 143482 114520 143488
rect 114376 141772 114428 141778
rect 114376 141714 114428 141720
rect 114284 108996 114336 109002
rect 114284 108938 114336 108944
rect 114100 104848 114152 104854
rect 114100 104790 114152 104796
rect 114466 98696 114522 98705
rect 114466 98631 114522 98640
rect 114480 96898 114508 98631
rect 114468 96892 114520 96898
rect 114468 96834 114520 96840
rect 115216 91662 115244 143550
rect 115940 143540 115992 143546
rect 115940 143482 115992 143488
rect 115952 143313 115980 143482
rect 115938 143304 115994 143313
rect 115938 143239 115994 143248
rect 115940 141772 115992 141778
rect 115940 141714 115992 141720
rect 115952 141409 115980 141714
rect 115938 141400 115994 141409
rect 115938 141335 115994 141344
rect 115940 140752 115992 140758
rect 115940 140694 115992 140700
rect 115952 139505 115980 140694
rect 115938 139496 115994 139505
rect 115938 139431 115994 139440
rect 116124 132456 116176 132462
rect 116124 132398 116176 132404
rect 116136 131753 116164 132398
rect 116122 131744 116178 131753
rect 116122 131679 116178 131688
rect 115940 131096 115992 131102
rect 115940 131038 115992 131044
rect 115952 129849 115980 131038
rect 115938 129840 115994 129849
rect 115938 129775 115994 129784
rect 116124 126948 116176 126954
rect 116124 126890 116176 126896
rect 116136 126041 116164 126890
rect 116122 126032 116178 126041
rect 116122 125967 116178 125976
rect 116124 124160 116176 124166
rect 116122 124128 116124 124137
rect 116176 124128 116178 124137
rect 116122 124063 116178 124072
rect 115940 122800 115992 122806
rect 115940 122742 115992 122748
rect 115952 122233 115980 122742
rect 115938 122224 115994 122233
rect 115938 122159 115994 122168
rect 115940 121440 115992 121446
rect 115940 121382 115992 121388
rect 115952 120193 115980 121382
rect 115938 120184 115994 120193
rect 115938 120119 115994 120128
rect 115296 118856 115348 118862
rect 115296 118798 115348 118804
rect 115204 91656 115256 91662
rect 115204 91598 115256 91604
rect 114466 87272 114522 87281
rect 114466 87207 114468 87216
rect 114520 87207 114522 87216
rect 114468 87178 114520 87184
rect 114008 86964 114060 86970
rect 114008 86906 114060 86912
rect 115308 83745 115336 118798
rect 116228 118289 116256 149806
rect 116400 145580 116452 145586
rect 116400 145522 116452 145528
rect 116412 137601 116440 145522
rect 116398 137592 116454 137601
rect 116398 137527 116454 137536
rect 116504 133657 116532 149874
rect 116582 149288 116638 149297
rect 116582 149223 116638 149232
rect 116490 133648 116546 133657
rect 116490 133583 116546 133592
rect 116214 118280 116270 118289
rect 116214 118215 116270 118224
rect 116032 117292 116084 117298
rect 116032 117234 116084 117240
rect 116044 116385 116072 117234
rect 116030 116376 116086 116385
rect 116030 116311 116086 116320
rect 116124 114504 116176 114510
rect 116122 114472 116124 114481
rect 116176 114472 116178 114481
rect 116122 114407 116178 114416
rect 116124 113144 116176 113150
rect 116124 113086 116176 113092
rect 116136 112577 116164 113086
rect 116122 112568 116178 112577
rect 116122 112503 116178 112512
rect 116124 111784 116176 111790
rect 116124 111726 116176 111732
rect 116136 110673 116164 111726
rect 116122 110664 116178 110673
rect 116122 110599 116178 110608
rect 115388 109608 115440 109614
rect 115388 109550 115440 109556
rect 115294 83736 115350 83745
rect 115294 83671 115350 83680
rect 115400 81841 115428 109550
rect 116400 108996 116452 109002
rect 116400 108938 116452 108944
rect 116412 108769 116440 108938
rect 116398 108760 116454 108769
rect 116398 108695 116454 108704
rect 115940 104848 115992 104854
rect 115938 104816 115940 104825
rect 115992 104816 115994 104825
rect 115938 104751 115994 104760
rect 116596 97209 116624 149223
rect 116582 97200 116638 97209
rect 116582 97135 116638 97144
rect 116688 95305 116716 151786
rect 118974 151056 119030 151065
rect 118974 150991 119030 151000
rect 117044 150476 117096 150482
rect 117044 150418 117096 150424
rect 116766 149424 116822 149433
rect 116766 149359 116822 149368
rect 116780 99113 116808 149359
rect 116860 147008 116912 147014
rect 116860 146950 116912 146956
rect 116872 101017 116900 146950
rect 116952 146940 117004 146946
rect 116952 146882 117004 146888
rect 116964 106865 116992 146882
rect 117056 135561 117084 150418
rect 118988 149954 119016 150991
rect 119816 150226 119844 151786
rect 120460 150226 120488 151786
rect 121104 150226 121132 155110
rect 122668 153746 122696 163254
rect 123114 163200 123170 164400
rect 124034 163200 124090 164400
rect 124862 163200 124918 164400
rect 125690 163200 125746 164400
rect 126518 163200 126574 164400
rect 127346 163200 127402 164400
rect 128174 163200 128230 164400
rect 129002 163200 129058 164400
rect 129922 163200 129978 164400
rect 130750 163200 130806 164400
rect 131578 163200 131634 164400
rect 132406 163200 132462 164400
rect 133234 163200 133290 164400
rect 134062 163200 134118 164400
rect 134890 163200 134946 164400
rect 135810 163200 135866 164400
rect 136638 163200 136694 164400
rect 137466 163200 137522 164400
rect 138294 163200 138350 164400
rect 139122 163200 139178 164400
rect 139950 163200 140006 164400
rect 140778 163200 140834 164400
rect 141698 163200 141754 164400
rect 142526 163200 142582 164400
rect 143354 163200 143410 164400
rect 144182 163200 144238 164400
rect 145010 163200 145066 164400
rect 145838 163200 145894 164400
rect 146666 163200 146722 164400
rect 147586 163200 147642 164400
rect 148414 163200 148470 164400
rect 149242 163200 149298 164400
rect 150070 163200 150126 164400
rect 150898 163200 150954 164400
rect 151726 163200 151782 164400
rect 152554 163200 152610 164400
rect 153474 163200 153530 164400
rect 154302 163200 154358 164400
rect 155130 163200 155186 164400
rect 155958 163200 156014 164400
rect 156786 163200 156842 164400
rect 157614 163200 157670 164400
rect 158442 163200 158498 164400
rect 159362 163200 159418 164400
rect 160190 163200 160246 164400
rect 161018 163200 161074 164400
rect 161124 163254 161428 163282
rect 122748 158840 122800 158846
rect 122748 158782 122800 158788
rect 121736 153740 121788 153746
rect 121736 153682 121788 153688
rect 122656 153740 122708 153746
rect 122656 153682 122708 153688
rect 121748 150226 121776 153682
rect 122380 152448 122432 152454
rect 122380 152390 122432 152396
rect 122392 150226 122420 152390
rect 122760 151706 122788 158782
rect 123128 157826 123156 163200
rect 124048 159798 124076 163200
rect 124876 160682 124904 163200
rect 125704 161474 125732 163200
rect 125704 161446 125824 161474
rect 124864 160676 124916 160682
rect 124864 160618 124916 160624
rect 124036 159792 124088 159798
rect 124036 159734 124088 159740
rect 124128 159384 124180 159390
rect 124128 159326 124180 159332
rect 123116 157820 123168 157826
rect 123116 157762 123168 157768
rect 123022 155272 123078 155281
rect 123022 155207 123078 155216
rect 122748 151700 122800 151706
rect 122748 151642 122800 151648
rect 119816 150198 119890 150226
rect 120460 150198 120534 150226
rect 121104 150198 121178 150226
rect 121748 150198 121822 150226
rect 122392 150198 122466 150226
rect 118988 149926 119324 149954
rect 119862 149940 119890 150198
rect 120506 149940 120534 150198
rect 121150 149940 121178 150198
rect 121794 149940 121822 150198
rect 122438 149940 122466 150198
rect 123036 150192 123064 155207
rect 123668 152516 123720 152522
rect 123668 152458 123720 152464
rect 123680 150192 123708 152458
rect 124140 152454 124168 159326
rect 125508 158976 125560 158982
rect 125508 158918 125560 158924
rect 124770 156632 124826 156641
rect 124770 156567 124826 156576
rect 124310 153776 124366 153785
rect 124310 153711 124366 153720
rect 124128 152448 124180 152454
rect 124128 152390 124180 152396
rect 124324 150192 124352 153711
rect 124784 151814 124812 156567
rect 125520 153785 125548 158918
rect 125692 156732 125744 156738
rect 125692 156674 125744 156680
rect 125600 155304 125652 155310
rect 125600 155246 125652 155252
rect 125506 153776 125562 153785
rect 125506 153711 125562 153720
rect 124784 151786 124996 151814
rect 124968 150226 124996 151786
rect 124968 150198 125042 150226
rect 123036 150164 123110 150192
rect 123680 150164 123754 150192
rect 124324 150164 124398 150192
rect 123082 149940 123110 150164
rect 123726 149940 123754 150164
rect 124370 149940 124398 150164
rect 125014 149940 125042 150198
rect 125612 150192 125640 155246
rect 125704 152522 125732 156674
rect 125796 155310 125824 161446
rect 126532 156738 126560 163200
rect 127360 159186 127388 163200
rect 127622 159352 127678 159361
rect 127622 159287 127678 159296
rect 127348 159180 127400 159186
rect 127348 159122 127400 159128
rect 127070 157992 127126 158001
rect 127070 157927 127126 157936
rect 126520 156732 126572 156738
rect 126520 156674 126572 156680
rect 125784 155304 125836 155310
rect 125784 155246 125836 155252
rect 126886 153912 126942 153921
rect 126886 153847 126942 153856
rect 125692 152516 125744 152522
rect 125692 152458 125744 152464
rect 126334 152416 126390 152425
rect 126334 152351 126390 152360
rect 126348 150226 126376 152351
rect 126302 150198 126376 150226
rect 125612 150164 125686 150192
rect 125658 149940 125686 150164
rect 126302 149940 126330 150198
rect 126900 150192 126928 153847
rect 127084 150210 127112 157927
rect 127532 152516 127584 152522
rect 127532 152458 127584 152464
rect 127072 150204 127124 150210
rect 126900 150164 126974 150192
rect 126946 149940 126974 150164
rect 127544 150192 127572 152458
rect 127636 151910 127664 159287
rect 128188 155106 128216 163200
rect 128360 159724 128412 159730
rect 128360 159666 128412 159672
rect 128176 155100 128228 155106
rect 128176 155042 128228 155048
rect 128372 153678 128400 159666
rect 129016 158846 129044 163200
rect 129832 159452 129884 159458
rect 129832 159394 129884 159400
rect 129004 158840 129056 158846
rect 129004 158782 129056 158788
rect 129740 156664 129792 156670
rect 129740 156606 129792 156612
rect 129464 153876 129516 153882
rect 129464 153818 129516 153824
rect 128360 153672 128412 153678
rect 128360 153614 128412 153620
rect 128820 152448 128872 152454
rect 128820 152390 128872 152396
rect 127624 151904 127676 151910
rect 127624 151846 127676 151852
rect 128222 150204 128274 150210
rect 127544 150164 127618 150192
rect 127072 150146 127124 150152
rect 127590 149940 127618 150164
rect 128832 150192 128860 152390
rect 129476 150192 129504 153818
rect 129752 151814 129780 156606
rect 129844 152454 129872 159394
rect 129936 156670 129964 163200
rect 130764 159730 130792 163200
rect 130752 159724 130804 159730
rect 130752 159666 130804 159672
rect 131592 158778 131620 163200
rect 132420 159390 132448 163200
rect 132408 159384 132460 159390
rect 132408 159326 132460 159332
rect 132132 158840 132184 158846
rect 132132 158782 132184 158788
rect 131580 158772 131632 158778
rect 131580 158714 131632 158720
rect 129924 156664 129976 156670
rect 129924 156606 129976 156612
rect 130292 155372 130344 155378
rect 130292 155314 130344 155320
rect 129832 152448 129884 152454
rect 129832 152390 129884 152396
rect 130304 151814 130332 155314
rect 132144 153950 132172 158782
rect 132408 158772 132460 158778
rect 132408 158714 132460 158720
rect 132040 153944 132092 153950
rect 132040 153886 132092 153892
rect 132132 153944 132184 153950
rect 132132 153886 132184 153892
rect 131394 152552 131450 152561
rect 131394 152487 131450 152496
rect 129752 151786 130148 151814
rect 130304 151786 130792 151814
rect 130120 150226 130148 151786
rect 130764 150226 130792 151786
rect 130120 150198 130194 150226
rect 130764 150198 130838 150226
rect 128832 150164 128906 150192
rect 129476 150164 129550 150192
rect 128222 150146 128274 150152
rect 128234 149940 128262 150146
rect 128878 149940 128906 150164
rect 129522 149940 129550 150164
rect 130166 149940 130194 150198
rect 130810 149940 130838 150198
rect 131408 150192 131436 152487
rect 132052 150192 132080 153886
rect 132420 151774 132448 158714
rect 132500 158092 132552 158098
rect 132500 158034 132552 158040
rect 132408 151768 132460 151774
rect 132408 151710 132460 151716
rect 132512 150210 132540 158034
rect 133248 158030 133276 163200
rect 133418 159624 133474 159633
rect 133418 159559 133474 159568
rect 133236 158024 133288 158030
rect 133236 157966 133288 157972
rect 132684 156800 132736 156806
rect 132684 156742 132736 156748
rect 132696 150226 132724 156742
rect 133432 156466 133460 159559
rect 133420 156460 133472 156466
rect 133420 156402 133472 156408
rect 134076 152522 134104 163200
rect 134904 155038 134932 163200
rect 135824 161474 135852 163200
rect 135732 161446 135852 161474
rect 135258 156768 135314 156777
rect 135258 156703 135314 156712
rect 134892 155032 134944 155038
rect 134892 154974 134944 154980
rect 134616 154012 134668 154018
rect 134616 153954 134668 153960
rect 134064 152516 134116 152522
rect 134064 152458 134116 152464
rect 133972 151904 134024 151910
rect 133972 151846 134024 151852
rect 133984 150226 134012 151846
rect 134628 150226 134656 153954
rect 135272 150226 135300 156703
rect 135732 153882 135760 161446
rect 135812 159384 135864 159390
rect 135812 159326 135864 159332
rect 135824 155378 135852 159326
rect 136652 156806 136680 163200
rect 137480 159633 137508 163200
rect 137466 159624 137522 159633
rect 137466 159559 137522 159568
rect 138018 159488 138074 159497
rect 138018 159423 138074 159432
rect 137836 156868 137888 156874
rect 137836 156810 137888 156816
rect 136640 156800 136692 156806
rect 136640 156742 136692 156748
rect 136732 155508 136784 155514
rect 136732 155450 136784 155456
rect 135904 155440 135956 155446
rect 135904 155382 135956 155388
rect 135812 155372 135864 155378
rect 135812 155314 135864 155320
rect 135720 153876 135772 153882
rect 135720 153818 135772 153824
rect 135916 150226 135944 155382
rect 136548 152584 136600 152590
rect 136548 152526 136600 152532
rect 136560 150226 136588 152526
rect 136744 151814 136772 155450
rect 136744 151786 137232 151814
rect 137204 150226 137232 151786
rect 137848 150226 137876 156810
rect 138032 151978 138060 159423
rect 138308 155514 138336 163200
rect 139136 159458 139164 163200
rect 139124 159452 139176 159458
rect 139124 159394 139176 159400
rect 139492 158228 139544 158234
rect 139492 158170 139544 158176
rect 139400 156936 139452 156942
rect 139400 156878 139452 156884
rect 138296 155508 138348 155514
rect 138296 155450 138348 155456
rect 138480 154080 138532 154086
rect 138480 154022 138532 154028
rect 138020 151972 138072 151978
rect 138020 151914 138072 151920
rect 138492 150226 138520 154022
rect 139124 152448 139176 152454
rect 139124 152390 139176 152396
rect 139136 150226 139164 152390
rect 132500 150204 132552 150210
rect 131408 150164 131482 150192
rect 132052 150164 132126 150192
rect 131454 149940 131482 150164
rect 132098 149940 132126 150164
rect 132696 150198 132770 150226
rect 132500 150146 132552 150152
rect 132742 149940 132770 150198
rect 133374 150204 133426 150210
rect 133984 150198 134058 150226
rect 134628 150198 134702 150226
rect 135272 150198 135346 150226
rect 135916 150198 135990 150226
rect 136560 150198 136634 150226
rect 137204 150198 137278 150226
rect 137848 150198 137922 150226
rect 138492 150198 138566 150226
rect 139136 150198 139210 150226
rect 139412 150210 139440 156878
rect 139504 151910 139532 158170
rect 139964 158098 139992 163200
rect 140792 159390 140820 163200
rect 141712 160614 141740 163200
rect 141700 160608 141752 160614
rect 141700 160550 141752 160556
rect 140872 159860 140924 159866
rect 140872 159802 140924 159808
rect 140780 159384 140832 159390
rect 140780 159326 140832 159332
rect 139952 158092 140004 158098
rect 139952 158034 140004 158040
rect 140884 156398 140912 159802
rect 140872 156392 140924 156398
rect 140872 156334 140924 156340
rect 142342 155544 142398 155553
rect 142342 155479 142398 155488
rect 139766 155408 139822 155417
rect 139766 155343 139822 155352
rect 139492 151904 139544 151910
rect 139492 151846 139544 151852
rect 139780 150226 139808 155343
rect 141698 152824 141754 152833
rect 141698 152759 141754 152768
rect 141054 151192 141110 151201
rect 141054 151127 141110 151136
rect 133374 150146 133426 150152
rect 133386 149940 133414 150146
rect 134030 149940 134058 150198
rect 134674 149940 134702 150198
rect 135318 149940 135346 150198
rect 135962 149940 135990 150198
rect 136606 149940 136634 150198
rect 137250 149940 137278 150198
rect 137894 149940 137922 150198
rect 138538 149940 138566 150198
rect 139182 149940 139210 150198
rect 139400 150204 139452 150210
rect 139780 150198 139854 150226
rect 139400 150146 139452 150152
rect 139826 149940 139854 150198
rect 140458 150204 140510 150210
rect 140458 150146 140510 150152
rect 140470 149940 140498 150146
rect 141068 150090 141096 151127
rect 141712 150226 141740 152759
rect 142356 150226 142384 155479
rect 142540 155281 142568 163200
rect 143080 159180 143132 159186
rect 143080 159122 143132 159128
rect 142526 155272 142582 155281
rect 142526 155207 142582 155216
rect 143092 152454 143120 159122
rect 143368 154018 143396 163200
rect 144196 159186 144224 163200
rect 144828 159588 144880 159594
rect 144828 159530 144880 159536
rect 144184 159180 144236 159186
rect 144184 159122 144236 159128
rect 143632 158160 143684 158166
rect 143632 158102 143684 158108
rect 143356 154012 143408 154018
rect 143356 153954 143408 153960
rect 143080 152448 143132 152454
rect 143080 152390 143132 152396
rect 142988 151904 143040 151910
rect 142988 151846 143040 151852
rect 143000 150226 143028 151846
rect 143644 150226 143672 158102
rect 144840 157758 144868 159530
rect 145024 158778 145052 163200
rect 145852 158846 145880 163200
rect 145840 158840 145892 158846
rect 145840 158782 145892 158788
rect 145012 158772 145064 158778
rect 145012 158714 145064 158720
rect 146208 158772 146260 158778
rect 146208 158714 146260 158720
rect 145102 158128 145158 158137
rect 145102 158063 145158 158072
rect 144828 157752 144880 157758
rect 144828 157694 144880 157700
rect 144828 154964 144880 154970
rect 144828 154906 144880 154912
rect 144840 152386 144868 154906
rect 144920 153128 144972 153134
rect 144920 153070 144972 153076
rect 144828 152380 144880 152386
rect 144828 152322 144880 152328
rect 144276 151972 144328 151978
rect 144276 151914 144328 151920
rect 144288 150226 144316 151914
rect 144932 150226 144960 153070
rect 141712 150198 141786 150226
rect 142356 150198 142430 150226
rect 143000 150198 143074 150226
rect 143644 150198 143718 150226
rect 144288 150198 144362 150226
rect 144932 150198 145006 150226
rect 145116 150210 145144 158063
rect 145564 154148 145616 154154
rect 145564 154090 145616 154096
rect 145576 150226 145604 154090
rect 146220 151026 146248 158714
rect 146680 155446 146708 163200
rect 146852 160744 146904 160750
rect 146852 160686 146904 160692
rect 146668 155440 146720 155446
rect 146668 155382 146720 155388
rect 146208 151020 146260 151026
rect 146208 150962 146260 150968
rect 146864 150226 146892 160686
rect 147600 152590 147628 163200
rect 148428 160750 148456 163200
rect 149152 160812 149204 160818
rect 149152 160754 149204 160760
rect 148416 160744 148468 160750
rect 148416 160686 148468 160692
rect 147772 159928 147824 159934
rect 147772 159870 147824 159876
rect 147680 157004 147732 157010
rect 147680 156946 147732 156952
rect 147588 152584 147640 152590
rect 147588 152526 147640 152532
rect 147496 151088 147548 151094
rect 147496 151030 147548 151036
rect 141068 150062 141142 150090
rect 141114 149940 141142 150062
rect 141758 149940 141786 150198
rect 142402 149940 142430 150198
rect 143046 149940 143074 150198
rect 143690 149940 143718 150198
rect 144334 149940 144362 150198
rect 144978 149940 145006 150198
rect 145104 150204 145156 150210
rect 145576 150198 145650 150226
rect 145104 150146 145156 150152
rect 145622 149940 145650 150198
rect 146254 150204 146306 150210
rect 146864 150198 146938 150226
rect 146254 150146 146306 150152
rect 146266 149940 146294 150146
rect 146910 149940 146938 150198
rect 147508 150090 147536 151030
rect 147692 150210 147720 156946
rect 147784 154154 147812 159870
rect 147772 154148 147824 154154
rect 147772 154090 147824 154096
rect 148138 154048 148194 154057
rect 148138 153983 148194 153992
rect 148152 150226 148180 153983
rect 147680 150204 147732 150210
rect 148152 150198 148226 150226
rect 149164 150210 149192 160754
rect 149256 160546 149284 163200
rect 149428 162580 149480 162586
rect 149428 162522 149480 162528
rect 149244 160540 149296 160546
rect 149244 160482 149296 160488
rect 149440 150226 149468 162522
rect 150084 156874 150112 163200
rect 150912 159934 150940 163200
rect 150900 159928 150952 159934
rect 150900 159870 150952 159876
rect 150440 158840 150492 158846
rect 150440 158782 150492 158788
rect 150072 156868 150124 156874
rect 150072 156810 150124 156816
rect 150452 155174 150480 158782
rect 150532 158296 150584 158302
rect 150532 158238 150584 158244
rect 150440 155168 150492 155174
rect 150440 155110 150492 155116
rect 147680 150146 147732 150152
rect 147508 150062 147582 150090
rect 147554 149940 147582 150062
rect 148198 149940 148226 150198
rect 148830 150204 148882 150210
rect 148830 150146 148882 150152
rect 149152 150204 149204 150210
rect 149440 150198 149514 150226
rect 150544 150210 150572 158238
rect 150624 155576 150676 155582
rect 150624 155518 150676 155524
rect 150636 150226 150664 155518
rect 151740 151094 151768 163200
rect 151912 162648 151964 162654
rect 151912 162590 151964 162596
rect 151728 151088 151780 151094
rect 151728 151030 151780 151036
rect 149152 150146 149204 150152
rect 148842 149940 148870 150146
rect 149486 149940 149514 150198
rect 150026 150204 150078 150210
rect 150026 150146 150078 150152
rect 150532 150204 150584 150210
rect 150636 150198 150710 150226
rect 150532 150146 150584 150152
rect 150038 149940 150066 150146
rect 150682 149940 150710 150198
rect 151314 150204 151366 150210
rect 151924 150192 151952 162590
rect 152568 158778 152596 163200
rect 152556 158772 152608 158778
rect 152556 158714 152608 158720
rect 153108 158772 153160 158778
rect 153108 158714 153160 158720
rect 152554 151328 152610 151337
rect 152554 151263 152610 151272
rect 151924 150164 151998 150192
rect 151314 150146 151366 150152
rect 151326 149940 151354 150146
rect 151970 149940 151998 150164
rect 152568 150090 152596 151263
rect 153120 150958 153148 158714
rect 153384 158364 153436 158370
rect 153384 158306 153436 158312
rect 153200 154216 153252 154222
rect 153200 154158 153252 154164
rect 153108 150952 153160 150958
rect 153108 150894 153160 150900
rect 153212 150192 153240 154158
rect 153396 151814 153424 158306
rect 153488 158166 153516 163200
rect 153476 158160 153528 158166
rect 153476 158102 153528 158108
rect 154210 155680 154266 155689
rect 154210 155615 154266 155624
rect 154224 151814 154252 155615
rect 154316 154222 154344 163200
rect 155040 160880 155092 160886
rect 155040 160822 155092 160828
rect 154672 155644 154724 155650
rect 154672 155586 154724 155592
rect 154304 154216 154356 154222
rect 154304 154158 154356 154164
rect 153396 151786 153884 151814
rect 154224 151786 154528 151814
rect 153856 150226 153884 151786
rect 154500 150226 154528 151786
rect 153856 150198 153930 150226
rect 154500 150198 154574 150226
rect 154684 150210 154712 155586
rect 155052 151814 155080 160822
rect 155144 160818 155172 163200
rect 155132 160812 155184 160818
rect 155132 160754 155184 160760
rect 155972 159118 156000 163200
rect 156052 159656 156104 159662
rect 156052 159598 156104 159604
rect 155960 159112 156012 159118
rect 155960 159054 156012 159060
rect 156064 158001 156092 159598
rect 156050 157992 156106 158001
rect 156050 157927 156106 157936
rect 156420 157072 156472 157078
rect 156420 157014 156472 157020
rect 155960 154284 156012 154290
rect 155960 154226 156012 154232
rect 155972 153134 156000 154226
rect 155960 153128 156012 153134
rect 155960 153070 156012 153076
rect 155052 151786 155172 151814
rect 155144 150226 155172 151786
rect 153212 150164 153286 150192
rect 152568 150062 152642 150090
rect 152614 149940 152642 150062
rect 153258 149940 153286 150164
rect 153902 149940 153930 150198
rect 154546 149940 154574 150198
rect 154672 150204 154724 150210
rect 155144 150198 155218 150226
rect 154672 150146 154724 150152
rect 155190 149940 155218 150198
rect 155822 150204 155874 150210
rect 156432 150192 156460 157014
rect 156800 155582 156828 163200
rect 157628 159662 157656 163200
rect 158456 161474 158484 163200
rect 158456 161446 158668 161474
rect 157616 159656 157668 159662
rect 157616 159598 157668 159604
rect 157432 159452 157484 159458
rect 157432 159394 157484 159400
rect 157340 155712 157392 155718
rect 157340 155654 157392 155660
rect 156788 155576 156840 155582
rect 156788 155518 156840 155524
rect 157352 152318 157380 155654
rect 157444 154970 157472 159394
rect 157432 154964 157484 154970
rect 157432 154906 157484 154912
rect 158352 153128 158404 153134
rect 158352 153070 158404 153076
rect 157064 152312 157116 152318
rect 157064 152254 157116 152260
rect 157340 152312 157392 152318
rect 157340 152254 157392 152260
rect 157076 150192 157104 152254
rect 157708 151156 157760 151162
rect 157708 151098 157760 151104
rect 156432 150164 156506 150192
rect 157076 150164 157150 150192
rect 155822 150146 155874 150152
rect 155834 149940 155862 150146
rect 156478 149940 156506 150164
rect 157122 149940 157150 150164
rect 157720 150090 157748 151098
rect 158364 150192 158392 153070
rect 158640 151162 158668 161446
rect 158720 159996 158772 160002
rect 158720 159938 158772 159944
rect 158732 158438 158760 159938
rect 159376 159361 159404 163200
rect 159362 159352 159418 159361
rect 159362 159287 159418 159296
rect 158720 158432 158772 158438
rect 158720 158374 158772 158380
rect 158996 158364 159048 158370
rect 158996 158306 159048 158312
rect 158628 151156 158680 151162
rect 158628 151098 158680 151104
rect 159008 150192 159036 158306
rect 160204 156942 160232 163200
rect 161032 163146 161060 163200
rect 161124 163146 161152 163254
rect 161032 163118 161152 163146
rect 160284 160948 160336 160954
rect 160284 160890 160336 160896
rect 160192 156936 160244 156942
rect 160192 156878 160244 156884
rect 159640 153672 159692 153678
rect 159640 153614 159692 153620
rect 159652 150192 159680 153614
rect 160296 150192 160324 160890
rect 161400 153134 161428 163254
rect 161846 163200 161902 164400
rect 162674 163200 162730 164400
rect 163502 163200 163558 164400
rect 164330 163200 164386 164400
rect 165250 163200 165306 164400
rect 166078 163200 166134 164400
rect 166906 163200 166962 164400
rect 167734 163200 167790 164400
rect 168562 163200 168618 164400
rect 169390 163200 169446 164400
rect 170218 163200 170274 164400
rect 171138 163200 171194 164400
rect 171966 163200 172022 164400
rect 172072 163254 172468 163282
rect 161480 161696 161532 161702
rect 161480 161638 161532 161644
rect 161388 153128 161440 153134
rect 161388 153070 161440 153076
rect 160928 152312 160980 152318
rect 160928 152254 160980 152260
rect 160940 150192 160968 152254
rect 161492 150210 161520 161638
rect 161860 160954 161888 163200
rect 161848 160948 161900 160954
rect 161848 160890 161900 160896
rect 161572 157140 161624 157146
rect 161572 157082 161624 157088
rect 161584 150226 161612 157082
rect 162688 156641 162716 163200
rect 163044 158500 163096 158506
rect 163044 158442 163096 158448
rect 162674 156632 162730 156641
rect 162674 156567 162730 156576
rect 162860 151224 162912 151230
rect 162860 151166 162912 151172
rect 161480 150204 161532 150210
rect 158364 150164 158438 150192
rect 159008 150164 159082 150192
rect 159652 150164 159726 150192
rect 160296 150164 160370 150192
rect 160940 150164 161014 150192
rect 157720 150062 157794 150090
rect 157766 149940 157794 150062
rect 158410 149940 158438 150164
rect 159054 149940 159082 150164
rect 159698 149940 159726 150164
rect 160342 149940 160370 150164
rect 160986 149940 161014 150164
rect 161584 150198 161658 150226
rect 161480 150146 161532 150152
rect 161630 149940 161658 150198
rect 162262 150204 162314 150210
rect 162262 150146 162314 150152
rect 162274 149940 162302 150146
rect 162872 150090 162900 151166
rect 163056 150210 163084 158442
rect 163516 158234 163544 163200
rect 164344 160002 164372 163200
rect 164332 159996 164384 160002
rect 164332 159938 164384 159944
rect 165264 158778 165292 163200
rect 165620 161628 165672 161634
rect 165620 161570 165672 161576
rect 165436 161016 165488 161022
rect 165436 160958 165488 160964
rect 165252 158772 165304 158778
rect 165252 158714 165304 158720
rect 163504 158228 163556 158234
rect 163504 158170 163556 158176
rect 164424 156460 164476 156466
rect 164424 156402 164476 156408
rect 163504 154352 163556 154358
rect 163504 154294 163556 154300
rect 163516 150226 163544 154294
rect 164436 151814 164464 156402
rect 164436 151786 164832 151814
rect 164804 150226 164832 151786
rect 165448 150226 165476 160958
rect 165528 160064 165580 160070
rect 165528 160006 165580 160012
rect 165540 158506 165568 160006
rect 165528 158500 165580 158506
rect 165528 158442 165580 158448
rect 165632 151814 165660 161570
rect 166092 160886 166120 163200
rect 166080 160880 166132 160886
rect 166080 160822 166132 160828
rect 166724 158568 166776 158574
rect 166724 158510 166776 158516
rect 165632 151786 166120 151814
rect 166092 150226 166120 151786
rect 166736 150226 166764 158510
rect 166920 150890 166948 163200
rect 167644 158772 167696 158778
rect 167644 158714 167696 158720
rect 167368 153196 167420 153202
rect 167368 153138 167420 153144
rect 166908 150884 166960 150890
rect 166908 150826 166960 150832
rect 167380 150226 167408 153138
rect 167656 151298 167684 158714
rect 167748 153202 167776 163200
rect 168472 161764 168524 161770
rect 168472 161706 168524 161712
rect 168380 158636 168432 158642
rect 168380 158578 168432 158584
rect 167736 153196 167788 153202
rect 167736 153138 167788 153144
rect 167644 151292 167696 151298
rect 167644 151234 167696 151240
rect 168012 151224 168064 151230
rect 168012 151166 168064 151172
rect 168104 151224 168156 151230
rect 168104 151166 168156 151172
rect 163044 150204 163096 150210
rect 163516 150198 163590 150226
rect 163044 150146 163096 150152
rect 162872 150062 162946 150090
rect 162918 149940 162946 150062
rect 163562 149940 163590 150198
rect 164194 150204 164246 150210
rect 164804 150198 164878 150226
rect 165448 150198 165522 150226
rect 166092 150198 166166 150226
rect 166736 150198 166810 150226
rect 167380 150198 167454 150226
rect 164194 150146 164246 150152
rect 164206 149940 164234 150146
rect 164850 149940 164878 150198
rect 165494 149940 165522 150198
rect 166138 149940 166166 150198
rect 166782 149940 166810 150198
rect 167426 149940 167454 150198
rect 168024 150090 168052 151166
rect 168116 150890 168144 151166
rect 168104 150884 168156 150890
rect 168104 150826 168156 150832
rect 168392 150210 168420 158578
rect 168484 151814 168512 161706
rect 168576 153610 168604 163200
rect 169404 157010 169432 163200
rect 169852 161084 169904 161090
rect 169852 161026 169904 161032
rect 169760 159520 169812 159526
rect 169760 159462 169812 159468
rect 169772 158642 169800 159462
rect 169760 158636 169812 158642
rect 169760 158578 169812 158584
rect 169392 157004 169444 157010
rect 169392 156946 169444 156952
rect 168564 153604 168616 153610
rect 168564 153546 168616 153552
rect 168484 151786 168696 151814
rect 168668 150226 168696 151786
rect 168380 150204 168432 150210
rect 168668 150198 168742 150226
rect 169864 150210 169892 161026
rect 170232 159594 170260 163200
rect 171152 159866 171180 163200
rect 171980 163146 172008 163200
rect 172072 163146 172100 163254
rect 171980 163118 172100 163146
rect 171324 161832 171376 161838
rect 171324 161774 171376 161780
rect 171140 159860 171192 159866
rect 171140 159802 171192 159808
rect 170220 159588 170272 159594
rect 170220 159530 170272 159536
rect 169944 157752 169996 157758
rect 169944 157694 169996 157700
rect 169956 150226 169984 157694
rect 171140 157276 171192 157282
rect 171140 157218 171192 157224
rect 168380 150146 168432 150152
rect 168024 150062 168098 150090
rect 168070 149940 168098 150062
rect 168714 149940 168742 150198
rect 169346 150204 169398 150210
rect 169346 150146 169398 150152
rect 169852 150204 169904 150210
rect 169956 150198 170030 150226
rect 171152 150210 171180 157218
rect 171336 150226 171364 161774
rect 172440 154086 172468 163254
rect 172794 163200 172850 164400
rect 173622 163200 173678 164400
rect 174450 163200 174506 164400
rect 175278 163200 175334 164400
rect 176106 163200 176162 164400
rect 177026 163200 177082 164400
rect 177854 163200 177910 164400
rect 178682 163200 178738 164400
rect 179510 163200 179566 164400
rect 180338 163200 180394 164400
rect 180444 163254 180748 163282
rect 172704 162036 172756 162042
rect 172704 161978 172756 161984
rect 172520 156392 172572 156398
rect 172520 156334 172572 156340
rect 172428 154080 172480 154086
rect 172428 154022 172480 154028
rect 169852 150146 169904 150152
rect 169358 149940 169386 150146
rect 170002 149940 170030 150198
rect 170634 150204 170686 150210
rect 170634 150146 170686 150152
rect 171140 150204 171192 150210
rect 171140 150146 171192 150152
rect 171290 150198 171364 150226
rect 172532 150226 172560 156334
rect 171922 150204 171974 150210
rect 170646 149940 170674 150146
rect 171290 149940 171318 150198
rect 172532 150198 172606 150226
rect 172716 150210 172744 161978
rect 172808 157146 172836 163200
rect 173636 158302 173664 163200
rect 174464 159050 174492 163200
rect 175292 161022 175320 163200
rect 175556 161900 175608 161906
rect 175556 161842 175608 161848
rect 175280 161016 175332 161022
rect 175280 160958 175332 160964
rect 175462 160712 175518 160721
rect 175462 160647 175518 160656
rect 174912 159384 174964 159390
rect 174912 159326 174964 159332
rect 174452 159044 174504 159050
rect 174452 158986 174504 158992
rect 173624 158296 173676 158302
rect 173624 158238 173676 158244
rect 172796 157140 172848 157146
rect 172796 157082 172848 157088
rect 174452 155780 174504 155786
rect 174452 155722 174504 155728
rect 173162 151464 173218 151473
rect 173162 151399 173218 151408
rect 171922 150146 171974 150152
rect 171934 149940 171962 150146
rect 172578 149940 172606 150198
rect 172704 150204 172756 150210
rect 172704 150146 172756 150152
rect 173176 150090 173204 151399
rect 174464 150226 174492 155722
rect 174924 152318 174952 159326
rect 175096 152652 175148 152658
rect 175096 152594 175148 152600
rect 174912 152312 174964 152318
rect 174912 152254 174964 152260
rect 175108 150226 175136 152594
rect 173854 150204 173906 150210
rect 174464 150198 174538 150226
rect 175108 150198 175182 150226
rect 173854 150146 173906 150152
rect 173176 150062 173250 150090
rect 173222 149940 173250 150062
rect 173866 149940 173894 150146
rect 174510 149940 174538 150198
rect 175154 149940 175182 150198
rect 175476 150192 175504 160647
rect 175568 151814 175596 161842
rect 176120 157078 176148 163200
rect 176660 159588 176712 159594
rect 176660 159530 176712 159536
rect 176108 157072 176160 157078
rect 176108 157014 176160 157020
rect 176672 156466 176700 159530
rect 177040 158370 177068 163200
rect 177868 159458 177896 163200
rect 178224 161968 178276 161974
rect 178224 161910 178276 161916
rect 177856 159452 177908 159458
rect 177856 159394 177908 159400
rect 177028 158364 177080 158370
rect 177028 158306 177080 158312
rect 177028 157344 177080 157350
rect 177028 157286 177080 157292
rect 176660 156460 176712 156466
rect 176660 156402 176712 156408
rect 175568 151786 176424 151814
rect 176396 150226 176424 151786
rect 177040 150226 177068 157286
rect 177672 154148 177724 154154
rect 177672 154090 177724 154096
rect 177684 150226 177712 154090
rect 178236 151814 178264 161910
rect 178696 153921 178724 163200
rect 179420 159316 179472 159322
rect 179420 159258 179472 159264
rect 179432 158001 179460 159258
rect 179418 157992 179474 158001
rect 179418 157927 179474 157936
rect 179418 157856 179474 157865
rect 179418 157791 179474 157800
rect 178682 153912 178738 153921
rect 178682 153847 178738 153856
rect 178236 151786 179000 151814
rect 178316 151360 178368 151366
rect 178316 151302 178368 151308
rect 176396 150198 176470 150226
rect 177040 150198 177114 150226
rect 177684 150198 177758 150226
rect 175476 150164 175826 150192
rect 175798 149940 175826 150164
rect 176442 149940 176470 150198
rect 177086 149940 177114 150198
rect 177730 149940 177758 150198
rect 178328 150090 178356 151302
rect 178972 150226 179000 151786
rect 178972 150198 179046 150226
rect 179432 150210 179460 157791
rect 179524 157282 179552 163200
rect 180352 163146 180380 163200
rect 180444 163146 180472 163254
rect 180352 163118 180472 163146
rect 179602 158264 179658 158273
rect 179602 158199 179658 158208
rect 179512 157276 179564 157282
rect 179512 157218 179564 157224
rect 179616 150226 179644 158199
rect 180720 151366 180748 163254
rect 181166 163200 181222 164400
rect 181994 163200 182050 164400
rect 182914 163200 182970 164400
rect 183742 163200 183798 164400
rect 184570 163200 184626 164400
rect 185398 163200 185454 164400
rect 186226 163200 186282 164400
rect 187054 163200 187110 164400
rect 187882 163200 187938 164400
rect 188802 163200 188858 164400
rect 189630 163200 189686 164400
rect 190458 163200 190514 164400
rect 191286 163200 191342 164400
rect 192114 163200 192170 164400
rect 192942 163200 192998 164400
rect 193770 163200 193826 164400
rect 194690 163200 194746 164400
rect 195518 163200 195574 164400
rect 195624 163254 195928 163282
rect 181076 162104 181128 162110
rect 181076 162046 181128 162052
rect 180892 161152 180944 161158
rect 180892 161094 180944 161100
rect 180708 151360 180760 151366
rect 180708 151302 180760 151308
rect 180904 150226 180932 161094
rect 180982 156904 181038 156913
rect 180982 156839 181038 156848
rect 178328 150062 178402 150090
rect 178374 149940 178402 150062
rect 179018 149940 179046 150198
rect 179420 150204 179472 150210
rect 179616 150198 179690 150226
rect 179420 150146 179472 150152
rect 179662 149940 179690 150198
rect 180294 150204 180346 150210
rect 180294 150146 180346 150152
rect 180858 150198 180932 150226
rect 180996 150210 181024 156839
rect 181088 151814 181116 162046
rect 181180 160070 181208 163200
rect 181168 160064 181220 160070
rect 181168 160006 181220 160012
rect 182008 154154 182036 163200
rect 182928 156777 182956 163200
rect 183756 161090 183784 163200
rect 183744 161084 183796 161090
rect 183744 161026 183796 161032
rect 184584 159526 184612 163200
rect 184572 159520 184624 159526
rect 184572 159462 184624 159468
rect 184848 159248 184900 159254
rect 184848 159190 184900 159196
rect 183560 158704 183612 158710
rect 183560 158646 183612 158652
rect 182914 156768 182970 156777
rect 182914 156703 182970 156712
rect 182364 154216 182416 154222
rect 182364 154158 182416 154164
rect 181996 154148 182048 154154
rect 181996 154090 182048 154096
rect 182376 152561 182404 154158
rect 182730 152688 182786 152697
rect 182730 152623 182786 152632
rect 182362 152552 182418 152561
rect 182362 152487 182418 152496
rect 181088 151786 181484 151814
rect 181456 150226 181484 151786
rect 180984 150204 181036 150210
rect 180306 149940 180334 150146
rect 180858 149940 180886 150198
rect 181456 150198 181530 150226
rect 180984 150146 181036 150152
rect 181502 149940 181530 150198
rect 182134 150204 182186 150210
rect 182744 150192 182772 152623
rect 183374 151600 183430 151609
rect 183374 151535 183430 151544
rect 182744 150164 182818 150192
rect 182134 150146 182186 150152
rect 182146 149940 182174 150146
rect 182790 149940 182818 150164
rect 183388 150090 183416 151535
rect 183572 150210 183600 158646
rect 184860 158137 184888 159190
rect 185032 158432 185084 158438
rect 185032 158374 185084 158380
rect 184846 158128 184902 158137
rect 184846 158063 184902 158072
rect 184020 155848 184072 155854
rect 184020 155790 184072 155796
rect 183560 150204 183612 150210
rect 184032 150192 184060 155790
rect 185044 151814 185072 158374
rect 185412 154222 185440 163200
rect 185950 160848 186006 160857
rect 185950 160783 186006 160792
rect 185400 154216 185452 154222
rect 185400 154158 185452 154164
rect 185044 151786 185348 151814
rect 185320 150226 185348 151786
rect 184710 150204 184762 150210
rect 184032 150164 184106 150192
rect 183560 150146 183612 150152
rect 183388 150062 183462 150090
rect 183434 149940 183462 150062
rect 184078 149940 184106 150164
rect 185320 150198 185394 150226
rect 184710 150146 184762 150152
rect 184722 149940 184750 150146
rect 185366 149940 185394 150198
rect 185964 150192 185992 160783
rect 186240 155650 186268 163200
rect 186320 162172 186372 162178
rect 186320 162114 186372 162120
rect 186228 155644 186280 155650
rect 186228 155586 186280 155592
rect 186332 151814 186360 162114
rect 187068 158438 187096 163200
rect 187700 159792 187752 159798
rect 187700 159734 187752 159740
rect 187056 158432 187108 158438
rect 187056 158374 187108 158380
rect 187240 155916 187292 155922
rect 187240 155858 187292 155864
rect 186332 151786 186636 151814
rect 186608 150226 186636 151786
rect 186608 150198 186682 150226
rect 185964 150164 186038 150192
rect 186010 149940 186038 150164
rect 186654 149940 186682 150198
rect 187252 150192 187280 155858
rect 187712 152425 187740 159734
rect 187896 159322 187924 163200
rect 187884 159316 187936 159322
rect 187884 159258 187936 159264
rect 188816 154290 188844 163200
rect 189172 162240 189224 162246
rect 189172 162182 189224 162188
rect 188804 154284 188856 154290
rect 188804 154226 188856 154232
rect 187884 152720 187936 152726
rect 187884 152662 187936 152668
rect 187698 152416 187754 152425
rect 187698 152351 187754 152360
rect 187896 150192 187924 152662
rect 188528 151428 188580 151434
rect 188528 151370 188580 151376
rect 187252 150164 187326 150192
rect 187896 150164 187970 150192
rect 187298 149940 187326 150164
rect 187942 149940 187970 150164
rect 188540 150090 188568 151370
rect 189184 150192 189212 162182
rect 189644 155417 189672 163200
rect 190472 158574 190500 163200
rect 190736 162376 190788 162382
rect 190736 162318 190788 162324
rect 190460 158568 190512 158574
rect 190460 158510 190512 158516
rect 190552 158500 190604 158506
rect 190552 158442 190604 158448
rect 189630 155408 189686 155417
rect 189630 155343 189686 155352
rect 189816 154420 189868 154426
rect 189816 154362 189868 154368
rect 189828 150192 189856 154362
rect 190564 150226 190592 158442
rect 190518 150198 190592 150226
rect 190748 150210 190776 162318
rect 191104 161220 191156 161226
rect 191104 161162 191156 161168
rect 191116 150226 191144 161162
rect 191300 159390 191328 163200
rect 191288 159384 191340 159390
rect 191288 159326 191340 159332
rect 192128 154358 192156 163200
rect 192392 156596 192444 156602
rect 192392 156538 192444 156544
rect 192116 154352 192168 154358
rect 192116 154294 192168 154300
rect 192404 150226 192432 156538
rect 192956 155718 192984 163200
rect 193404 162308 193456 162314
rect 193404 162250 193456 162256
rect 193128 159180 193180 159186
rect 193128 159122 193180 159128
rect 192944 155712 192996 155718
rect 192944 155654 192996 155660
rect 193140 152794 193168 159122
rect 193036 152788 193088 152794
rect 193036 152730 193088 152736
rect 193128 152788 193180 152794
rect 193128 152730 193180 152736
rect 193048 150226 193076 152730
rect 193416 151814 193444 162250
rect 193784 157350 193812 163200
rect 194704 159798 194732 163200
rect 195532 163146 195560 163200
rect 195624 163146 195652 163254
rect 195532 163118 195652 163146
rect 194692 159792 194744 159798
rect 194692 159734 194744 159740
rect 195244 159724 195296 159730
rect 195244 159666 195296 159672
rect 195256 158710 195284 159666
rect 195244 158704 195296 158710
rect 195244 158646 195296 158652
rect 194600 158636 194652 158642
rect 194600 158578 194652 158584
rect 193772 157344 193824 157350
rect 193772 157286 193824 157292
rect 194324 156528 194376 156534
rect 194324 156470 194376 156476
rect 194336 151910 194364 156470
rect 194324 151904 194376 151910
rect 194324 151846 194376 151852
rect 193416 151786 194364 151814
rect 193680 151496 193732 151502
rect 193680 151438 193732 151444
rect 190736 150204 190788 150210
rect 189184 150164 189258 150192
rect 189828 150164 189902 150192
rect 188540 150062 188614 150090
rect 188586 149940 188614 150062
rect 189230 149940 189258 150164
rect 189874 149940 189902 150164
rect 190518 149940 190546 150198
rect 191116 150198 191190 150226
rect 190736 150146 190788 150152
rect 191162 149940 191190 150198
rect 191794 150204 191846 150210
rect 192404 150198 192478 150226
rect 193048 150198 193122 150226
rect 191794 150146 191846 150152
rect 191806 149940 191834 150146
rect 192450 149940 192478 150198
rect 193094 149940 193122 150198
rect 193692 150090 193720 151438
rect 194336 150226 194364 151786
rect 194336 150198 194410 150226
rect 194612 150210 194640 158578
rect 194968 157956 195020 157962
rect 194968 157898 195020 157904
rect 194980 150226 195008 157898
rect 195900 151434 195928 163254
rect 196346 163200 196402 164400
rect 197174 163200 197230 164400
rect 198002 163200 198058 164400
rect 198830 163200 198886 164400
rect 199658 163200 199714 164400
rect 200578 163200 200634 164400
rect 201406 163200 201462 164400
rect 202234 163200 202290 164400
rect 203062 163200 203118 164400
rect 203890 163200 203946 164400
rect 204718 163200 204774 164400
rect 205546 163200 205602 164400
rect 206466 163200 206522 164400
rect 207294 163200 207350 164400
rect 208122 163200 208178 164400
rect 208950 163200 209006 164400
rect 209778 163200 209834 164400
rect 210606 163200 210662 164400
rect 211434 163200 211490 164400
rect 212354 163200 212410 164400
rect 213182 163200 213238 164400
rect 214010 163200 214066 164400
rect 214838 163200 214894 164400
rect 215666 163200 215722 164400
rect 216494 163200 216550 164400
rect 217322 163200 217378 164400
rect 218242 163200 218298 164400
rect 219070 163200 219126 164400
rect 219898 163200 219954 164400
rect 220726 163200 220782 164400
rect 221554 163200 221610 164400
rect 222382 163200 222438 164400
rect 223210 163200 223266 164400
rect 224130 163200 224186 164400
rect 224958 163200 225014 164400
rect 225786 163200 225842 164400
rect 226614 163200 226670 164400
rect 227442 163200 227498 164400
rect 228270 163200 228326 164400
rect 229098 163200 229154 164400
rect 230018 163200 230074 164400
rect 230846 163200 230902 164400
rect 231674 163200 231730 164400
rect 232502 163200 232558 164400
rect 233330 163200 233386 164400
rect 234158 163200 234214 164400
rect 234986 163200 235042 164400
rect 235906 163200 235962 164400
rect 236734 163200 236790 164400
rect 237562 163200 237618 164400
rect 238390 163200 238446 164400
rect 239218 163200 239274 164400
rect 240046 163200 240102 164400
rect 240874 163200 240930 164400
rect 241794 163200 241850 164400
rect 242622 163200 242678 164400
rect 243450 163200 243506 164400
rect 244278 163200 244334 164400
rect 245106 163200 245162 164400
rect 245934 163200 245990 164400
rect 246762 163200 246818 164400
rect 247682 163200 247738 164400
rect 248510 163200 248566 164400
rect 249338 163200 249394 164400
rect 250166 163200 250222 164400
rect 250994 163200 251050 164400
rect 251822 163200 251878 164400
rect 252650 163200 252706 164400
rect 253570 163200 253626 164400
rect 254398 163200 254454 164400
rect 255226 163200 255282 164400
rect 256054 163200 256110 164400
rect 256882 163200 256938 164400
rect 257710 163200 257766 164400
rect 258538 163200 258594 164400
rect 259458 163200 259514 164400
rect 260286 163200 260342 164400
rect 261114 163200 261170 164400
rect 261942 163200 261998 164400
rect 262770 163200 262826 164400
rect 263598 163200 263654 164400
rect 264426 163200 264482 164400
rect 265346 163200 265402 164400
rect 266174 163200 266230 164400
rect 267002 163200 267058 164400
rect 267830 163200 267886 164400
rect 268658 163200 268714 164400
rect 269486 163200 269542 164400
rect 270314 163200 270370 164400
rect 271234 163200 271290 164400
rect 272062 163200 272118 164400
rect 272890 163200 272946 164400
rect 273718 163200 273774 164400
rect 274546 163200 274602 164400
rect 275374 163200 275430 164400
rect 276202 163200 276258 164400
rect 277122 163200 277178 164400
rect 277950 163200 278006 164400
rect 278778 163200 278834 164400
rect 279606 163200 279662 164400
rect 280434 163200 280490 164400
rect 281262 163200 281318 164400
rect 282090 163200 282146 164400
rect 283010 163200 283066 164400
rect 283838 163200 283894 164400
rect 284666 163200 284722 164400
rect 285494 163200 285550 164400
rect 286322 163200 286378 164400
rect 287150 163200 287206 164400
rect 287978 163200 288034 164400
rect 288898 163200 288954 164400
rect 289726 163200 289782 164400
rect 290554 163200 290610 164400
rect 291382 163200 291438 164400
rect 292210 163200 292266 164400
rect 293038 163200 293094 164400
rect 293866 163200 293922 164400
rect 294786 163200 294842 164400
rect 295614 163200 295670 164400
rect 295720 163254 295932 163282
rect 196256 161288 196308 161294
rect 196256 161230 196308 161236
rect 195888 151428 195940 151434
rect 195888 151370 195940 151376
rect 196268 150226 196296 161230
rect 196360 158778 196388 163200
rect 196900 162444 196952 162450
rect 196900 162386 196952 162392
rect 196348 158772 196400 158778
rect 196348 158714 196400 158720
rect 196912 150226 196940 162386
rect 197188 158506 197216 163200
rect 198016 159594 198044 163200
rect 198844 161158 198872 163200
rect 198832 161152 198884 161158
rect 198832 161094 198884 161100
rect 198004 159588 198056 159594
rect 198004 159530 198056 159536
rect 197360 159112 197412 159118
rect 197360 159054 197412 159060
rect 197176 158500 197228 158506
rect 197176 158442 197228 158448
rect 197372 153542 197400 159054
rect 198740 158772 198792 158778
rect 198740 158714 198792 158720
rect 198096 155100 198148 155106
rect 198096 155042 198148 155048
rect 197544 154488 197596 154494
rect 197544 154430 197596 154436
rect 197360 153536 197412 153542
rect 197360 153478 197412 153484
rect 197556 150226 197584 154430
rect 198108 153066 198136 155042
rect 198752 154426 198780 158714
rect 199672 155786 199700 163200
rect 200304 161356 200356 161362
rect 200304 161298 200356 161304
rect 200120 157888 200172 157894
rect 200120 157830 200172 157836
rect 199660 155780 199712 155786
rect 199660 155722 199712 155728
rect 199476 154556 199528 154562
rect 199476 154498 199528 154504
rect 198740 154420 198792 154426
rect 198740 154362 198792 154368
rect 198004 153060 198056 153066
rect 198004 153002 198056 153008
rect 198096 153060 198148 153066
rect 198096 153002 198148 153008
rect 198016 151814 198044 153002
rect 198016 151786 198228 151814
rect 198200 150226 198228 151786
rect 198832 151564 198884 151570
rect 198832 151506 198884 151512
rect 193692 150062 193766 150090
rect 193738 149940 193766 150062
rect 194382 149940 194410 150198
rect 194600 150204 194652 150210
rect 194980 150198 195054 150226
rect 194600 150146 194652 150152
rect 195026 149940 195054 150198
rect 195658 150204 195710 150210
rect 196268 150198 196342 150226
rect 196912 150198 196986 150226
rect 197556 150198 197630 150226
rect 198200 150198 198274 150226
rect 195658 150146 195710 150152
rect 195670 149940 195698 150146
rect 196314 149940 196342 150198
rect 196958 149940 196986 150198
rect 197602 149940 197630 150198
rect 198246 149940 198274 150198
rect 198844 150090 198872 151506
rect 199488 150226 199516 154498
rect 200132 150226 200160 157830
rect 199488 150198 199562 150226
rect 200132 150198 200206 150226
rect 200316 150210 200344 161298
rect 200592 158642 200620 163200
rect 201314 159624 201370 159633
rect 201314 159559 201370 159568
rect 200580 158636 200632 158642
rect 200580 158578 200632 158584
rect 201328 157758 201356 159559
rect 201420 159186 201448 163200
rect 202052 162512 202104 162518
rect 202052 162454 202104 162460
rect 201408 159180 201460 159186
rect 201408 159122 201460 159128
rect 201316 157752 201368 157758
rect 201316 157694 201368 157700
rect 201868 155032 201920 155038
rect 201868 154974 201920 154980
rect 200764 152856 200816 152862
rect 200764 152798 200816 152804
rect 200776 150226 200804 152798
rect 201880 152726 201908 154974
rect 201868 152720 201920 152726
rect 201868 152662 201920 152668
rect 202064 150226 202092 162454
rect 202248 158778 202276 163200
rect 203076 158778 203104 163200
rect 202236 158772 202288 158778
rect 202236 158714 202288 158720
rect 202788 158772 202840 158778
rect 202788 158714 202840 158720
rect 203064 158772 203116 158778
rect 203064 158714 203116 158720
rect 202696 151904 202748 151910
rect 202696 151846 202748 151852
rect 202708 150226 202736 151846
rect 202800 151502 202828 158714
rect 203338 157992 203394 158001
rect 203338 157927 203394 157936
rect 202788 151496 202840 151502
rect 202788 151438 202840 151444
rect 203352 150226 203380 157927
rect 203904 155922 203932 163200
rect 204260 161492 204312 161498
rect 204260 161434 204312 161440
rect 204168 159044 204220 159050
rect 204168 158986 204220 158992
rect 203892 155916 203944 155922
rect 203892 155858 203944 155864
rect 204180 152250 204208 158986
rect 204168 152244 204220 152250
rect 204168 152186 204220 152192
rect 204272 151814 204300 161434
rect 204732 159497 204760 163200
rect 205560 161226 205588 163200
rect 205548 161220 205600 161226
rect 205548 161162 205600 161168
rect 204718 159488 204774 159497
rect 204718 159423 204774 159432
rect 205272 157208 205324 157214
rect 205272 157150 205324 157156
rect 204272 151786 204668 151814
rect 203984 151632 204036 151638
rect 203984 151574 204036 151580
rect 198844 150062 198918 150090
rect 198890 149940 198918 150062
rect 199534 149940 199562 150198
rect 200178 149940 200206 150198
rect 200304 150204 200356 150210
rect 200776 150198 200850 150226
rect 200304 150146 200356 150152
rect 200822 149940 200850 150198
rect 201454 150204 201506 150210
rect 202064 150198 202138 150226
rect 202708 150198 202782 150226
rect 203352 150198 203426 150226
rect 201454 150146 201506 150152
rect 201466 149940 201494 150146
rect 202110 149940 202138 150198
rect 202754 149940 202782 150198
rect 203398 149940 203426 150198
rect 203996 150090 204024 151574
rect 204640 150226 204668 151786
rect 205284 150226 205312 157150
rect 206480 155854 206508 163200
rect 207020 161560 207072 161566
rect 207020 161502 207072 161508
rect 206560 161424 206612 161430
rect 206560 161366 206612 161372
rect 206468 155848 206520 155854
rect 206468 155790 206520 155796
rect 205916 152924 205968 152930
rect 205916 152866 205968 152872
rect 205928 150226 205956 152866
rect 206572 150226 206600 161366
rect 207032 151814 207060 161502
rect 207112 159928 207164 159934
rect 207112 159870 207164 159876
rect 207124 157962 207152 159870
rect 207308 158001 207336 163200
rect 208136 159254 208164 163200
rect 208964 159934 208992 163200
rect 208952 159928 209004 159934
rect 208952 159870 209004 159876
rect 208124 159248 208176 159254
rect 208124 159190 208176 159196
rect 208492 158772 208544 158778
rect 208492 158714 208544 158720
rect 207294 157992 207350 158001
rect 207112 157956 207164 157962
rect 207294 157927 207350 157936
rect 207112 157898 207164 157904
rect 207112 157820 207164 157826
rect 207112 157762 207164 157768
rect 207124 152862 207152 157762
rect 207572 155236 207624 155242
rect 207572 155178 207624 155184
rect 207112 152856 207164 152862
rect 207112 152798 207164 152804
rect 207584 151814 207612 155178
rect 208400 153808 208452 153814
rect 208400 153750 208452 153756
rect 208412 151842 208440 153750
rect 208504 153678 208532 158714
rect 209792 157214 209820 163200
rect 210620 159050 210648 163200
rect 211448 159730 211476 163200
rect 212368 161474 212396 163200
rect 212368 161446 212488 161474
rect 211436 159724 211488 159730
rect 211436 159666 211488 159672
rect 210884 159316 210936 159322
rect 210884 159258 210936 159264
rect 210608 159044 210660 159050
rect 210608 158986 210660 158992
rect 209962 158128 210018 158137
rect 209962 158063 210018 158072
rect 209780 157208 209832 157214
rect 209780 157150 209832 157156
rect 209778 153776 209834 153785
rect 209778 153711 209834 153720
rect 208492 153672 208544 153678
rect 208492 153614 208544 153620
rect 208492 152992 208544 152998
rect 208492 152934 208544 152940
rect 208400 151836 208452 151842
rect 207032 151786 207244 151814
rect 207584 151786 207888 151814
rect 207216 150226 207244 151786
rect 207860 150226 207888 151786
rect 208400 151778 208452 151784
rect 208504 150226 208532 152934
rect 209136 152380 209188 152386
rect 209136 152322 209188 152328
rect 209148 150226 209176 152322
rect 209792 150226 209820 153711
rect 204640 150198 204714 150226
rect 205284 150198 205358 150226
rect 205928 150198 206002 150226
rect 206572 150198 206646 150226
rect 207216 150198 207290 150226
rect 207860 150198 207934 150226
rect 208504 150198 208578 150226
rect 209148 150198 209222 150226
rect 209792 150198 209866 150226
rect 209976 150210 210004 158063
rect 210896 152930 210924 159258
rect 212356 159180 212408 159186
rect 212356 159122 212408 159128
rect 212264 153740 212316 153746
rect 212264 153682 212316 153688
rect 210884 152924 210936 152930
rect 210884 152866 210936 152872
rect 210424 151836 210476 151842
rect 210424 151778 210476 151784
rect 210436 150226 210464 151778
rect 211620 151700 211672 151706
rect 211620 151642 211672 151648
rect 203996 150062 204070 150090
rect 204042 149940 204070 150062
rect 204686 149940 204714 150198
rect 205330 149940 205358 150198
rect 205974 149940 206002 150198
rect 206618 149940 206646 150198
rect 207262 149940 207290 150198
rect 207906 149940 207934 150198
rect 208550 149940 208578 150198
rect 209194 149940 209222 150198
rect 209838 149940 209866 150198
rect 209964 150204 210016 150210
rect 210436 150198 210510 150226
rect 209964 150146 210016 150152
rect 210482 149940 210510 150198
rect 211114 150204 211166 150210
rect 211114 150146 211166 150152
rect 211126 149940 211154 150146
rect 211632 150090 211660 151642
rect 212276 150226 212304 153682
rect 212368 152658 212396 159122
rect 212356 152652 212408 152658
rect 212356 152594 212408 152600
rect 212460 151570 212488 161446
rect 212632 159792 212684 159798
rect 212632 159734 212684 159740
rect 212644 152998 212672 159734
rect 213196 154494 213224 163200
rect 213920 160676 213972 160682
rect 213920 160618 213972 160624
rect 213184 154488 213236 154494
rect 213184 154430 213236 154436
rect 212632 152992 212684 152998
rect 212632 152934 212684 152940
rect 212908 152856 212960 152862
rect 212908 152798 212960 152804
rect 212448 151564 212500 151570
rect 212448 151506 212500 151512
rect 212920 150226 212948 152798
rect 213550 152416 213606 152425
rect 213550 152351 213606 152360
rect 213564 150226 213592 152351
rect 213932 151814 213960 160618
rect 214024 159118 214052 163200
rect 214852 159322 214880 163200
rect 214840 159316 214892 159322
rect 214840 159258 214892 159264
rect 214012 159112 214064 159118
rect 214012 159054 214064 159060
rect 215024 159044 215076 159050
rect 215024 158986 215076 158992
rect 215036 156602 215064 158986
rect 215484 156732 215536 156738
rect 215484 156674 215536 156680
rect 215024 156596 215076 156602
rect 215024 156538 215076 156544
rect 214840 155304 214892 155310
rect 214840 155246 214892 155252
rect 213932 151786 214236 151814
rect 214208 150226 214236 151786
rect 214852 150226 214880 155246
rect 215496 150226 215524 156674
rect 215680 154562 215708 163200
rect 216508 155242 216536 163200
rect 216864 159656 216916 159662
rect 216864 159598 216916 159604
rect 216680 159112 216732 159118
rect 216680 159054 216732 159060
rect 216692 156738 216720 159054
rect 216680 156732 216732 156738
rect 216680 156674 216732 156680
rect 216496 155236 216548 155242
rect 216496 155178 216548 155184
rect 215668 154556 215720 154562
rect 215668 154498 215720 154504
rect 216220 153604 216272 153610
rect 216220 153546 216272 153552
rect 216232 152454 216260 153546
rect 216876 153066 216904 159598
rect 217336 159118 217364 163200
rect 218256 159798 218284 163200
rect 218244 159792 218296 159798
rect 218244 159734 218296 159740
rect 217324 159112 217376 159118
rect 217324 159054 217376 159060
rect 218704 158704 218756 158710
rect 218704 158646 218756 158652
rect 218060 156664 218112 156670
rect 218060 156606 218112 156612
rect 217416 153944 217468 153950
rect 217416 153886 217468 153892
rect 216772 153060 216824 153066
rect 216772 153002 216824 153008
rect 216864 153060 216916 153066
rect 216864 153002 216916 153008
rect 216128 152448 216180 152454
rect 216128 152390 216180 152396
rect 216220 152448 216272 152454
rect 216220 152390 216272 152396
rect 216140 150226 216168 152390
rect 216784 150226 216812 153002
rect 217428 150226 217456 153886
rect 218072 150226 218100 156606
rect 218716 150226 218744 158646
rect 219084 155310 219112 163200
rect 219532 155372 219584 155378
rect 219532 155314 219584 155320
rect 219072 155304 219124 155310
rect 219072 155246 219124 155252
rect 219544 151814 219572 155314
rect 219912 153950 219940 163200
rect 220176 159928 220228 159934
rect 220176 159870 220228 159876
rect 220188 158710 220216 159870
rect 220740 158778 220768 163200
rect 220728 158772 220780 158778
rect 220728 158714 220780 158720
rect 220176 158704 220228 158710
rect 220176 158646 220228 158652
rect 220636 158024 220688 158030
rect 220636 157966 220688 157972
rect 219900 153944 219952 153950
rect 219900 153886 219952 153892
rect 219544 151786 220032 151814
rect 219348 151768 219400 151774
rect 219348 151710 219400 151716
rect 212276 150198 212350 150226
rect 212920 150198 212994 150226
rect 213564 150198 213638 150226
rect 214208 150198 214282 150226
rect 214852 150198 214926 150226
rect 215496 150198 215570 150226
rect 216140 150198 216214 150226
rect 216784 150198 216858 150226
rect 217428 150198 217502 150226
rect 218072 150198 218146 150226
rect 218716 150198 218790 150226
rect 211632 150062 211706 150090
rect 211678 149940 211706 150062
rect 212322 149940 212350 150198
rect 212966 149940 212994 150198
rect 213610 149940 213638 150198
rect 214254 149940 214282 150198
rect 214898 149940 214926 150198
rect 215542 149940 215570 150198
rect 216186 149940 216214 150198
rect 216830 149940 216858 150198
rect 217474 149940 217502 150198
rect 218118 149940 218146 150198
rect 218762 149940 218790 150198
rect 219360 150090 219388 151710
rect 220004 150226 220032 151786
rect 220004 150198 220078 150226
rect 219360 150062 219434 150090
rect 219406 149940 219434 150062
rect 220050 149940 220078 150198
rect 220648 150192 220676 157966
rect 221568 157894 221596 163200
rect 222016 159996 222068 160002
rect 222016 159938 222068 159944
rect 221556 157888 221608 157894
rect 221556 157830 221608 157836
rect 221740 155508 221792 155514
rect 221740 155450 221792 155456
rect 221752 152862 221780 155450
rect 221740 152856 221792 152862
rect 221740 152798 221792 152804
rect 221924 152720 221976 152726
rect 221924 152662 221976 152668
rect 221280 152516 221332 152522
rect 221280 152458 221332 152464
rect 221292 150192 221320 152458
rect 221936 150192 221964 152662
rect 222028 152522 222056 159938
rect 222396 159934 222424 163200
rect 222384 159928 222436 159934
rect 222384 159870 222436 159876
rect 222108 159248 222160 159254
rect 222108 159190 222160 159196
rect 222016 152516 222068 152522
rect 222016 152458 222068 152464
rect 222120 152425 222148 159190
rect 222752 156800 222804 156806
rect 222752 156742 222804 156748
rect 222568 153876 222620 153882
rect 222568 153818 222620 153824
rect 222106 152416 222162 152425
rect 222106 152351 222162 152360
rect 222580 150192 222608 153818
rect 222764 151814 222792 156742
rect 223224 155378 223252 163200
rect 223948 159316 224000 159322
rect 223948 159258 224000 159264
rect 223488 159112 223540 159118
rect 223488 159054 223540 159060
rect 223212 155372 223264 155378
rect 223212 155314 223264 155320
rect 223500 153785 223528 159054
rect 223856 157752 223908 157758
rect 223856 157694 223908 157700
rect 223486 153776 223542 153785
rect 223486 153711 223542 153720
rect 222764 151786 223252 151814
rect 223224 150226 223252 151786
rect 223224 150198 223298 150226
rect 220648 150164 220722 150192
rect 221292 150164 221366 150192
rect 221936 150164 222010 150192
rect 222580 150164 222654 150192
rect 220694 149940 220722 150164
rect 221338 149940 221366 150164
rect 221982 149940 222010 150164
rect 222626 149940 222654 150164
rect 223270 149940 223298 150198
rect 223868 150192 223896 157694
rect 223960 152726 223988 159258
rect 224144 158982 224172 163200
rect 224972 159662 225000 163200
rect 225696 159928 225748 159934
rect 225696 159870 225748 159876
rect 224960 159656 225012 159662
rect 224960 159598 225012 159604
rect 224132 158976 224184 158982
rect 224132 158918 224184 158924
rect 224960 158092 225012 158098
rect 224960 158034 225012 158040
rect 224500 152856 224552 152862
rect 224500 152798 224552 152804
rect 224592 152856 224644 152862
rect 224592 152798 224644 152804
rect 223948 152720 224000 152726
rect 223948 152662 224000 152668
rect 224512 150192 224540 152798
rect 224604 152522 224632 152798
rect 224592 152516 224644 152522
rect 224592 152458 224644 152464
rect 224972 150210 225000 158034
rect 225708 158030 225736 159870
rect 225696 158024 225748 158030
rect 225696 157966 225748 157972
rect 225800 155514 225828 163200
rect 225788 155508 225840 155514
rect 225788 155450 225840 155456
rect 226628 155106 226656 163200
rect 227076 160608 227128 160614
rect 227076 160550 227128 160556
rect 226616 155100 226668 155106
rect 226616 155042 226668 155048
rect 225144 154964 225196 154970
rect 225144 154906 225196 154912
rect 224960 150204 225012 150210
rect 223868 150164 223942 150192
rect 224512 150164 224586 150192
rect 223914 149940 223942 150164
rect 224558 149940 224586 150164
rect 225156 150192 225184 154906
rect 226432 152312 226484 152318
rect 226432 152254 226484 152260
rect 225834 150204 225886 150210
rect 225156 150164 225230 150192
rect 224960 150146 225012 150152
rect 225202 149940 225230 150164
rect 226444 150192 226472 152254
rect 227088 150192 227116 160550
rect 227456 159322 227484 163200
rect 227444 159316 227496 159322
rect 227444 159258 227496 159264
rect 228284 159254 228312 163200
rect 228272 159248 228324 159254
rect 228272 159190 228324 159196
rect 227720 158976 227772 158982
rect 227720 158918 227772 158924
rect 227732 156534 227760 158918
rect 227904 158772 227956 158778
rect 227904 158714 227956 158720
rect 227720 156528 227772 156534
rect 227720 156470 227772 156476
rect 227916 155281 227944 158714
rect 229112 158098 229140 163200
rect 229100 158092 229152 158098
rect 229100 158034 229152 158040
rect 227718 155272 227774 155281
rect 227718 155207 227774 155216
rect 227902 155272 227958 155281
rect 227902 155207 227958 155216
rect 227732 150192 227760 155207
rect 230032 155174 230060 163200
rect 230756 160064 230808 160070
rect 230756 160006 230808 160012
rect 230388 159928 230440 159934
rect 230388 159870 230440 159876
rect 229192 155168 229244 155174
rect 229192 155110 229244 155116
rect 230020 155168 230072 155174
rect 230020 155110 230072 155116
rect 228364 154012 228416 154018
rect 228364 153954 228416 153960
rect 228376 150192 228404 153954
rect 229008 152788 229060 152794
rect 229008 152730 229060 152736
rect 229020 150226 229048 152730
rect 229020 150198 229094 150226
rect 229204 150210 229232 155110
rect 230400 152794 230428 159870
rect 230388 152788 230440 152794
rect 230388 152730 230440 152736
rect 230768 152386 230796 160006
rect 230860 158778 230888 163200
rect 231688 159866 231716 163200
rect 231952 160744 232004 160750
rect 231952 160686 232004 160692
rect 231676 159860 231728 159866
rect 231676 159802 231728 159808
rect 230848 158772 230900 158778
rect 230848 158714 230900 158720
rect 230940 155440 230992 155446
rect 230940 155382 230992 155388
rect 230756 152380 230808 152386
rect 230756 152322 230808 152328
rect 229652 151020 229704 151026
rect 229652 150962 229704 150968
rect 226444 150164 226518 150192
rect 227088 150164 227162 150192
rect 227732 150164 227806 150192
rect 228376 150164 228450 150192
rect 225834 150146 225886 150152
rect 225846 149940 225874 150146
rect 226490 149940 226518 150164
rect 227134 149940 227162 150164
rect 227778 149940 227806 150164
rect 228422 149940 228450 150164
rect 229066 149940 229094 150198
rect 229192 150204 229244 150210
rect 229192 150146 229244 150152
rect 229664 150090 229692 150962
rect 230952 150226 230980 155382
rect 231584 152584 231636 152590
rect 231584 152526 231636 152532
rect 231596 150226 231624 152526
rect 231964 151814 231992 160686
rect 232516 155446 232544 163200
rect 232872 160540 232924 160546
rect 232872 160482 232924 160488
rect 232504 155440 232556 155446
rect 232504 155382 232556 155388
rect 231964 151786 232268 151814
rect 232240 150226 232268 151786
rect 232884 150226 232912 160482
rect 233240 157956 233292 157962
rect 233240 157898 233292 157904
rect 230342 150204 230394 150210
rect 230952 150198 231026 150226
rect 231596 150198 231670 150226
rect 232240 150198 232314 150226
rect 232884 150198 232958 150226
rect 233252 150210 233280 157898
rect 233344 153882 233372 163200
rect 234172 160002 234200 163200
rect 234160 159996 234212 160002
rect 234160 159938 234212 159944
rect 233516 156868 233568 156874
rect 233516 156810 233568 156816
rect 233332 153876 233384 153882
rect 233332 153818 233384 153824
rect 233528 150226 233556 156810
rect 235000 152522 235028 163200
rect 235920 158137 235948 163200
rect 236092 158160 236144 158166
rect 235906 158128 235962 158137
rect 236092 158102 236144 158108
rect 235906 158063 235962 158072
rect 234988 152516 235040 152522
rect 234988 152458 235040 152464
rect 234804 151088 234856 151094
rect 234804 151030 234856 151036
rect 230342 150146 230394 150152
rect 229664 150062 229738 150090
rect 229710 149940 229738 150062
rect 230354 149940 230382 150146
rect 230998 149940 231026 150198
rect 231642 149940 231670 150198
rect 232286 149940 232314 150198
rect 232930 149940 232958 150198
rect 233240 150204 233292 150210
rect 233528 150198 233602 150226
rect 233240 150146 233292 150152
rect 233574 149940 233602 150198
rect 234206 150204 234258 150210
rect 234206 150146 234258 150152
rect 234218 149940 234246 150146
rect 234816 150090 234844 151030
rect 235448 150952 235500 150958
rect 235448 150894 235500 150900
rect 235460 150090 235488 150894
rect 236104 150226 236132 158102
rect 236748 156670 236776 163200
rect 237380 160812 237432 160818
rect 237380 160754 237432 160760
rect 236736 156664 236788 156670
rect 236736 156606 236788 156612
rect 236734 152552 236790 152561
rect 236734 152487 236790 152496
rect 236748 150226 236776 152487
rect 237392 150226 237420 160754
rect 237470 159352 237526 159361
rect 237470 159287 237526 159296
rect 237484 153270 237512 159287
rect 237576 159186 237604 163200
rect 238404 159934 238432 163200
rect 238392 159928 238444 159934
rect 238392 159870 238444 159876
rect 237564 159180 237616 159186
rect 237564 159122 237616 159128
rect 238024 158772 238076 158778
rect 238024 158714 238076 158720
rect 238036 155582 238064 158714
rect 239232 157962 239260 163200
rect 239956 159248 240008 159254
rect 239956 159190 240008 159196
rect 239220 157956 239272 157962
rect 239220 157898 239272 157904
rect 237932 155576 237984 155582
rect 237932 155518 237984 155524
rect 238024 155576 238076 155582
rect 238024 155518 238076 155524
rect 237840 153536 237892 153542
rect 237840 153478 237892 153484
rect 237472 153264 237524 153270
rect 237472 153206 237524 153212
rect 237852 150498 237880 153478
rect 237944 151814 237972 155518
rect 239968 153066 239996 159190
rect 240060 156806 240088 163200
rect 240888 160070 240916 163200
rect 240876 160064 240928 160070
rect 240876 160006 240928 160012
rect 241808 158846 241836 163200
rect 242072 160948 242124 160954
rect 242072 160890 242124 160896
rect 241796 158840 241848 158846
rect 241796 158782 241848 158788
rect 240140 156936 240192 156942
rect 240140 156878 240192 156884
rect 240048 156800 240100 156806
rect 240048 156742 240100 156748
rect 239312 153060 239364 153066
rect 239312 153002 239364 153008
rect 239956 153060 240008 153066
rect 239956 153002 240008 153008
rect 237944 151786 238708 151814
rect 237852 150470 238064 150498
rect 238036 150226 238064 150470
rect 238680 150226 238708 151786
rect 239324 150226 239352 153002
rect 239956 151156 240008 151162
rect 239956 151098 240008 151104
rect 236104 150198 236178 150226
rect 236748 150198 236822 150226
rect 237392 150198 237466 150226
rect 238036 150198 238110 150226
rect 238680 150198 238754 150226
rect 239324 150198 239398 150226
rect 234816 150062 234890 150090
rect 235460 150062 235534 150090
rect 234862 149940 234890 150062
rect 235506 149940 235534 150062
rect 236150 149940 236178 150198
rect 236794 149940 236822 150198
rect 237438 149940 237466 150198
rect 238082 149940 238110 150198
rect 238726 149940 238754 150198
rect 239370 149940 239398 150198
rect 239968 150090 239996 151098
rect 240152 150210 240180 156878
rect 240600 153264 240652 153270
rect 240600 153206 240652 153212
rect 240612 150226 240640 153206
rect 241888 153128 241940 153134
rect 241888 153070 241940 153076
rect 241900 150226 241928 153070
rect 242084 151814 242112 160890
rect 242440 159452 242492 159458
rect 242440 159394 242492 159400
rect 242452 152590 242480 159394
rect 242636 158166 242664 163200
rect 242900 158228 242952 158234
rect 242900 158170 242952 158176
rect 242624 158160 242676 158166
rect 242624 158102 242676 158108
rect 242440 152584 242492 152590
rect 242440 152526 242492 152532
rect 242084 151786 242480 151814
rect 242452 150226 242480 151786
rect 240140 150204 240192 150210
rect 240612 150198 240686 150226
rect 240140 150146 240192 150152
rect 239968 150062 240042 150090
rect 240014 149940 240042 150062
rect 240658 149940 240686 150198
rect 241290 150204 241342 150210
rect 241900 150198 241974 150226
rect 242452 150198 242526 150226
rect 242912 150210 242940 158170
rect 243082 156632 243138 156641
rect 243082 156567 243138 156576
rect 243096 150226 243124 156567
rect 243464 154018 243492 163200
rect 243452 154012 243504 154018
rect 243452 153954 243504 153960
rect 244292 153814 244320 163200
rect 245120 159458 245148 163200
rect 245752 160880 245804 160886
rect 245752 160822 245804 160828
rect 245108 159452 245160 159458
rect 245108 159394 245160 159400
rect 244556 158840 244608 158846
rect 244556 158782 244608 158788
rect 244280 153808 244332 153814
rect 244280 153750 244332 153756
rect 244568 152862 244596 158782
rect 245660 157888 245712 157894
rect 245660 157830 245712 157836
rect 245672 153134 245700 157830
rect 245660 153128 245712 153134
rect 245660 153070 245712 153076
rect 244372 152856 244424 152862
rect 244372 152798 244424 152804
rect 244556 152856 244608 152862
rect 244556 152798 244608 152804
rect 244384 150226 244412 152798
rect 245016 151292 245068 151298
rect 245016 151234 245068 151240
rect 241290 150146 241342 150152
rect 241302 149940 241330 150146
rect 241946 149940 241974 150198
rect 242498 149940 242526 150198
rect 242900 150204 242952 150210
rect 243096 150198 243170 150226
rect 242900 150146 242952 150152
rect 243142 149940 243170 150198
rect 243774 150204 243826 150210
rect 244384 150198 244458 150226
rect 243774 150146 243826 150152
rect 243786 149940 243814 150146
rect 244430 149940 244458 150198
rect 245028 150090 245056 151234
rect 245764 150226 245792 160822
rect 245948 158234 245976 163200
rect 245936 158228 245988 158234
rect 245936 158170 245988 158176
rect 246776 156874 246804 163200
rect 247224 159520 247276 159526
rect 247224 159462 247276 159468
rect 247040 159316 247092 159322
rect 247040 159258 247092 159264
rect 246764 156868 246816 156874
rect 246764 156810 246816 156816
rect 247052 156641 247080 159258
rect 247132 157004 247184 157010
rect 247132 156946 247184 156952
rect 247038 156632 247094 156641
rect 247038 156567 247094 156576
rect 246948 153196 247000 153202
rect 246948 153138 247000 153144
rect 246304 151224 246356 151230
rect 246304 151166 246356 151172
rect 245718 150198 245792 150226
rect 245028 150062 245102 150090
rect 245074 149940 245102 150062
rect 245718 149940 245746 150198
rect 246316 150090 246344 151166
rect 246960 150226 246988 153138
rect 246960 150198 247034 150226
rect 247144 150210 247172 156946
rect 247236 153202 247264 159462
rect 247696 159118 247724 163200
rect 247684 159112 247736 159118
rect 247684 159054 247736 159060
rect 248524 158778 248552 163200
rect 248512 158772 248564 158778
rect 248512 158714 248564 158720
rect 249352 156942 249380 163200
rect 250180 161474 250208 163200
rect 250180 161446 250300 161474
rect 249616 158772 249668 158778
rect 249616 158714 249668 158720
rect 249340 156936 249392 156942
rect 249340 156878 249392 156884
rect 248880 156460 248932 156466
rect 248880 156402 248932 156408
rect 247224 153196 247276 153202
rect 247224 153138 247276 153144
rect 247592 152448 247644 152454
rect 247592 152390 247644 152396
rect 247604 150226 247632 152390
rect 248892 150226 248920 156402
rect 249628 152794 249656 158714
rect 250272 154086 250300 161446
rect 251008 159254 251036 163200
rect 251836 159526 251864 163200
rect 251824 159520 251876 159526
rect 251824 159462 251876 159468
rect 250996 159248 251048 159254
rect 250996 159190 251048 159196
rect 251732 159180 251784 159186
rect 251732 159122 251784 159128
rect 251456 158296 251508 158302
rect 251456 158238 251508 158244
rect 250812 157140 250864 157146
rect 250812 157082 250864 157088
rect 250168 154080 250220 154086
rect 250168 154022 250220 154028
rect 250260 154080 250312 154086
rect 250260 154022 250312 154028
rect 249524 152788 249576 152794
rect 249524 152730 249576 152736
rect 249616 152788 249668 152794
rect 249616 152730 249668 152736
rect 249536 150226 249564 152730
rect 250180 150226 250208 154022
rect 250824 150226 250852 157082
rect 251468 150226 251496 158238
rect 251744 156466 251772 159122
rect 252664 158302 252692 163200
rect 252744 161016 252796 161022
rect 252744 160958 252796 160964
rect 252652 158296 252704 158302
rect 252652 158238 252704 158244
rect 252560 157072 252612 157078
rect 252560 157014 252612 157020
rect 251732 156460 251784 156466
rect 251732 156402 251784 156408
rect 252100 152244 252152 152250
rect 252100 152186 252152 152192
rect 252112 150226 252140 152186
rect 246316 150062 246390 150090
rect 246362 149940 246390 150062
rect 247006 149940 247034 150198
rect 247132 150204 247184 150210
rect 247604 150198 247678 150226
rect 247132 150146 247184 150152
rect 247650 149940 247678 150198
rect 248282 150204 248334 150210
rect 248892 150198 248966 150226
rect 249536 150198 249610 150226
rect 250180 150198 250254 150226
rect 250824 150198 250898 150226
rect 251468 150198 251542 150226
rect 252112 150198 252186 150226
rect 252572 150210 252600 157014
rect 252756 150226 252784 160958
rect 253584 157010 253612 163200
rect 254032 158364 254084 158370
rect 254032 158306 254084 158312
rect 253572 157004 253624 157010
rect 253572 156946 253624 156952
rect 254044 150226 254072 158306
rect 254412 157078 254440 163200
rect 254400 157072 254452 157078
rect 254400 157014 254452 157020
rect 255240 152590 255268 163200
rect 255504 159996 255556 160002
rect 255504 159938 255556 159944
rect 255516 153921 255544 159938
rect 256068 158370 256096 163200
rect 256792 159384 256844 159390
rect 256792 159326 256844 159332
rect 256056 158364 256108 158370
rect 256056 158306 256108 158312
rect 256700 157956 256752 157962
rect 256700 157898 256752 157904
rect 255872 157276 255924 157282
rect 255872 157218 255924 157224
rect 255318 153912 255374 153921
rect 255318 153847 255374 153856
rect 255502 153912 255558 153921
rect 255502 153847 255558 153856
rect 254676 152584 254728 152590
rect 254676 152526 254728 152532
rect 255228 152584 255280 152590
rect 255228 152526 255280 152532
rect 254688 150226 254716 152526
rect 255332 150226 255360 153847
rect 255884 151814 255912 157218
rect 256712 152454 256740 157898
rect 256700 152448 256752 152454
rect 256700 152390 256752 152396
rect 256804 152318 256832 159326
rect 256896 158778 256924 163200
rect 257724 159186 257752 163200
rect 258080 161084 258132 161090
rect 258080 161026 258132 161032
rect 257712 159180 257764 159186
rect 257712 159122 257764 159128
rect 256884 158772 256936 158778
rect 256884 158714 256936 158720
rect 257988 158772 258040 158778
rect 257988 158714 258040 158720
rect 258000 154154 258028 158714
rect 257896 154148 257948 154154
rect 257896 154090 257948 154096
rect 257988 154148 258040 154154
rect 257988 154090 258040 154096
rect 257252 152380 257304 152386
rect 257252 152322 257304 152328
rect 256792 152312 256844 152318
rect 256792 152254 256844 152260
rect 255884 151786 256004 151814
rect 255976 150226 256004 151786
rect 256608 151360 256660 151366
rect 256608 151302 256660 151308
rect 248282 150146 248334 150152
rect 248294 149940 248322 150146
rect 248938 149940 248966 150198
rect 249582 149940 249610 150198
rect 250226 149940 250254 150198
rect 250870 149940 250898 150198
rect 251514 149940 251542 150198
rect 252158 149940 252186 150198
rect 252560 150204 252612 150210
rect 252756 150198 252830 150226
rect 252560 150146 252612 150152
rect 252802 149940 252830 150198
rect 253434 150204 253486 150210
rect 254044 150198 254118 150226
rect 254688 150198 254762 150226
rect 255332 150198 255406 150226
rect 255976 150198 256050 150226
rect 253434 150146 253486 150152
rect 253446 149940 253474 150146
rect 254090 149940 254118 150198
rect 254734 149940 254762 150198
rect 255378 149940 255406 150198
rect 256022 149940 256050 150198
rect 256620 150090 256648 151302
rect 257264 150226 257292 152322
rect 257908 150226 257936 154090
rect 257264 150198 257338 150226
rect 257908 150198 257982 150226
rect 258092 150210 258120 161026
rect 258552 160002 258580 163200
rect 258540 159996 258592 160002
rect 258540 159938 258592 159944
rect 259472 157894 259500 163200
rect 259460 157888 259512 157894
rect 259460 157830 259512 157836
rect 260300 157146 260328 163200
rect 260748 159588 260800 159594
rect 260748 159530 260800 159536
rect 260288 157140 260340 157146
rect 260288 157082 260340 157088
rect 258538 156768 258594 156777
rect 258538 156703 258594 156712
rect 258552 150226 258580 156703
rect 260472 154216 260524 154222
rect 260472 154158 260524 154164
rect 259828 153196 259880 153202
rect 259828 153138 259880 153144
rect 259840 150226 259868 153138
rect 260484 150226 260512 154158
rect 260760 152386 260788 159530
rect 261128 159322 261156 163200
rect 261956 159390 261984 163200
rect 261944 159384 261996 159390
rect 261944 159326 261996 159332
rect 261116 159316 261168 159322
rect 261116 159258 261168 159264
rect 262128 159112 262180 159118
rect 262128 159054 262180 159060
rect 260840 158432 260892 158438
rect 260840 158374 260892 158380
rect 260748 152380 260800 152386
rect 260748 152322 260800 152328
rect 256620 150062 256694 150090
rect 256666 149940 256694 150062
rect 257310 149940 257338 150198
rect 257954 149940 257982 150198
rect 258080 150204 258132 150210
rect 258552 150198 258626 150226
rect 258080 150146 258132 150152
rect 258598 149940 258626 150198
rect 259230 150204 259282 150210
rect 259840 150198 259914 150226
rect 260484 150198 260558 150226
rect 260852 150210 260880 158374
rect 261116 155644 261168 155650
rect 261116 155586 261168 155592
rect 261128 150226 261156 155586
rect 262140 154970 262168 159054
rect 262784 157962 262812 163200
rect 263508 159384 263560 159390
rect 263508 159326 263560 159332
rect 262772 157956 262824 157962
rect 262772 157898 262824 157904
rect 262128 154964 262180 154970
rect 262128 154906 262180 154912
rect 263048 154284 263100 154290
rect 263048 154226 263100 154232
rect 262404 152924 262456 152930
rect 262404 152866 262456 152872
rect 262416 150226 262444 152866
rect 263060 150226 263088 154226
rect 263520 152930 263548 159326
rect 263612 154222 263640 163200
rect 263876 160064 263928 160070
rect 263876 160006 263928 160012
rect 263784 158568 263836 158574
rect 263784 158510 263836 158516
rect 263690 155408 263746 155417
rect 263690 155343 263746 155352
rect 263600 154216 263652 154222
rect 263600 154158 263652 154164
rect 263600 153740 263652 153746
rect 263600 153682 263652 153688
rect 263508 152924 263560 152930
rect 263508 152866 263560 152872
rect 259230 150146 259282 150152
rect 259242 149940 259270 150146
rect 259886 149940 259914 150198
rect 260530 149940 260558 150198
rect 260840 150204 260892 150210
rect 261128 150198 261202 150226
rect 260840 150146 260892 150152
rect 261174 149940 261202 150198
rect 261806 150204 261858 150210
rect 262416 150198 262490 150226
rect 263060 150198 263134 150226
rect 263612 150210 263640 153682
rect 263704 150226 263732 155343
rect 263796 153746 263824 158510
rect 263888 155417 263916 160006
rect 264440 159118 264468 163200
rect 265360 160070 265388 163200
rect 265348 160064 265400 160070
rect 265348 160006 265400 160012
rect 265070 159488 265126 159497
rect 265070 159423 265126 159432
rect 264428 159112 264480 159118
rect 264428 159054 264480 159060
rect 263874 155408 263930 155417
rect 263874 155343 263930 155352
rect 263784 153740 263836 153746
rect 263784 153682 263836 153688
rect 265084 152318 265112 159423
rect 266188 158438 266216 163200
rect 266176 158432 266228 158438
rect 266176 158374 266228 158380
rect 266912 157344 266964 157350
rect 266912 157286 266964 157292
rect 265164 155712 265216 155718
rect 265164 155654 265216 155660
rect 264980 152312 265032 152318
rect 264980 152254 265032 152260
rect 265072 152312 265124 152318
rect 265072 152254 265124 152260
rect 264992 150226 265020 152254
rect 261806 150146 261858 150152
rect 261818 149940 261846 150146
rect 262462 149940 262490 150198
rect 263106 149940 263134 150198
rect 263600 150204 263652 150210
rect 263704 150198 263778 150226
rect 263600 150146 263652 150152
rect 263750 149940 263778 150198
rect 264382 150204 264434 150210
rect 264992 150198 265066 150226
rect 265176 150210 265204 155654
rect 265716 154352 265768 154358
rect 265716 154294 265768 154300
rect 265728 150226 265756 154294
rect 264382 150146 264434 150152
rect 264394 149940 264422 150146
rect 265038 149940 265066 150198
rect 265164 150204 265216 150210
rect 265164 150146 265216 150152
rect 265682 150198 265756 150226
rect 266924 150226 266952 157286
rect 267016 154290 267044 163200
rect 267844 159050 267872 163200
rect 267832 159044 267884 159050
rect 267832 158986 267884 158992
rect 268672 158778 268700 163200
rect 268936 159724 268988 159730
rect 268936 159666 268988 159672
rect 268660 158772 268712 158778
rect 268660 158714 268712 158720
rect 268844 154420 268896 154426
rect 268844 154362 268896 154368
rect 267004 154284 267056 154290
rect 267004 154226 267056 154232
rect 267556 152992 267608 152998
rect 267556 152934 267608 152940
rect 267568 150226 267596 152934
rect 268200 151428 268252 151434
rect 268200 151370 268252 151376
rect 266314 150204 266366 150210
rect 265682 149940 265710 150198
rect 266924 150198 266998 150226
rect 267568 150198 267642 150226
rect 266314 150146 266366 150152
rect 266326 149940 266354 150146
rect 266970 149940 266998 150198
rect 267614 149940 267642 150198
rect 268212 150090 268240 151370
rect 268856 150226 268884 154362
rect 268948 153202 268976 159666
rect 269028 159316 269080 159322
rect 269028 159258 269080 159264
rect 269040 155038 269068 159258
rect 269396 158500 269448 158506
rect 269396 158442 269448 158448
rect 269028 155032 269080 155038
rect 269028 154974 269080 154980
rect 268936 153196 268988 153202
rect 268936 153138 268988 153144
rect 269408 151814 269436 158442
rect 269500 157826 269528 163200
rect 269488 157820 269540 157826
rect 269488 157762 269540 157768
rect 270328 154358 270356 163200
rect 270500 161152 270552 161158
rect 270500 161094 270552 161100
rect 270316 154352 270368 154358
rect 270316 154294 270368 154300
rect 270132 152380 270184 152386
rect 270132 152322 270184 152328
rect 269408 151786 269528 151814
rect 269500 150226 269528 151786
rect 270144 150226 270172 152322
rect 270512 151814 270540 161094
rect 271248 159322 271276 163200
rect 272076 159594 272104 163200
rect 272524 159792 272576 159798
rect 272524 159734 272576 159740
rect 272064 159588 272116 159594
rect 272064 159530 272116 159536
rect 271236 159316 271288 159322
rect 271236 159258 271288 159264
rect 271696 158772 271748 158778
rect 271696 158714 271748 158720
rect 271052 155780 271104 155786
rect 271052 155722 271104 155728
rect 271064 151814 271092 155722
rect 271708 152998 271736 158714
rect 272064 158636 272116 158642
rect 272064 158578 272116 158584
rect 271696 152992 271748 152998
rect 271696 152934 271748 152940
rect 270512 151786 270816 151814
rect 271064 151786 271460 151814
rect 270788 150226 270816 151786
rect 271432 150226 271460 151786
rect 272076 150226 272104 158578
rect 272536 152386 272564 159734
rect 272904 158506 272932 163200
rect 272892 158500 272944 158506
rect 272892 158442 272944 158448
rect 273444 155916 273496 155922
rect 273444 155858 273496 155864
rect 272708 152652 272760 152658
rect 272708 152594 272760 152600
rect 272524 152380 272576 152386
rect 272524 152322 272576 152328
rect 272720 150226 272748 152594
rect 273260 151496 273312 151502
rect 273260 151438 273312 151444
rect 268856 150198 268930 150226
rect 269500 150198 269574 150226
rect 270144 150198 270218 150226
rect 270788 150198 270862 150226
rect 271432 150198 271506 150226
rect 272076 150198 272150 150226
rect 272720 150198 272794 150226
rect 268212 150062 268286 150090
rect 268258 149940 268286 150062
rect 268902 149940 268930 150198
rect 269546 149940 269574 150198
rect 270190 149940 270218 150198
rect 270834 149940 270862 150198
rect 271478 149940 271506 150198
rect 272122 149940 272150 150198
rect 272766 149940 272794 150198
rect 273272 150090 273300 151438
rect 273456 150210 273484 155858
rect 273732 155718 273760 163200
rect 274560 158574 274588 163200
rect 274640 159248 274692 159254
rect 274640 159190 274692 159196
rect 274548 158568 274600 158574
rect 274548 158510 274600 158516
rect 273720 155712 273772 155718
rect 273720 155654 273772 155660
rect 274652 153746 274680 159190
rect 275388 158914 275416 163200
rect 275836 161220 275888 161226
rect 275836 161162 275888 161168
rect 275376 158908 275428 158914
rect 275376 158850 275428 158856
rect 274640 153740 274692 153746
rect 274640 153682 274692 153688
rect 273904 153672 273956 153678
rect 273904 153614 273956 153620
rect 273916 150226 273944 153614
rect 275284 152312 275336 152318
rect 275284 152254 275336 152260
rect 275296 150226 275324 152254
rect 273444 150204 273496 150210
rect 273916 150198 273990 150226
rect 273444 150146 273496 150152
rect 273272 150062 273346 150090
rect 273318 149940 273346 150062
rect 273962 149940 273990 150198
rect 274594 150204 274646 150210
rect 274594 150146 274646 150152
rect 275250 150198 275324 150226
rect 275848 150226 275876 161162
rect 276018 157992 276074 158001
rect 276018 157927 276074 157936
rect 275848 150198 275922 150226
rect 276032 150210 276060 157927
rect 276216 157282 276244 163200
rect 276204 157276 276256 157282
rect 276204 157218 276256 157224
rect 276480 155848 276532 155854
rect 276480 155790 276532 155796
rect 276492 150226 276520 155790
rect 277136 155650 277164 163200
rect 277964 159798 277992 163200
rect 277952 159792 278004 159798
rect 277952 159734 278004 159740
rect 278792 158982 278820 163200
rect 279516 159044 279568 159050
rect 279516 158986 279568 158992
rect 278780 158976 278832 158982
rect 278780 158918 278832 158924
rect 278688 158908 278740 158914
rect 278688 158850 278740 158856
rect 277952 158704 278004 158710
rect 277952 158646 278004 158652
rect 277124 155644 277176 155650
rect 277124 155586 277176 155592
rect 277766 152416 277822 152425
rect 277766 152351 277822 152360
rect 277780 150226 277808 152351
rect 277964 151814 277992 158646
rect 278700 152658 278728 158850
rect 278780 157208 278832 157214
rect 278780 157150 278832 157156
rect 278688 152652 278740 152658
rect 278688 152594 278740 152600
rect 278792 151814 278820 157150
rect 279332 156596 279384 156602
rect 279332 156538 279384 156544
rect 279344 151814 279372 156538
rect 279528 156398 279556 158986
rect 279620 158642 279648 163200
rect 279884 159180 279936 159186
rect 279884 159122 279936 159128
rect 279608 158636 279660 158642
rect 279608 158578 279660 158584
rect 279516 156392 279568 156398
rect 279516 156334 279568 156340
rect 279896 153678 279924 159122
rect 280448 155786 280476 163200
rect 281172 159656 281224 159662
rect 281172 159598 281224 159604
rect 280436 155780 280488 155786
rect 280436 155722 280488 155728
rect 279884 153672 279936 153678
rect 279884 153614 279936 153620
rect 281184 153202 281212 159598
rect 281276 158794 281304 163200
rect 282104 159730 282132 163200
rect 282092 159724 282144 159730
rect 282092 159666 282144 159672
rect 281276 158766 281580 158794
rect 281552 154426 281580 158766
rect 283024 156738 283052 163200
rect 282092 156732 282144 156738
rect 282092 156674 282144 156680
rect 283012 156732 283064 156738
rect 283012 156674 283064 156680
rect 281632 154488 281684 154494
rect 281632 154430 281684 154436
rect 281540 154420 281592 154426
rect 281540 154362 281592 154368
rect 280344 153196 280396 153202
rect 280344 153138 280396 153144
rect 281172 153196 281224 153202
rect 281172 153138 281224 153144
rect 277964 151786 278452 151814
rect 278792 151786 279096 151814
rect 279344 151786 279740 151814
rect 278424 150226 278452 151786
rect 279068 150226 279096 151786
rect 279712 150226 279740 151786
rect 280356 150226 280384 153138
rect 280988 151564 281040 151570
rect 280988 151506 281040 151512
rect 274606 149940 274634 150146
rect 275250 149940 275278 150198
rect 275894 149940 275922 150198
rect 276020 150204 276072 150210
rect 276492 150198 276566 150226
rect 276020 150146 276072 150152
rect 276538 149940 276566 150198
rect 277170 150204 277222 150210
rect 277780 150198 277854 150226
rect 278424 150198 278498 150226
rect 279068 150198 279142 150226
rect 279712 150198 279786 150226
rect 280356 150198 280430 150226
rect 277170 150146 277222 150152
rect 277182 149940 277210 150146
rect 277826 149940 277854 150198
rect 278470 149940 278498 150198
rect 279114 149940 279142 150198
rect 279758 149940 279786 150198
rect 280402 149940 280430 150198
rect 281000 150090 281028 151506
rect 281644 150226 281672 154430
rect 282104 151814 282132 156674
rect 283852 155242 283880 163200
rect 284392 159860 284444 159866
rect 284392 159802 284444 159808
rect 284300 159112 284352 159118
rect 284300 159054 284352 159060
rect 283104 155236 283156 155242
rect 283104 155178 283156 155184
rect 283840 155236 283892 155242
rect 283840 155178 283892 155184
rect 282920 152720 282972 152726
rect 282920 152662 282972 152668
rect 282104 151786 282316 151814
rect 282288 150226 282316 151786
rect 282932 150226 282960 152662
rect 281644 150198 281718 150226
rect 282288 150198 282362 150226
rect 282932 150198 283006 150226
rect 283116 150210 283144 155178
rect 284312 154562 284340 159054
rect 283564 154556 283616 154562
rect 283564 154498 283616 154504
rect 284300 154556 284352 154562
rect 284300 154498 284352 154504
rect 283576 150226 283604 154498
rect 284404 152726 284432 159802
rect 284680 159254 284708 163200
rect 285508 159662 285536 163200
rect 285496 159656 285548 159662
rect 285496 159598 285548 159604
rect 284668 159248 284720 159254
rect 284668 159190 284720 159196
rect 286336 158778 286364 163200
rect 287060 159792 287112 159798
rect 287060 159734 287112 159740
rect 287072 159390 287100 159734
rect 287060 159384 287112 159390
rect 287060 159326 287112 159332
rect 286324 158772 286376 158778
rect 286324 158714 286376 158720
rect 286876 158772 286928 158778
rect 286876 158714 286928 158720
rect 286140 155304 286192 155310
rect 286140 155246 286192 155252
rect 284850 153776 284906 153785
rect 284850 153711 284906 153720
rect 284392 152720 284444 152726
rect 284392 152662 284444 152668
rect 284864 150226 284892 153711
rect 285496 152380 285548 152386
rect 285496 152322 285548 152328
rect 285508 150226 285536 152322
rect 286152 150226 286180 155246
rect 286888 153950 286916 158714
rect 287164 155854 287192 163200
rect 287992 159798 288020 163200
rect 288256 159928 288308 159934
rect 288256 159870 288308 159876
rect 287980 159792 288032 159798
rect 287980 159734 288032 159740
rect 287152 155848 287204 155854
rect 287152 155790 287204 155796
rect 287426 155272 287482 155281
rect 287426 155207 287482 155216
rect 286784 153944 286836 153950
rect 286784 153886 286836 153892
rect 286876 153944 286928 153950
rect 286876 153886 286928 153892
rect 286796 150226 286824 153886
rect 287440 150226 287468 155207
rect 288072 153128 288124 153134
rect 288072 153070 288124 153076
rect 288084 150226 288112 153070
rect 288268 152318 288296 159870
rect 288624 159792 288676 159798
rect 288624 159734 288676 159740
rect 288440 158024 288492 158030
rect 288440 157966 288492 157972
rect 288256 152312 288308 152318
rect 288256 152254 288308 152260
rect 288452 151814 288480 157966
rect 288636 157214 288664 159734
rect 288912 158778 288940 163200
rect 288900 158772 288952 158778
rect 288900 158714 288952 158720
rect 289740 158030 289768 163200
rect 289728 158024 289780 158030
rect 289728 157966 289780 157972
rect 288624 157208 288676 157214
rect 288624 157150 288676 157156
rect 290004 156528 290056 156534
rect 290004 156470 290056 156476
rect 289360 155372 289412 155378
rect 289360 155314 289412 155320
rect 288452 151786 288756 151814
rect 288728 150226 288756 151786
rect 289372 150226 289400 155314
rect 290016 150226 290044 156470
rect 290568 155310 290596 163200
rect 291396 159934 291424 163200
rect 291384 159928 291436 159934
rect 291384 159870 291436 159876
rect 292224 159730 292252 163200
rect 291108 159724 291160 159730
rect 291108 159666 291160 159672
rect 292212 159724 292264 159730
rect 292212 159666 292264 159672
rect 290556 155304 290608 155310
rect 290556 155246 290608 155252
rect 291120 153202 291148 159666
rect 291476 159384 291528 159390
rect 291476 159326 291528 159332
rect 291292 155508 291344 155514
rect 291292 155450 291344 155456
rect 291200 155100 291252 155106
rect 291200 155042 291252 155048
rect 290648 153196 290700 153202
rect 290648 153138 290700 153144
rect 291108 153196 291160 153202
rect 291108 153138 291160 153144
rect 290660 150226 290688 153138
rect 281000 150062 281074 150090
rect 281046 149940 281074 150062
rect 281690 149940 281718 150198
rect 282334 149940 282362 150198
rect 282978 149940 283006 150198
rect 283104 150204 283156 150210
rect 283576 150198 283650 150226
rect 283104 150146 283156 150152
rect 283622 149940 283650 150198
rect 284254 150204 284306 150210
rect 284864 150198 284938 150226
rect 285508 150198 285582 150226
rect 286152 150198 286226 150226
rect 286796 150198 286870 150226
rect 287440 150198 287514 150226
rect 288084 150198 288158 150226
rect 288728 150198 288802 150226
rect 289372 150198 289446 150226
rect 290016 150198 290090 150226
rect 290660 150198 290734 150226
rect 291212 150210 291240 155042
rect 291304 150226 291332 155450
rect 291488 155106 291516 159326
rect 292304 158772 292356 158778
rect 292304 158714 292356 158720
rect 291476 155100 291528 155106
rect 291476 155042 291528 155048
rect 292316 153134 292344 158714
rect 293052 158098 293080 163200
rect 292764 158092 292816 158098
rect 292764 158034 292816 158040
rect 293040 158092 293092 158098
rect 293040 158034 293092 158040
rect 292578 156632 292634 156641
rect 292578 156567 292634 156576
rect 292304 153128 292356 153134
rect 292304 153070 292356 153076
rect 292592 150226 292620 156567
rect 284254 150146 284306 150152
rect 284266 149940 284294 150146
rect 284910 149940 284938 150198
rect 285554 149940 285582 150198
rect 286198 149940 286226 150198
rect 286842 149940 286870 150198
rect 287486 149940 287514 150198
rect 288130 149940 288158 150198
rect 288774 149940 288802 150198
rect 289418 149940 289446 150198
rect 290062 149940 290090 150198
rect 290706 149940 290734 150198
rect 291200 150204 291252 150210
rect 291304 150198 291378 150226
rect 291200 150146 291252 150152
rect 291350 149940 291378 150198
rect 291982 150204 292034 150210
rect 292592 150198 292666 150226
rect 292776 150210 292804 158034
rect 293880 155514 293908 163200
rect 294800 155582 294828 163200
rect 295628 163146 295656 163200
rect 295720 163146 295748 163254
rect 295628 163118 295748 163146
rect 294788 155576 294840 155582
rect 294788 155518 294840 155524
rect 293868 155508 293920 155514
rect 293868 155450 293920 155456
rect 295156 155440 295208 155446
rect 295156 155382 295208 155388
rect 294052 155168 294104 155174
rect 294052 155110 294104 155116
rect 293224 153060 293276 153066
rect 293224 153002 293276 153008
rect 293236 150226 293264 153002
rect 294064 151814 294092 155110
rect 294064 151786 294552 151814
rect 294524 150226 294552 151786
rect 295168 150226 295196 155382
rect 295904 152726 295932 163254
rect 296442 163200 296498 164400
rect 297270 163200 297326 164400
rect 298098 163200 298154 164400
rect 298926 163200 298982 164400
rect 299754 163200 299810 164400
rect 300674 163200 300730 164400
rect 301502 163200 301558 164400
rect 302330 163200 302386 164400
rect 303158 163200 303214 164400
rect 303986 163200 304042 164400
rect 304814 163200 304870 164400
rect 305642 163200 305698 164400
rect 306562 163200 306618 164400
rect 307390 163200 307446 164400
rect 308218 163200 308274 164400
rect 309046 163200 309102 164400
rect 309874 163200 309930 164400
rect 310702 163200 310758 164400
rect 311530 163200 311586 164400
rect 312450 163200 312506 164400
rect 313278 163200 313334 164400
rect 314106 163200 314162 164400
rect 314934 163200 314990 164400
rect 315762 163200 315818 164400
rect 316590 163200 316646 164400
rect 317418 163200 317474 164400
rect 318338 163200 318394 164400
rect 319166 163200 319222 164400
rect 319994 163200 320050 164400
rect 320822 163200 320878 164400
rect 321650 163200 321706 164400
rect 322478 163200 322534 164400
rect 322584 163254 322796 163282
rect 296456 157350 296484 163200
rect 296812 159316 296864 159322
rect 296812 159258 296864 159264
rect 296444 157344 296496 157350
rect 296444 157286 296496 157292
rect 296628 155848 296680 155854
rect 296628 155790 296680 155796
rect 296444 155372 296496 155378
rect 296444 155314 296496 155320
rect 295800 152720 295852 152726
rect 295800 152662 295852 152668
rect 295892 152720 295944 152726
rect 295892 152662 295944 152668
rect 295812 150226 295840 152662
rect 296456 150226 296484 155314
rect 296640 155310 296668 155790
rect 296628 155304 296680 155310
rect 296628 155246 296680 155252
rect 296824 153610 296852 159258
rect 297284 155854 297312 163200
rect 298112 159322 298140 163200
rect 298940 159798 298968 163200
rect 298928 159792 298980 159798
rect 298928 159734 298980 159740
rect 299388 159452 299440 159458
rect 299388 159394 299440 159400
rect 298100 159316 298152 159322
rect 298100 159258 298152 159264
rect 298650 158128 298706 158137
rect 298650 158063 298706 158072
rect 297272 155848 297324 155854
rect 297272 155790 297324 155796
rect 297730 153912 297786 153921
rect 297088 153876 297140 153882
rect 297730 153847 297786 153856
rect 297088 153818 297140 153824
rect 296812 153604 296864 153610
rect 296812 153546 296864 153552
rect 297100 150226 297128 153818
rect 297744 150226 297772 153847
rect 298376 152516 298428 152522
rect 298376 152458 298428 152464
rect 298388 150226 298416 152458
rect 298664 151814 298692 158063
rect 299400 153066 299428 159394
rect 299768 156670 299796 163200
rect 299664 156664 299716 156670
rect 299664 156606 299716 156612
rect 299756 156664 299808 156670
rect 299756 156606 299808 156612
rect 299480 156460 299532 156466
rect 299480 156402 299532 156408
rect 299388 153060 299440 153066
rect 299388 153002 299440 153008
rect 298664 151786 299060 151814
rect 299032 150226 299060 151786
rect 291982 150146 292034 150152
rect 291994 149940 292022 150146
rect 292638 149940 292666 150198
rect 292764 150204 292816 150210
rect 293236 150198 293310 150226
rect 292764 150146 292816 150152
rect 293282 149940 293310 150198
rect 293914 150204 293966 150210
rect 294524 150198 294598 150226
rect 295168 150198 295242 150226
rect 295812 150198 295886 150226
rect 296456 150198 296530 150226
rect 297100 150198 297174 150226
rect 297744 150198 297818 150226
rect 298388 150198 298462 150226
rect 299032 150198 299106 150226
rect 299492 150210 299520 156402
rect 299676 150226 299704 156606
rect 300688 155446 300716 163200
rect 301516 158778 301544 163200
rect 301688 159520 301740 159526
rect 301688 159462 301740 159468
rect 301504 158772 301556 158778
rect 301504 158714 301556 158720
rect 300676 155440 300728 155446
rect 300676 155382 300728 155388
rect 301700 152454 301728 159462
rect 302240 156800 302292 156806
rect 302240 156742 302292 156748
rect 301596 152448 301648 152454
rect 301596 152390 301648 152396
rect 301688 152448 301740 152454
rect 301688 152390 301740 152396
rect 300952 152312 301004 152318
rect 300952 152254 301004 152260
rect 300964 150226 300992 152254
rect 301608 150226 301636 152390
rect 293914 150146 293966 150152
rect 293926 149940 293954 150146
rect 294570 149940 294598 150198
rect 295214 149940 295242 150198
rect 295858 149940 295886 150198
rect 296502 149940 296530 150198
rect 297146 149940 297174 150198
rect 297790 149940 297818 150198
rect 298434 149940 298462 150198
rect 299078 149940 299106 150198
rect 299480 150204 299532 150210
rect 299676 150198 299750 150226
rect 299480 150146 299532 150152
rect 299722 149940 299750 150198
rect 300354 150204 300406 150210
rect 300964 150198 301038 150226
rect 301608 150198 301682 150226
rect 300354 150146 300406 150152
rect 300366 149940 300394 150146
rect 301010 149940 301038 150198
rect 301654 149940 301682 150198
rect 302252 150090 302280 156742
rect 302344 152522 302372 163200
rect 303172 156806 303200 163200
rect 303160 156800 303212 156806
rect 303160 156742 303212 156748
rect 304000 156602 304028 163200
rect 304828 159186 304856 163200
rect 305000 159996 305052 160002
rect 305000 159938 305052 159944
rect 304816 159180 304868 159186
rect 304816 159122 304868 159128
rect 304816 158772 304868 158778
rect 304816 158714 304868 158720
rect 304080 158160 304132 158166
rect 304080 158102 304132 158108
rect 303988 156596 304040 156602
rect 303988 156538 304040 156544
rect 302882 155408 302938 155417
rect 302882 155343 302938 155352
rect 302332 152516 302384 152522
rect 302332 152458 302384 152464
rect 302896 150090 302924 155343
rect 303528 152856 303580 152862
rect 303528 152798 303580 152804
rect 303540 150090 303568 152798
rect 304092 150226 304120 158102
rect 304828 154018 304856 158714
rect 304724 154012 304776 154018
rect 304724 153954 304776 153960
rect 304816 154012 304868 154018
rect 304816 153954 304868 153960
rect 304092 150198 304166 150226
rect 302252 150062 302326 150090
rect 302896 150062 302970 150090
rect 303540 150062 303614 150090
rect 302298 149940 302326 150062
rect 302942 149940 302970 150062
rect 303586 149940 303614 150062
rect 304138 149940 304166 150198
rect 304736 150090 304764 153954
rect 305012 152862 305040 159938
rect 305656 159866 305684 163200
rect 306576 161474 306604 163200
rect 306576 161446 306696 161474
rect 305644 159860 305696 159866
rect 305644 159802 305696 159808
rect 305460 159248 305512 159254
rect 305460 159190 305512 159196
rect 305472 153814 305500 159190
rect 306380 158228 306432 158234
rect 306380 158170 306432 158176
rect 306392 157334 306420 158170
rect 306392 157306 306604 157334
rect 306380 156936 306432 156942
rect 306380 156878 306432 156884
rect 306392 156466 306420 156878
rect 306380 156460 306432 156466
rect 306380 156402 306432 156408
rect 305368 153808 305420 153814
rect 305368 153750 305420 153756
rect 305460 153808 305512 153814
rect 305460 153750 305512 153756
rect 305000 152856 305052 152862
rect 305000 152798 305052 152804
rect 305380 150090 305408 153750
rect 306012 153060 306064 153066
rect 306012 153002 306064 153008
rect 306024 150090 306052 153002
rect 306576 150226 306604 157306
rect 306668 156874 306696 161446
rect 307404 158166 307432 163200
rect 308232 159526 308260 163200
rect 308220 159520 308272 159526
rect 308220 159462 308272 159468
rect 307392 158160 307444 158166
rect 307392 158102 307444 158108
rect 307024 157004 307076 157010
rect 307024 156946 307076 156952
rect 306656 156868 306708 156874
rect 306656 156810 306708 156816
rect 307036 156534 307064 156946
rect 307300 156936 307352 156942
rect 307300 156878 307352 156884
rect 307024 156528 307076 156534
rect 307024 156470 307076 156476
rect 306576 150198 306742 150226
rect 304736 150062 304810 150090
rect 305380 150062 305454 150090
rect 306024 150062 306098 150090
rect 304782 149940 304810 150062
rect 305426 149940 305454 150062
rect 306070 149940 306098 150062
rect 306714 149940 306742 150198
rect 307312 150090 307340 156878
rect 307944 154964 307996 154970
rect 307944 154906 307996 154912
rect 307956 150090 307984 154906
rect 309060 152794 309088 163200
rect 309888 161474 309916 163200
rect 309888 161446 310008 161474
rect 309232 156460 309284 156466
rect 309232 156402 309284 156408
rect 308588 152788 308640 152794
rect 308588 152730 308640 152736
rect 309048 152788 309100 152794
rect 309048 152730 309100 152736
rect 308600 150090 308628 152730
rect 309244 150090 309272 156402
rect 309876 154080 309928 154086
rect 309876 154022 309928 154028
rect 309888 150090 309916 154022
rect 309980 153882 310008 161446
rect 310612 158296 310664 158302
rect 310612 158238 310664 158244
rect 309968 153876 310020 153882
rect 309968 153818 310020 153824
rect 310520 153740 310572 153746
rect 310520 153682 310572 153688
rect 310532 150090 310560 153682
rect 310624 150210 310652 158238
rect 310716 156942 310744 163200
rect 311072 160064 311124 160070
rect 311072 160006 311124 160012
rect 310704 156936 310756 156942
rect 310704 156878 310756 156884
rect 311084 152318 311112 160006
rect 311544 160002 311572 163200
rect 311532 159996 311584 160002
rect 311532 159938 311584 159944
rect 311900 159928 311952 159934
rect 311900 159870 311952 159876
rect 311912 157758 311940 159870
rect 312464 159458 312492 163200
rect 312452 159452 312504 159458
rect 312452 159394 312504 159400
rect 311992 159316 312044 159322
rect 311992 159258 312044 159264
rect 311900 157752 311952 157758
rect 311900 157694 311952 157700
rect 311900 157072 311952 157078
rect 311900 157014 311952 157020
rect 311164 152448 311216 152454
rect 311164 152390 311216 152396
rect 311072 152312 311124 152318
rect 311072 152254 311124 152260
rect 310612 150204 310664 150210
rect 310612 150146 310664 150152
rect 311176 150090 311204 152390
rect 311912 151814 311940 157014
rect 312004 156466 312032 159258
rect 312452 156528 312504 156534
rect 312452 156470 312504 156476
rect 311992 156460 312044 156466
rect 311992 156402 312044 156408
rect 311912 151786 312032 151814
rect 312004 150210 312032 151786
rect 312464 150226 312492 156470
rect 313292 154494 313320 163200
rect 314120 158234 314148 163200
rect 314384 158364 314436 158370
rect 314384 158306 314436 158312
rect 314108 158228 314160 158234
rect 314108 158170 314160 158176
rect 313280 154488 313332 154494
rect 313280 154430 313332 154436
rect 313740 152584 313792 152590
rect 313740 152526 313792 152532
rect 313752 150226 313780 152526
rect 314396 150226 314424 158306
rect 314948 152590 314976 163200
rect 315776 158846 315804 163200
rect 315764 158840 315816 158846
rect 315764 158782 315816 158788
rect 315028 154148 315080 154154
rect 315028 154090 315080 154096
rect 314936 152584 314988 152590
rect 314936 152526 314988 152532
rect 315040 150226 315068 154090
rect 316604 154086 316632 163200
rect 317432 158302 317460 163200
rect 318352 160070 318380 163200
rect 318340 160064 318392 160070
rect 318340 160006 318392 160012
rect 319180 159526 319208 163200
rect 317788 159520 317840 159526
rect 317788 159462 317840 159468
rect 319168 159520 319220 159526
rect 319168 159462 319220 159468
rect 317420 158296 317472 158302
rect 317420 158238 317472 158244
rect 316960 157888 317012 157894
rect 316960 157830 317012 157836
rect 316592 154080 316644 154086
rect 316592 154022 316644 154028
rect 315672 153672 315724 153678
rect 315672 153614 315724 153620
rect 315684 150226 315712 153614
rect 316316 152856 316368 152862
rect 316316 152798 316368 152804
rect 316328 150226 316356 152798
rect 316972 150226 317000 157830
rect 317420 157140 317472 157146
rect 317420 157082 317472 157088
rect 317432 151814 317460 157082
rect 317800 156534 317828 159462
rect 318708 158840 318760 158846
rect 318708 158782 318760 158788
rect 317788 156528 317840 156534
rect 317788 156470 317840 156476
rect 317972 155032 318024 155038
rect 317972 154974 318024 154980
rect 317984 151814 318012 154974
rect 318720 153066 318748 158782
rect 319536 157956 319588 157962
rect 319536 157898 319588 157904
rect 318708 153060 318760 153066
rect 318708 153002 318760 153008
rect 318892 152924 318944 152930
rect 318892 152866 318944 152872
rect 317432 151786 317644 151814
rect 317984 151786 318288 151814
rect 317616 150226 317644 151786
rect 318260 150226 318288 151786
rect 318904 150226 318932 152866
rect 319548 150226 319576 157898
rect 320008 154154 320036 163200
rect 320732 159588 320784 159594
rect 320732 159530 320784 159536
rect 320180 154216 320232 154222
rect 320180 154158 320232 154164
rect 319996 154148 320048 154154
rect 319996 154090 320048 154096
rect 320192 150226 320220 154158
rect 320744 151910 320772 159530
rect 320836 158370 320864 163200
rect 321664 158710 321692 163200
rect 322492 163146 322520 163200
rect 322584 163146 322612 163254
rect 322492 163118 322612 163146
rect 321652 158704 321704 158710
rect 321652 158646 321704 158652
rect 322112 158432 322164 158438
rect 322112 158374 322164 158380
rect 320824 158364 320876 158370
rect 320824 158306 320876 158312
rect 320916 154556 320968 154562
rect 320916 154498 320968 154504
rect 320732 151904 320784 151910
rect 320732 151846 320784 151852
rect 320928 150226 320956 154498
rect 321468 152448 321520 152454
rect 321468 152390 321520 152396
rect 311854 150204 311906 150210
rect 311854 150146 311906 150152
rect 311992 150204 312044 150210
rect 312464 150198 312538 150226
rect 311992 150146 312044 150152
rect 307312 150062 307386 150090
rect 307956 150062 308030 150090
rect 308600 150062 308674 150090
rect 309244 150062 309318 150090
rect 309888 150062 309962 150090
rect 310532 150062 310606 150090
rect 311176 150062 311250 150090
rect 307358 149940 307386 150062
rect 308002 149940 308030 150062
rect 308646 149940 308674 150062
rect 309290 149940 309318 150062
rect 309934 149940 309962 150062
rect 310578 149940 310606 150062
rect 311222 149940 311250 150062
rect 311866 149940 311894 150146
rect 312510 149940 312538 150198
rect 313142 150204 313194 150210
rect 313752 150198 313826 150226
rect 314396 150198 314470 150226
rect 315040 150198 315114 150226
rect 315684 150198 315758 150226
rect 316328 150198 316402 150226
rect 316972 150198 317046 150226
rect 317616 150198 317690 150226
rect 318260 150198 318334 150226
rect 318904 150198 318978 150226
rect 319548 150198 319622 150226
rect 320192 150198 320266 150226
rect 313142 150146 313194 150152
rect 313154 149940 313182 150146
rect 313798 149940 313826 150198
rect 314442 149940 314470 150198
rect 315086 149940 315114 150198
rect 315730 149940 315758 150198
rect 316374 149940 316402 150198
rect 317018 149940 317046 150198
rect 317662 149940 317690 150198
rect 318306 149940 318334 150198
rect 318950 149940 318978 150198
rect 319594 149940 319622 150198
rect 320238 149940 320266 150198
rect 320882 150198 320956 150226
rect 321480 150226 321508 152390
rect 322124 150226 322152 158374
rect 322768 152862 322796 163254
rect 323306 163200 323362 164400
rect 324226 163200 324282 164400
rect 325054 163200 325110 164400
rect 325882 163200 325938 164400
rect 326710 163200 326766 164400
rect 326816 163254 327028 163282
rect 322848 154284 322900 154290
rect 322848 154226 322900 154232
rect 322756 152856 322808 152862
rect 322756 152798 322808 152804
rect 322860 150226 322888 154226
rect 323320 154222 323348 163200
rect 323400 156392 323452 156398
rect 323400 156334 323452 156340
rect 323308 154216 323360 154222
rect 323308 154158 323360 154164
rect 321480 150198 321554 150226
rect 322124 150198 322198 150226
rect 320882 149940 320910 150198
rect 321526 149940 321554 150198
rect 322170 149940 322198 150198
rect 322814 150198 322888 150226
rect 323412 150226 323440 156334
rect 324240 155922 324268 163200
rect 325068 159322 325096 163200
rect 325896 159934 325924 163200
rect 326724 163146 326752 163200
rect 326816 163146 326844 163254
rect 326724 163118 326844 163146
rect 325884 159928 325936 159934
rect 325884 159870 325936 159876
rect 325056 159316 325108 159322
rect 325056 159258 325108 159264
rect 324320 159180 324372 159186
rect 324320 159122 324372 159128
rect 324332 157962 324360 159122
rect 324320 157956 324372 157962
rect 324320 157898 324372 157904
rect 324688 157820 324740 157826
rect 324688 157762 324740 157768
rect 324228 155916 324280 155922
rect 324228 155858 324280 155864
rect 324044 152992 324096 152998
rect 324044 152934 324096 152940
rect 324056 150226 324084 152934
rect 324700 150226 324728 157762
rect 325332 154352 325384 154358
rect 325332 154294 325384 154300
rect 325344 150226 325372 154294
rect 327000 154290 327028 163254
rect 327538 163200 327594 164400
rect 328366 163200 328422 164400
rect 329194 163200 329250 164400
rect 330114 163200 330170 164400
rect 330942 163200 330998 164400
rect 331770 163200 331826 164400
rect 332598 163200 332654 164400
rect 333426 163200 333482 164400
rect 334254 163200 334310 164400
rect 335082 163200 335138 164400
rect 336002 163200 336058 164400
rect 336830 163200 336886 164400
rect 337658 163200 337714 164400
rect 337764 163254 338068 163282
rect 327552 158982 327580 163200
rect 328380 161474 328408 163200
rect 328288 161446 328408 161474
rect 329208 161474 329236 163200
rect 329208 161446 329328 161474
rect 327540 158976 327592 158982
rect 327540 158918 327592 158924
rect 327080 158500 327132 158506
rect 327080 158442 327132 158448
rect 326988 154284 327040 154290
rect 326988 154226 327040 154232
rect 325976 153604 326028 153610
rect 325976 153546 326028 153552
rect 325988 150226 326016 153546
rect 326620 151904 326672 151910
rect 326620 151846 326672 151852
rect 326632 150226 326660 151846
rect 327092 151814 327120 158442
rect 327908 155712 327960 155718
rect 327908 155654 327960 155660
rect 327092 151786 327304 151814
rect 327276 150226 327304 151786
rect 327920 150226 327948 155654
rect 328288 152930 328316 161446
rect 328368 158976 328420 158982
rect 328368 158918 328420 158924
rect 328380 155718 328408 158918
rect 328552 158568 328604 158574
rect 328552 158510 328604 158516
rect 328368 155712 328420 155718
rect 328368 155654 328420 155660
rect 328276 152924 328328 152930
rect 328276 152866 328328 152872
rect 328564 150226 328592 158510
rect 329300 152658 329328 161446
rect 330128 158438 330156 163200
rect 330208 159996 330260 160002
rect 330208 159938 330260 159944
rect 330116 158432 330168 158438
rect 330116 158374 330168 158380
rect 329840 157276 329892 157282
rect 329840 157218 329892 157224
rect 329196 152652 329248 152658
rect 329196 152594 329248 152600
rect 329288 152652 329340 152658
rect 329288 152594 329340 152600
rect 329208 150226 329236 152594
rect 329852 150226 329880 157218
rect 330220 155174 330248 159938
rect 330956 157010 330984 163200
rect 331784 159390 331812 163200
rect 332612 160002 332640 163200
rect 332600 159996 332652 160002
rect 332600 159938 332652 159944
rect 332600 159656 332652 159662
rect 332600 159598 332652 159604
rect 331772 159384 331824 159390
rect 331772 159326 331824 159332
rect 331772 158908 331824 158914
rect 331772 158850 331824 158856
rect 331312 158636 331364 158642
rect 331312 158578 331364 158584
rect 330944 157004 330996 157010
rect 330944 156946 330996 156952
rect 330484 155644 330536 155650
rect 330484 155586 330536 155592
rect 330208 155168 330260 155174
rect 330208 155110 330260 155116
rect 330024 155100 330076 155106
rect 330024 155042 330076 155048
rect 323412 150198 323486 150226
rect 324056 150198 324130 150226
rect 324700 150198 324774 150226
rect 325344 150198 325418 150226
rect 325988 150198 326062 150226
rect 326632 150198 326706 150226
rect 327276 150198 327350 150226
rect 327920 150198 327994 150226
rect 328564 150198 328638 150226
rect 329208 150198 329282 150226
rect 329852 150198 329926 150226
rect 330036 150210 330064 155042
rect 330496 150226 330524 155586
rect 322814 149940 322842 150198
rect 323458 149940 323486 150198
rect 324102 149940 324130 150198
rect 324746 149940 324774 150198
rect 325390 149940 325418 150198
rect 326034 149940 326062 150198
rect 326678 149940 326706 150198
rect 327322 149940 327350 150198
rect 327966 149940 327994 150198
rect 328610 149940 328638 150198
rect 329254 149940 329282 150198
rect 329898 149940 329926 150198
rect 330024 150204 330076 150210
rect 330496 150198 330570 150226
rect 331324 150210 331352 158578
rect 331784 150226 331812 158850
rect 332612 151910 332640 159598
rect 333060 155780 333112 155786
rect 333060 155722 333112 155728
rect 332600 151904 332652 151910
rect 332600 151846 332652 151852
rect 333072 150226 333100 155722
rect 333440 154358 333468 163200
rect 334268 155650 334296 163200
rect 334900 156732 334952 156738
rect 334900 156674 334952 156680
rect 334256 155644 334308 155650
rect 334256 155586 334308 155592
rect 333704 154420 333756 154426
rect 333704 154362 333756 154368
rect 333428 154352 333480 154358
rect 333428 154294 333480 154300
rect 333716 150226 333744 154362
rect 334348 153196 334400 153202
rect 334348 153138 334400 153144
rect 334360 150226 334388 153138
rect 334912 150226 334940 156674
rect 335096 154426 335124 163200
rect 336016 158778 336044 163200
rect 336648 160064 336700 160070
rect 336648 160006 336700 160012
rect 336004 158772 336056 158778
rect 336004 158714 336056 158720
rect 336660 155786 336688 160006
rect 336844 157078 336872 163200
rect 337672 163146 337700 163200
rect 337764 163146 337792 163254
rect 337672 163118 337792 163146
rect 337752 158772 337804 158778
rect 337752 158714 337804 158720
rect 336832 157072 336884 157078
rect 336832 157014 336884 157020
rect 336648 155780 336700 155786
rect 336648 155722 336700 155728
rect 335544 155236 335596 155242
rect 335544 155178 335596 155184
rect 335084 154420 335136 154426
rect 335084 154362 335136 154368
rect 335556 150226 335584 155178
rect 337476 153944 337528 153950
rect 337476 153886 337528 153892
rect 336188 153808 336240 153814
rect 336188 153750 336240 153756
rect 336200 150226 336228 153750
rect 336832 151904 336884 151910
rect 336832 151846 336884 151852
rect 336844 150226 336872 151846
rect 337488 150226 337516 153886
rect 337764 152998 337792 158714
rect 338040 153950 338068 163254
rect 338486 163200 338542 164400
rect 339314 163200 339370 164400
rect 340142 163200 340198 164400
rect 340970 163200 341026 164400
rect 341890 163200 341946 164400
rect 342718 163200 342774 164400
rect 343546 163200 343602 164400
rect 344374 163200 344430 164400
rect 345202 163200 345258 164400
rect 346030 163200 346086 164400
rect 346858 163200 346914 164400
rect 347778 163200 347834 164400
rect 348606 163200 348662 164400
rect 349434 163200 349490 164400
rect 350262 163200 350318 164400
rect 351090 163200 351146 164400
rect 351918 163200 351974 164400
rect 352746 163200 352802 164400
rect 353666 163200 353722 164400
rect 354494 163200 354550 164400
rect 355322 163200 355378 164400
rect 356150 163200 356206 164400
rect 356978 163200 357034 164400
rect 357084 163254 357388 163282
rect 338396 159724 338448 159730
rect 338396 159666 338448 159672
rect 338120 155304 338172 155310
rect 338120 155246 338172 155252
rect 338028 153944 338080 153950
rect 338028 153886 338080 153892
rect 337752 152992 337804 152998
rect 337752 152934 337804 152940
rect 338132 150226 338160 155246
rect 338408 154562 338436 159666
rect 338500 158506 338528 163200
rect 339328 159594 339356 163200
rect 339316 159588 339368 159594
rect 339316 159530 339368 159536
rect 338488 158500 338540 158506
rect 338488 158442 338540 158448
rect 340156 158030 340184 163200
rect 340052 158024 340104 158030
rect 340052 157966 340104 157972
rect 340144 158024 340196 158030
rect 340144 157966 340196 157972
rect 338672 157208 338724 157214
rect 338672 157150 338724 157156
rect 338396 154556 338448 154562
rect 338396 154498 338448 154504
rect 338684 151814 338712 157150
rect 339592 155372 339644 155378
rect 339592 155314 339644 155320
rect 338948 154420 339000 154426
rect 338948 154362 339000 154368
rect 338960 153202 338988 154362
rect 338948 153196 339000 153202
rect 338948 153138 339000 153144
rect 339408 153128 339460 153134
rect 339408 153070 339460 153076
rect 338684 151786 338804 151814
rect 338776 150226 338804 151786
rect 339420 150226 339448 153070
rect 330024 150146 330076 150152
rect 330542 149940 330570 150198
rect 331174 150204 331226 150210
rect 331174 150146 331226 150152
rect 331312 150204 331364 150210
rect 331784 150198 331858 150226
rect 331312 150146 331364 150152
rect 331186 149940 331214 150146
rect 331830 149940 331858 150198
rect 332462 150204 332514 150210
rect 333072 150198 333146 150226
rect 333716 150198 333790 150226
rect 334360 150198 334434 150226
rect 334912 150198 334986 150226
rect 335556 150198 335630 150226
rect 336200 150198 336274 150226
rect 336844 150198 336918 150226
rect 337488 150198 337562 150226
rect 338132 150198 338206 150226
rect 338776 150198 338850 150226
rect 339420 150198 339494 150226
rect 339604 150210 339632 155314
rect 340064 150226 340092 157966
rect 340984 154426 341012 163200
rect 341340 157752 341392 157758
rect 341340 157694 341392 157700
rect 340972 154420 341024 154426
rect 340972 154362 341024 154368
rect 341352 150226 341380 157694
rect 341904 156738 341932 163200
rect 342732 160070 342760 163200
rect 342720 160064 342772 160070
rect 342720 160006 342772 160012
rect 342260 158092 342312 158098
rect 342260 158034 342312 158040
rect 341892 156732 341944 156738
rect 341892 156674 341944 156680
rect 341984 154556 342036 154562
rect 341984 154498 342036 154504
rect 341996 150226 342024 154498
rect 342272 151814 342300 158034
rect 343272 155508 343324 155514
rect 343272 155450 343324 155456
rect 342272 151786 342668 151814
rect 342640 150226 342668 151786
rect 343284 150226 343312 155450
rect 343560 155242 343588 163200
rect 343640 159792 343692 159798
rect 343640 159734 343692 159740
rect 343548 155236 343600 155242
rect 343548 155178 343600 155184
rect 343652 151910 343680 159734
rect 343916 155576 343968 155582
rect 343916 155518 343968 155524
rect 343640 151904 343692 151910
rect 343640 151846 343692 151852
rect 343928 150226 343956 155518
rect 344388 155310 344416 163200
rect 345020 157344 345072 157350
rect 345020 157286 345072 157292
rect 344376 155304 344428 155310
rect 344376 155246 344428 155252
rect 344560 152720 344612 152726
rect 344560 152662 344612 152668
rect 344572 150226 344600 152662
rect 345032 151814 345060 157286
rect 345216 155378 345244 163200
rect 345940 159860 345992 159866
rect 345940 159802 345992 159808
rect 345952 155854 345980 159802
rect 346044 159730 346072 163200
rect 346032 159724 346084 159730
rect 346032 159666 346084 159672
rect 346872 157146 346900 163200
rect 347792 157214 347820 163200
rect 347780 157208 347832 157214
rect 347780 157150 347832 157156
rect 346860 157140 346912 157146
rect 346860 157082 346912 157088
rect 348620 156670 348648 163200
rect 349252 156800 349304 156806
rect 349252 156742 349304 156748
rect 347780 156664 347832 156670
rect 347780 156606 347832 156612
rect 348608 156664 348660 156670
rect 348608 156606 348660 156612
rect 346492 156460 346544 156466
rect 346492 156402 346544 156408
rect 345848 155848 345900 155854
rect 345848 155790 345900 155796
rect 345940 155848 345992 155854
rect 345940 155790 345992 155796
rect 345204 155372 345256 155378
rect 345204 155314 345256 155320
rect 345032 151786 345244 151814
rect 345216 150226 345244 151786
rect 345860 150226 345888 155790
rect 346504 150226 346532 156402
rect 347136 151904 347188 151910
rect 347136 151846 347188 151852
rect 347148 150226 347176 151846
rect 347792 150226 347820 156606
rect 348424 155440 348476 155446
rect 348424 155382 348476 155388
rect 348436 150226 348464 155382
rect 349068 154012 349120 154018
rect 349068 153954 349120 153960
rect 349080 150226 349108 153954
rect 332462 150146 332514 150152
rect 332474 149940 332502 150146
rect 333118 149940 333146 150198
rect 333762 149940 333790 150198
rect 334406 149940 334434 150198
rect 334958 149940 334986 150198
rect 335602 149940 335630 150198
rect 336246 149940 336274 150198
rect 336890 149940 336918 150198
rect 337534 149940 337562 150198
rect 338178 149940 338206 150198
rect 338822 149940 338850 150198
rect 339466 149940 339494 150198
rect 339592 150204 339644 150210
rect 340064 150198 340138 150226
rect 339592 150146 339644 150152
rect 340110 149940 340138 150198
rect 340742 150204 340794 150210
rect 341352 150198 341426 150226
rect 341996 150198 342070 150226
rect 342640 150198 342714 150226
rect 343284 150198 343358 150226
rect 343928 150198 344002 150226
rect 344572 150198 344646 150226
rect 345216 150198 345290 150226
rect 345860 150198 345934 150226
rect 346504 150198 346578 150226
rect 347148 150198 347222 150226
rect 347792 150198 347866 150226
rect 348436 150198 348510 150226
rect 349080 150198 349154 150226
rect 349264 150210 349292 156742
rect 349448 152454 349476 163200
rect 350276 158098 350304 163200
rect 351104 158574 351132 163200
rect 351932 158642 351960 163200
rect 352760 159662 352788 163200
rect 352748 159656 352800 159662
rect 352748 159598 352800 159604
rect 352012 159316 352064 159322
rect 352012 159258 352064 159264
rect 351920 158636 351972 158642
rect 351920 158578 351972 158584
rect 351092 158568 351144 158574
rect 351092 158510 351144 158516
rect 350264 158092 350316 158098
rect 350264 158034 350316 158040
rect 350540 157956 350592 157962
rect 350540 157898 350592 157904
rect 349712 152516 349764 152522
rect 349712 152458 349764 152464
rect 349436 152448 349488 152454
rect 349436 152390 349488 152396
rect 349724 150226 349752 152458
rect 340742 150146 340794 150152
rect 340754 149940 340782 150146
rect 341398 149940 341426 150198
rect 342042 149940 342070 150198
rect 342686 149940 342714 150198
rect 343330 149940 343358 150198
rect 343974 149940 344002 150198
rect 344618 149940 344646 150198
rect 345262 149940 345290 150198
rect 345906 149940 345934 150198
rect 346550 149940 346578 150198
rect 347194 149940 347222 150198
rect 347838 149940 347866 150198
rect 348482 149940 348510 150198
rect 349126 149940 349154 150198
rect 349252 150204 349304 150210
rect 349724 150198 349798 150226
rect 350552 150210 350580 157898
rect 352024 157282 352052 159258
rect 353300 158160 353352 158166
rect 353300 158102 353352 158108
rect 352012 157276 352064 157282
rect 352012 157218 352064 157224
rect 351920 156868 351972 156874
rect 351920 156810 351972 156816
rect 351000 156596 351052 156602
rect 351000 156538 351052 156544
rect 351012 150226 351040 156538
rect 349252 150146 349304 150152
rect 349770 149940 349798 150198
rect 350402 150204 350454 150210
rect 350402 150146 350454 150152
rect 350540 150204 350592 150210
rect 351012 150198 351086 150226
rect 351932 150210 351960 156810
rect 352288 155848 352340 155854
rect 352288 155790 352340 155796
rect 352300 150226 352328 155790
rect 353312 151814 353340 158102
rect 353680 155514 353708 163200
rect 354220 156528 354272 156534
rect 354220 156470 354272 156476
rect 353668 155508 353720 155514
rect 353668 155450 353720 155456
rect 353312 151786 353616 151814
rect 353588 150226 353616 151786
rect 354232 150226 354260 156470
rect 354508 155446 354536 163200
rect 354496 155440 354548 155446
rect 354496 155382 354548 155388
rect 355336 153814 355364 163200
rect 355692 159452 355744 159458
rect 355692 159394 355744 159400
rect 355508 153876 355560 153882
rect 355508 153818 355560 153824
rect 355324 153808 355376 153814
rect 355324 153750 355376 153756
rect 354864 152788 354916 152794
rect 354864 152730 354916 152736
rect 354876 150226 354904 152730
rect 355520 150226 355548 153818
rect 355704 153202 355732 159394
rect 356164 157350 356192 163200
rect 356992 163146 357020 163200
rect 357084 163146 357112 163254
rect 356992 163118 357112 163146
rect 356152 157344 356204 157350
rect 356152 157286 356204 157292
rect 356152 156936 356204 156942
rect 356152 156878 356204 156884
rect 355692 153196 355744 153202
rect 355692 153138 355744 153144
rect 356164 150226 356192 156878
rect 356796 155168 356848 155174
rect 356796 155110 356848 155116
rect 356808 150226 356836 155110
rect 357360 153882 357388 163254
rect 357806 163200 357862 164400
rect 358634 163200 358690 164400
rect 359554 163200 359610 164400
rect 360382 163200 360438 164400
rect 361210 163200 361266 164400
rect 362038 163200 362094 164400
rect 362866 163200 362922 164400
rect 363694 163200 363750 164400
rect 364522 163200 364578 164400
rect 365442 163200 365498 164400
rect 366270 163200 366326 164400
rect 367098 163200 367154 164400
rect 367926 163200 367982 164400
rect 368032 163254 368428 163282
rect 357624 158228 357676 158234
rect 357624 158170 357676 158176
rect 357348 153876 357400 153882
rect 357348 153818 357400 153824
rect 357440 153196 357492 153202
rect 357440 153138 357492 153144
rect 357452 150226 357480 153138
rect 350540 150146 350592 150152
rect 350414 149940 350442 150146
rect 351058 149940 351086 150198
rect 351690 150204 351742 150210
rect 351690 150146 351742 150152
rect 351920 150204 351972 150210
rect 352300 150198 352374 150226
rect 351920 150146 351972 150152
rect 351702 149940 351730 150146
rect 352346 149940 352374 150198
rect 352978 150204 353030 150210
rect 353588 150198 353662 150226
rect 354232 150198 354306 150226
rect 354876 150198 354950 150226
rect 355520 150198 355594 150226
rect 356164 150198 356238 150226
rect 356808 150198 356882 150226
rect 357452 150198 357526 150226
rect 357636 150210 357664 158170
rect 357820 156806 357848 163200
rect 358648 158166 358676 163200
rect 359568 159458 359596 163200
rect 359556 159452 359608 159458
rect 359556 159394 359608 159400
rect 359464 158704 359516 158710
rect 359464 158646 359516 158652
rect 358636 158160 358688 158166
rect 358636 158102 358688 158108
rect 358912 157344 358964 157350
rect 358912 157286 358964 157292
rect 357808 156800 357860 156806
rect 357808 156742 357860 156748
rect 358084 154488 358136 154494
rect 358084 154430 358136 154436
rect 358096 150226 358124 154430
rect 358924 152794 358952 157286
rect 358912 152788 358964 152794
rect 358912 152730 358964 152736
rect 359372 152584 359424 152590
rect 359372 152526 359424 152532
rect 359384 150226 359412 152526
rect 359476 151910 359504 158646
rect 360200 158296 360252 158302
rect 360200 158238 360252 158244
rect 360016 153060 360068 153066
rect 360016 153002 360068 153008
rect 359464 151904 359516 151910
rect 359464 151846 359516 151852
rect 360028 150226 360056 153002
rect 352978 150146 353030 150152
rect 352990 149940 353018 150146
rect 353634 149940 353662 150198
rect 354278 149940 354306 150198
rect 354922 149940 354950 150198
rect 355566 149940 355594 150198
rect 356210 149940 356238 150198
rect 356854 149940 356882 150198
rect 357498 149940 357526 150198
rect 357624 150204 357676 150210
rect 358096 150198 358170 150226
rect 357624 150146 357676 150152
rect 358142 149940 358170 150198
rect 358774 150204 358826 150210
rect 359384 150198 359458 150226
rect 360028 150198 360102 150226
rect 360212 150210 360240 158238
rect 360396 154018 360424 163200
rect 361224 158234 361252 163200
rect 361580 159520 361632 159526
rect 361580 159462 361632 159468
rect 361212 158228 361264 158234
rect 361212 158170 361264 158176
rect 360660 154080 360712 154086
rect 360660 154022 360712 154028
rect 360384 154012 360436 154018
rect 360384 153954 360436 153960
rect 360672 150226 360700 154022
rect 360844 153944 360896 153950
rect 361028 153944 361080 153950
rect 360896 153892 361028 153898
rect 360844 153886 361080 153892
rect 360856 153870 361068 153886
rect 358774 150146 358826 150152
rect 358786 149940 358814 150146
rect 359430 149940 359458 150198
rect 360074 149940 360102 150198
rect 360200 150204 360252 150210
rect 360672 150198 360746 150226
rect 361592 150210 361620 159462
rect 362052 158982 362080 163200
rect 362132 159928 362184 159934
rect 362132 159870 362184 159876
rect 362040 158976 362092 158982
rect 362040 158918 362092 158924
rect 362144 155786 362172 159870
rect 362880 158794 362908 163200
rect 362880 158766 363000 158794
rect 361948 155780 362000 155786
rect 361948 155722 362000 155728
rect 362132 155780 362184 155786
rect 362132 155722 362184 155728
rect 361960 150226 361988 155722
rect 362972 152726 363000 158766
rect 363512 158364 363564 158370
rect 363512 158306 363564 158312
rect 363236 154148 363288 154154
rect 363236 154090 363288 154096
rect 362960 152720 363012 152726
rect 362960 152662 363012 152668
rect 363248 150226 363276 154090
rect 363524 151814 363552 158306
rect 363708 156874 363736 163200
rect 363696 156868 363748 156874
rect 363696 156810 363748 156816
rect 364536 155582 364564 163200
rect 364524 155576 364576 155582
rect 364524 155518 364576 155524
rect 365168 152856 365220 152862
rect 365168 152798 365220 152804
rect 364524 151904 364576 151910
rect 364524 151846 364576 151852
rect 363524 151786 363920 151814
rect 363892 150226 363920 151786
rect 364536 150226 364564 151846
rect 365180 150226 365208 152798
rect 365456 152590 365484 163200
rect 366284 159526 366312 163200
rect 366272 159520 366324 159526
rect 366272 159462 366324 159468
rect 366824 158976 366876 158982
rect 366824 158918 366876 158924
rect 365904 157276 365956 157282
rect 365904 157218 365956 157224
rect 365720 154216 365772 154222
rect 365720 154158 365772 154164
rect 365444 152584 365496 152590
rect 365444 152526 365496 152532
rect 365732 150226 365760 154158
rect 360200 150146 360252 150152
rect 360718 149940 360746 150198
rect 361350 150204 361402 150210
rect 361350 150146 361402 150152
rect 361580 150204 361632 150210
rect 361960 150198 362034 150226
rect 361580 150146 361632 150152
rect 361362 149940 361390 150146
rect 362006 149940 362034 150198
rect 362638 150204 362690 150210
rect 363248 150198 363322 150226
rect 363892 150198 363966 150226
rect 364536 150198 364610 150226
rect 365180 150198 365254 150226
rect 365732 150198 365806 150226
rect 365916 150210 365944 157218
rect 366272 155916 366324 155922
rect 366272 155858 366324 155864
rect 366284 151814 366312 155858
rect 366836 154494 366864 158918
rect 367112 158302 367140 163200
rect 367940 163146 367968 163200
rect 368032 163146 368060 163254
rect 367940 163118 368060 163146
rect 367100 158296 367152 158302
rect 367100 158238 367152 158244
rect 367652 155780 367704 155786
rect 367652 155722 367704 155728
rect 366824 154488 366876 154494
rect 366824 154430 366876 154436
rect 366284 151786 366404 151814
rect 366376 150226 366404 151786
rect 367664 150226 367692 155722
rect 368296 154284 368348 154290
rect 368296 154226 368348 154232
rect 368308 150226 368336 154226
rect 368400 154154 368428 163254
rect 368754 163200 368810 164400
rect 369582 163200 369638 164400
rect 370410 163200 370466 164400
rect 371330 163200 371386 164400
rect 372158 163200 372214 164400
rect 372986 163200 373042 164400
rect 373814 163200 373870 164400
rect 374642 163200 374698 164400
rect 375470 163200 375526 164400
rect 376298 163200 376354 164400
rect 376404 163254 376708 163282
rect 368572 159996 368624 160002
rect 368572 159938 368624 159944
rect 368388 154148 368440 154154
rect 368388 154090 368440 154096
rect 368584 153202 368612 159938
rect 368768 159798 368796 163200
rect 368756 159792 368808 159798
rect 368756 159734 368808 159740
rect 369596 155718 369624 163200
rect 370424 155786 370452 163200
rect 370872 158432 370924 158438
rect 370872 158374 370924 158380
rect 370412 155780 370464 155786
rect 370412 155722 370464 155728
rect 368940 155712 368992 155718
rect 368940 155654 368992 155660
rect 369584 155712 369636 155718
rect 369584 155654 369636 155660
rect 368572 153196 368624 153202
rect 368572 153138 368624 153144
rect 368952 150226 368980 155654
rect 369584 152924 369636 152930
rect 369584 152866 369636 152872
rect 369596 150226 369624 152866
rect 370228 152652 370280 152658
rect 370228 152594 370280 152600
rect 370240 150226 370268 152594
rect 370884 150226 370912 158374
rect 371240 157004 371292 157010
rect 371240 156946 371292 156952
rect 371252 151814 371280 156946
rect 371344 154222 371372 163200
rect 372068 159384 372120 159390
rect 372068 159326 372120 159332
rect 371332 154216 371384 154222
rect 371332 154158 371384 154164
rect 372080 151814 372108 159326
rect 372172 158982 372200 163200
rect 372620 160064 372672 160070
rect 372620 160006 372672 160012
rect 372160 158976 372212 158982
rect 372160 158918 372212 158924
rect 372632 152930 372660 160006
rect 373000 159390 373028 163200
rect 372988 159384 373040 159390
rect 372988 159326 373040 159332
rect 373828 156942 373856 163200
rect 374276 158976 374328 158982
rect 374276 158918 374328 158924
rect 373816 156936 373868 156942
rect 373816 156878 373868 156884
rect 374092 155644 374144 155650
rect 374092 155586 374144 155592
rect 373448 154352 373500 154358
rect 373448 154294 373500 154300
rect 372804 153196 372856 153202
rect 372804 153138 372856 153144
rect 372620 152924 372672 152930
rect 372620 152866 372672 152872
rect 371252 151786 371556 151814
rect 372080 151786 372200 151814
rect 371528 150226 371556 151786
rect 372172 150226 372200 151786
rect 372816 150226 372844 153138
rect 373460 150226 373488 154294
rect 374104 150226 374132 155586
rect 374288 152862 374316 158918
rect 374656 157010 374684 163200
rect 375484 159866 375512 163200
rect 376312 163146 376340 163200
rect 376404 163146 376432 163254
rect 376312 163118 376432 163146
rect 375472 159860 375524 159866
rect 375472 159802 375524 159808
rect 376024 157072 376076 157078
rect 376024 157014 376076 157020
rect 374644 157004 374696 157010
rect 374644 156946 374696 156952
rect 374736 153128 374788 153134
rect 374736 153070 374788 153076
rect 374276 152856 374328 152862
rect 374276 152798 374328 152804
rect 374748 150226 374776 153070
rect 375380 152992 375432 152998
rect 375380 152934 375432 152940
rect 375392 150226 375420 152934
rect 376036 150226 376064 157014
rect 376576 153944 376628 153950
rect 376576 153886 376628 153892
rect 376588 151814 376616 153886
rect 376680 152658 376708 163254
rect 377218 163200 377274 164400
rect 378046 163200 378102 164400
rect 378874 163200 378930 164400
rect 379702 163200 379758 164400
rect 380530 163200 380586 164400
rect 380636 163254 380848 163282
rect 377232 158506 377260 163200
rect 377956 159588 378008 159594
rect 377956 159530 378008 159536
rect 376852 158500 376904 158506
rect 376852 158442 376904 158448
rect 377220 158500 377272 158506
rect 377220 158442 377272 158448
rect 376668 152652 376720 152658
rect 376668 152594 376720 152600
rect 376864 151814 376892 158442
rect 376588 151786 376708 151814
rect 376864 151786 377352 151814
rect 376680 150226 376708 151786
rect 377324 150226 377352 151786
rect 377968 150226 377996 159530
rect 378060 158370 378088 163200
rect 378324 159724 378376 159730
rect 378324 159666 378376 159672
rect 378048 158364 378100 158370
rect 378048 158306 378100 158312
rect 378336 155650 378364 159666
rect 378888 158846 378916 163200
rect 379716 159594 379744 163200
rect 380544 163146 380572 163200
rect 380636 163146 380664 163254
rect 380544 163118 380664 163146
rect 379704 159588 379756 159594
rect 379704 159530 379756 159536
rect 378876 158840 378928 158846
rect 378876 158782 378928 158788
rect 378600 158024 378652 158030
rect 378600 157966 378652 157972
rect 378324 155644 378376 155650
rect 378324 155586 378376 155592
rect 378612 150226 378640 157966
rect 379888 156732 379940 156738
rect 379888 156674 379940 156680
rect 379244 154420 379296 154426
rect 379244 154362 379296 154368
rect 379256 150226 379284 154362
rect 379900 150226 379928 156674
rect 380820 153950 380848 163254
rect 381358 163200 381414 164400
rect 382186 163200 382242 164400
rect 383106 163200 383162 164400
rect 383934 163200 383990 164400
rect 384762 163200 384818 164400
rect 385590 163200 385646 164400
rect 386418 163200 386474 164400
rect 387246 163200 387302 164400
rect 388074 163200 388130 164400
rect 388994 163200 389050 164400
rect 389822 163200 389878 164400
rect 390650 163200 390706 164400
rect 391478 163200 391534 164400
rect 391584 163254 391796 163282
rect 380992 158840 381044 158846
rect 380992 158782 381044 158788
rect 380900 155236 380952 155242
rect 380900 155178 380952 155184
rect 380808 153944 380860 153950
rect 380808 153886 380860 153892
rect 380532 152924 380584 152930
rect 380532 152866 380584 152872
rect 380544 150226 380572 152866
rect 380912 151814 380940 155178
rect 381004 152930 381032 158782
rect 381372 155242 381400 163200
rect 382200 159730 382228 163200
rect 382188 159724 382240 159730
rect 382188 159666 382240 159672
rect 383120 157078 383148 163200
rect 383660 157208 383712 157214
rect 383660 157150 383712 157156
rect 383108 157072 383160 157078
rect 383108 157014 383160 157020
rect 383108 155644 383160 155650
rect 383108 155586 383160 155592
rect 382280 155372 382332 155378
rect 382280 155314 382332 155320
rect 381452 155304 381504 155310
rect 381452 155246 381504 155252
rect 381360 155236 381412 155242
rect 381360 155178 381412 155184
rect 380992 152924 381044 152930
rect 380992 152866 381044 152872
rect 381464 151814 381492 155246
rect 382292 151814 382320 155314
rect 380912 151786 381216 151814
rect 381464 151786 381860 151814
rect 382292 151786 382504 151814
rect 381188 150226 381216 151786
rect 381832 150226 381860 151786
rect 382476 150226 382504 151786
rect 383120 150226 383148 155586
rect 362638 150146 362690 150152
rect 362650 149940 362678 150146
rect 363294 149940 363322 150198
rect 363938 149940 363966 150198
rect 364582 149940 364610 150198
rect 365226 149940 365254 150198
rect 365778 149940 365806 150198
rect 365904 150204 365956 150210
rect 366376 150198 366450 150226
rect 365904 150146 365956 150152
rect 366422 149940 366450 150198
rect 367054 150204 367106 150210
rect 367664 150198 367738 150226
rect 368308 150198 368382 150226
rect 368952 150198 369026 150226
rect 369596 150198 369670 150226
rect 370240 150198 370314 150226
rect 370884 150198 370958 150226
rect 371528 150198 371602 150226
rect 372172 150198 372246 150226
rect 372816 150198 372890 150226
rect 373460 150198 373534 150226
rect 374104 150198 374178 150226
rect 374748 150198 374822 150226
rect 375392 150198 375466 150226
rect 376036 150198 376110 150226
rect 376680 150198 376754 150226
rect 377324 150198 377398 150226
rect 377968 150198 378042 150226
rect 378612 150198 378686 150226
rect 379256 150198 379330 150226
rect 379900 150198 379974 150226
rect 380544 150198 380618 150226
rect 381188 150198 381262 150226
rect 381832 150198 381906 150226
rect 382476 150198 382550 150226
rect 383120 150198 383194 150226
rect 383672 150210 383700 157150
rect 383752 157140 383804 157146
rect 383752 157082 383804 157088
rect 383764 150226 383792 157082
rect 383948 155310 383976 163200
rect 384776 156738 384804 163200
rect 385604 158778 385632 163200
rect 386432 160002 386460 163200
rect 386420 159996 386472 160002
rect 386420 159938 386472 159944
rect 385960 159656 386012 159662
rect 385960 159598 386012 159604
rect 385592 158772 385644 158778
rect 385592 158714 385644 158720
rect 385224 158092 385276 158098
rect 385224 158034 385276 158040
rect 384764 156732 384816 156738
rect 384764 156674 384816 156680
rect 385040 156664 385092 156670
rect 385040 156606 385092 156612
rect 383936 155304 383988 155310
rect 383936 155246 383988 155252
rect 385052 150226 385080 156606
rect 367054 150146 367106 150152
rect 367066 149940 367094 150146
rect 367710 149940 367738 150198
rect 368354 149940 368382 150198
rect 368998 149940 369026 150198
rect 369642 149940 369670 150198
rect 370286 149940 370314 150198
rect 370930 149940 370958 150198
rect 371574 149940 371602 150198
rect 372218 149940 372246 150198
rect 372862 149940 372890 150198
rect 373506 149940 373534 150198
rect 374150 149940 374178 150198
rect 374794 149940 374822 150198
rect 375438 149940 375466 150198
rect 376082 149940 376110 150198
rect 376726 149940 376754 150198
rect 377370 149940 377398 150198
rect 378014 149940 378042 150198
rect 378658 149940 378686 150198
rect 379302 149940 379330 150198
rect 379946 149940 379974 150198
rect 380590 149940 380618 150198
rect 381234 149940 381262 150198
rect 381878 149940 381906 150198
rect 382522 149940 382550 150198
rect 383166 149940 383194 150198
rect 383660 150204 383712 150210
rect 383764 150198 383838 150226
rect 383660 150146 383712 150152
rect 383810 149940 383838 150198
rect 384442 150204 384494 150210
rect 385052 150198 385126 150226
rect 385236 150210 385264 158034
rect 385972 153202 386000 159598
rect 386512 158636 386564 158642
rect 386512 158578 386564 158584
rect 385960 153196 386012 153202
rect 385960 153138 386012 153144
rect 385592 152516 385644 152522
rect 385592 152458 385644 152464
rect 385604 151814 385632 152458
rect 385604 151786 385724 151814
rect 385696 150226 385724 151786
rect 384442 150146 384494 150152
rect 384454 149940 384482 150146
rect 385098 149940 385126 150198
rect 385224 150204 385276 150210
rect 385696 150198 385770 150226
rect 386524 150210 386552 158578
rect 386972 158568 387024 158574
rect 386972 158510 387024 158516
rect 386984 150226 387012 158510
rect 387260 156670 387288 163200
rect 388088 158030 388116 163200
rect 389008 159662 389036 163200
rect 388996 159656 389048 159662
rect 388996 159598 389048 159604
rect 389836 158846 389864 163200
rect 390664 159050 390692 163200
rect 391492 163146 391520 163200
rect 391584 163146 391612 163254
rect 391492 163118 391612 163146
rect 390652 159044 390704 159050
rect 390652 158986 390704 158992
rect 389824 158840 389876 158846
rect 389824 158782 389876 158788
rect 391572 158840 391624 158846
rect 391572 158782 391624 158788
rect 389088 158772 389140 158778
rect 389088 158714 389140 158720
rect 388076 158024 388128 158030
rect 388076 157966 388128 157972
rect 387248 156664 387300 156670
rect 387248 156606 387300 156612
rect 388352 155508 388404 155514
rect 388352 155450 388404 155456
rect 388260 153196 388312 153202
rect 388260 153138 388312 153144
rect 388272 150226 388300 153138
rect 388364 151814 388392 155450
rect 389100 152998 389128 158714
rect 389548 155440 389600 155446
rect 389548 155382 389600 155388
rect 389088 152992 389140 152998
rect 389088 152934 389140 152940
rect 388364 151786 388944 151814
rect 388916 150226 388944 151786
rect 389560 150226 389588 155382
rect 391480 154012 391532 154018
rect 391480 153954 391532 153960
rect 390192 153876 390244 153882
rect 390192 153818 390244 153824
rect 390204 150226 390232 153818
rect 390836 152788 390888 152794
rect 390836 152730 390888 152736
rect 390848 150226 390876 152730
rect 391492 150226 391520 153954
rect 391584 152794 391612 158782
rect 391768 153882 391796 163254
rect 392306 163200 392362 164400
rect 393134 163200 393190 164400
rect 393962 163200 394018 164400
rect 394882 163200 394938 164400
rect 395710 163200 395766 164400
rect 396538 163200 396594 164400
rect 397366 163200 397422 164400
rect 398194 163200 398250 164400
rect 399022 163200 399078 164400
rect 399850 163200 399906 164400
rect 400770 163200 400826 164400
rect 401598 163200 401654 164400
rect 402426 163200 402482 164400
rect 403254 163200 403310 164400
rect 404082 163200 404138 164400
rect 404910 163200 404966 164400
rect 405738 163200 405794 164400
rect 406658 163200 406714 164400
rect 407486 163200 407542 164400
rect 408314 163200 408370 164400
rect 409142 163200 409198 164400
rect 409970 163200 410026 164400
rect 410798 163200 410854 164400
rect 411626 163200 411682 164400
rect 412546 163200 412602 164400
rect 413374 163200 413430 164400
rect 414202 163200 414258 164400
rect 415030 163200 415086 164400
rect 415858 163200 415914 164400
rect 416686 163200 416742 164400
rect 417514 163200 417570 164400
rect 418434 163200 418490 164400
rect 419262 163200 419318 164400
rect 420090 163200 420146 164400
rect 420918 163200 420974 164400
rect 421746 163200 421802 164400
rect 422574 163200 422630 164400
rect 423402 163200 423458 164400
rect 424322 163200 424378 164400
rect 425150 163200 425206 164400
rect 425978 163200 426034 164400
rect 426806 163200 426862 164400
rect 427634 163200 427690 164400
rect 428462 163200 428518 164400
rect 429290 163200 429346 164400
rect 430210 163200 430266 164400
rect 431038 163200 431094 164400
rect 431866 163200 431922 164400
rect 432694 163200 432750 164400
rect 433522 163200 433578 164400
rect 434350 163200 434406 164400
rect 435178 163200 435234 164400
rect 436098 163200 436154 164400
rect 436926 163200 436982 164400
rect 437032 163254 437428 163282
rect 391848 159044 391900 159050
rect 391848 158986 391900 158992
rect 391860 154018 391888 158986
rect 391940 158160 391992 158166
rect 391940 158102 391992 158108
rect 391848 154012 391900 154018
rect 391848 153954 391900 153960
rect 391756 153876 391808 153882
rect 391756 153818 391808 153824
rect 391572 152788 391624 152794
rect 391572 152730 391624 152736
rect 385224 150146 385276 150152
rect 385742 149940 385770 150198
rect 386374 150204 386426 150210
rect 386374 150146 386426 150152
rect 386512 150204 386564 150210
rect 386984 150198 387058 150226
rect 386512 150146 386564 150152
rect 386386 149940 386414 150146
rect 387030 149940 387058 150198
rect 387662 150204 387714 150210
rect 388272 150198 388346 150226
rect 388916 150198 388990 150226
rect 389560 150198 389634 150226
rect 390204 150198 390278 150226
rect 390848 150198 390922 150226
rect 391492 150198 391566 150226
rect 391952 150210 391980 158102
rect 392124 156800 392176 156806
rect 392124 156742 392176 156748
rect 392136 150226 392164 156742
rect 392320 152522 392348 163200
rect 393148 159934 393176 163200
rect 393136 159928 393188 159934
rect 393136 159870 393188 159876
rect 393412 159452 393464 159458
rect 393412 159394 393464 159400
rect 392308 152516 392360 152522
rect 392308 152458 392360 152464
rect 393424 150226 393452 159394
rect 393976 158098 394004 163200
rect 394700 158228 394752 158234
rect 394700 158170 394752 158176
rect 393964 158092 394016 158098
rect 393964 158034 394016 158040
rect 394056 154080 394108 154086
rect 394056 154022 394108 154028
rect 394068 150226 394096 154022
rect 394712 150226 394740 158170
rect 394896 155446 394924 163200
rect 395724 159458 395752 163200
rect 396552 161474 396580 163200
rect 396552 161446 396672 161474
rect 395712 159452 395764 159458
rect 395712 159394 395764 159400
rect 396540 156868 396592 156874
rect 396540 156810 396592 156816
rect 396172 155576 396224 155582
rect 396172 155518 396224 155524
rect 394884 155440 394936 155446
rect 394884 155382 394936 155388
rect 395344 154488 395396 154494
rect 395344 154430 395396 154436
rect 395356 150226 395384 154430
rect 395988 152720 396040 152726
rect 395988 152662 396040 152668
rect 396000 150226 396028 152662
rect 387662 150146 387714 150152
rect 387674 149940 387702 150146
rect 388318 149940 388346 150198
rect 388962 149940 388990 150198
rect 389606 149940 389634 150198
rect 390250 149940 390278 150198
rect 390894 149940 390922 150198
rect 391538 149940 391566 150198
rect 391940 150204 391992 150210
rect 392136 150198 392210 150226
rect 391940 150146 391992 150152
rect 392182 149940 392210 150198
rect 392814 150204 392866 150210
rect 393424 150198 393498 150226
rect 394068 150198 394142 150226
rect 394712 150198 394786 150226
rect 395356 150198 395430 150226
rect 396000 150198 396074 150226
rect 396184 150210 396212 155518
rect 396552 150226 396580 156810
rect 396644 152726 396672 161446
rect 397380 155378 397408 163200
rect 397368 155372 397420 155378
rect 397368 155314 397420 155320
rect 398208 154086 398236 163200
rect 398472 159520 398524 159526
rect 398472 159462 398524 159468
rect 398196 154080 398248 154086
rect 398196 154022 398248 154028
rect 396632 152720 396684 152726
rect 396632 152662 396684 152668
rect 397828 152584 397880 152590
rect 397828 152526 397880 152532
rect 397840 150226 397868 152526
rect 398484 150226 398512 159462
rect 399036 152590 399064 163200
rect 399864 159526 399892 163200
rect 400404 159792 400456 159798
rect 400404 159734 400456 159740
rect 399852 159520 399904 159526
rect 399852 159462 399904 159468
rect 399116 158296 399168 158302
rect 399116 158238 399168 158244
rect 399024 152584 399076 152590
rect 399024 152526 399076 152532
rect 399128 150226 399156 158238
rect 400220 155712 400272 155718
rect 400220 155654 400272 155660
rect 399760 154148 399812 154154
rect 399760 154090 399812 154096
rect 399772 150226 399800 154090
rect 392814 150146 392866 150152
rect 392826 149940 392854 150146
rect 393470 149940 393498 150198
rect 394114 149940 394142 150198
rect 394758 149940 394786 150198
rect 395402 149940 395430 150198
rect 396046 149940 396074 150198
rect 396172 150204 396224 150210
rect 396552 150198 396626 150226
rect 396172 150146 396224 150152
rect 396598 149940 396626 150198
rect 397230 150204 397282 150210
rect 397840 150198 397914 150226
rect 398484 150198 398558 150226
rect 399128 150198 399202 150226
rect 399772 150198 399846 150226
rect 400232 150210 400260 155654
rect 400416 150226 400444 159734
rect 400784 156874 400812 163200
rect 400772 156868 400824 156874
rect 400772 156810 400824 156816
rect 401612 156806 401640 163200
rect 402440 159798 402468 163200
rect 402428 159792 402480 159798
rect 402428 159734 402480 159740
rect 403164 159384 403216 159390
rect 403164 159326 403216 159332
rect 401600 156800 401652 156806
rect 401600 156742 401652 156748
rect 401692 155780 401744 155786
rect 401692 155722 401744 155728
rect 401704 150226 401732 155722
rect 402336 154216 402388 154222
rect 402336 154158 402388 154164
rect 402348 150226 402376 154158
rect 402980 152856 403032 152862
rect 402980 152798 403032 152804
rect 402992 150226 403020 152798
rect 403176 151814 403204 159326
rect 403268 152862 403296 163200
rect 404096 158166 404124 163200
rect 404924 158234 404952 163200
rect 405556 159860 405608 159866
rect 405556 159802 405608 159808
rect 404912 158228 404964 158234
rect 404912 158170 404964 158176
rect 404084 158160 404136 158166
rect 404084 158102 404136 158108
rect 404452 157004 404504 157010
rect 404452 156946 404504 156952
rect 404084 156936 404136 156942
rect 404084 156878 404136 156884
rect 403256 152856 403308 152862
rect 403256 152798 403308 152804
rect 404096 151814 404124 156878
rect 404464 151814 404492 156946
rect 403176 151786 403664 151814
rect 404096 151786 404308 151814
rect 404464 151786 404952 151814
rect 403636 150226 403664 151786
rect 404280 150226 404308 151786
rect 404924 150226 404952 151786
rect 405568 150226 405596 159802
rect 405752 158846 405780 163200
rect 406672 159866 406700 163200
rect 406660 159860 406712 159866
rect 406660 159802 406712 159808
rect 405740 158840 405792 158846
rect 405740 158782 405792 158788
rect 406936 158840 406988 158846
rect 406936 158782 406988 158788
rect 406844 158500 406896 158506
rect 406844 158442 406896 158448
rect 406200 152652 406252 152658
rect 406200 152594 406252 152600
rect 406212 150226 406240 152594
rect 406856 150226 406884 158442
rect 406948 152658 406976 158782
rect 407396 158364 407448 158370
rect 407396 158306 407448 158312
rect 406936 152652 406988 152658
rect 406936 152594 406988 152600
rect 407408 151814 407436 158306
rect 407500 154154 407528 163200
rect 408328 155514 408356 163200
rect 409156 160070 409184 163200
rect 409144 160064 409196 160070
rect 409144 160006 409196 160012
rect 408500 159724 408552 159730
rect 408500 159666 408552 159672
rect 408316 155508 408368 155514
rect 408316 155450 408368 155456
rect 407488 154148 407540 154154
rect 407488 154090 407540 154096
rect 408512 153202 408540 159666
rect 408776 159588 408828 159594
rect 408776 159530 408828 159536
rect 408500 153196 408552 153202
rect 408500 153138 408552 153144
rect 408132 152924 408184 152930
rect 408132 152866 408184 152872
rect 407408 151786 407528 151814
rect 407500 150226 407528 151786
rect 408144 150226 408172 152866
rect 408788 150226 408816 159530
rect 409420 153944 409472 153950
rect 409420 153886 409472 153892
rect 409432 150226 409460 153886
rect 409984 153066 410012 163200
rect 410812 155242 410840 163200
rect 411352 157072 411404 157078
rect 411352 157014 411404 157020
rect 410064 155236 410116 155242
rect 410064 155178 410116 155184
rect 410800 155236 410852 155242
rect 410800 155178 410852 155184
rect 409972 153060 410024 153066
rect 409972 153002 410024 153008
rect 410076 150226 410104 155178
rect 410708 153196 410760 153202
rect 410708 153138 410760 153144
rect 410720 150226 410748 153138
rect 411364 150226 411392 157014
rect 411640 156942 411668 163200
rect 411628 156936 411680 156942
rect 411628 156878 411680 156884
rect 411996 155304 412048 155310
rect 411996 155246 412048 155252
rect 412008 150226 412036 155246
rect 412560 152930 412588 163200
rect 412824 159996 412876 160002
rect 412824 159938 412876 159944
rect 412640 156732 412692 156738
rect 412640 156674 412692 156680
rect 412548 152924 412600 152930
rect 412548 152866 412600 152872
rect 412652 150226 412680 156674
rect 397230 150146 397282 150152
rect 397242 149940 397270 150146
rect 397886 149940 397914 150198
rect 398530 149940 398558 150198
rect 399174 149940 399202 150198
rect 399818 149940 399846 150198
rect 400220 150204 400272 150210
rect 400416 150198 400490 150226
rect 400220 150146 400272 150152
rect 400462 149940 400490 150198
rect 401094 150204 401146 150210
rect 401704 150198 401778 150226
rect 402348 150198 402422 150226
rect 402992 150198 403066 150226
rect 403636 150198 403710 150226
rect 404280 150198 404354 150226
rect 404924 150198 404998 150226
rect 405568 150198 405642 150226
rect 406212 150198 406286 150226
rect 406856 150198 406930 150226
rect 407500 150198 407574 150226
rect 408144 150198 408218 150226
rect 408788 150198 408862 150226
rect 409432 150198 409506 150226
rect 410076 150198 410150 150226
rect 410720 150198 410794 150226
rect 411364 150198 411438 150226
rect 412008 150198 412082 150226
rect 412652 150198 412726 150226
rect 412836 150210 412864 159938
rect 413388 159730 413416 163200
rect 413376 159724 413428 159730
rect 413376 159666 413428 159672
rect 414216 156670 414244 163200
rect 414296 159656 414348 159662
rect 414296 159598 414348 159604
rect 414112 156664 414164 156670
rect 414112 156606 414164 156612
rect 414204 156664 414256 156670
rect 414204 156606 414256 156612
rect 413284 152992 413336 152998
rect 413284 152934 413336 152940
rect 413296 150226 413324 152934
rect 414124 151814 414152 156606
rect 414308 152454 414336 159598
rect 415044 158030 415072 163200
rect 414572 158024 414624 158030
rect 414572 157966 414624 157972
rect 415032 158024 415084 158030
rect 415032 157966 415084 157972
rect 414296 152448 414348 152454
rect 414296 152390 414348 152396
rect 414584 151814 414612 157966
rect 415872 152998 415900 163200
rect 415860 152992 415912 152998
rect 415860 152934 415912 152940
rect 416700 152794 416728 163200
rect 417148 154012 417200 154018
rect 417148 153954 417200 153960
rect 416504 152788 416556 152794
rect 416504 152730 416556 152736
rect 416688 152788 416740 152794
rect 416688 152730 416740 152736
rect 415860 152448 415912 152454
rect 415860 152390 415912 152396
rect 414124 151786 414520 151814
rect 414584 151786 415256 151814
rect 414492 150226 414520 151786
rect 415228 150226 415256 151786
rect 415872 150226 415900 152390
rect 416516 150226 416544 152730
rect 417160 150226 417188 153954
rect 417528 153950 417556 163200
rect 418448 153950 418476 163200
rect 419080 159928 419132 159934
rect 419080 159870 419132 159876
rect 417516 153944 417568 153950
rect 417516 153886 417568 153892
rect 418436 153944 418488 153950
rect 418436 153886 418488 153892
rect 417792 153876 417844 153882
rect 417792 153818 417844 153824
rect 417804 150226 417832 153818
rect 418436 152516 418488 152522
rect 418436 152458 418488 152464
rect 418448 150226 418476 152458
rect 419092 150226 419120 159870
rect 419276 156738 419304 163200
rect 420104 159662 420132 163200
rect 420092 159656 420144 159662
rect 420092 159598 420144 159604
rect 420932 158098 420960 163200
rect 421104 159452 421156 159458
rect 421104 159394 421156 159400
rect 419540 158092 419592 158098
rect 419540 158034 419592 158040
rect 420920 158092 420972 158098
rect 420920 158034 420972 158040
rect 419264 156732 419316 156738
rect 419264 156674 419316 156680
rect 419552 151814 419580 158034
rect 420368 155440 420420 155446
rect 420368 155382 420420 155388
rect 419552 151786 419764 151814
rect 419736 150226 419764 151786
rect 420380 150226 420408 155382
rect 421116 150226 421144 159394
rect 421760 155310 421788 163200
rect 422300 155372 422352 155378
rect 422300 155314 422352 155320
rect 421748 155304 421800 155310
rect 421748 155246 421800 155252
rect 421656 152720 421708 152726
rect 421656 152662 421708 152668
rect 401094 150146 401146 150152
rect 401106 149940 401134 150146
rect 401750 149940 401778 150198
rect 402394 149940 402422 150198
rect 403038 149940 403066 150198
rect 403682 149940 403710 150198
rect 404326 149940 404354 150198
rect 404970 149940 404998 150198
rect 405614 149940 405642 150198
rect 406258 149940 406286 150198
rect 406902 149940 406930 150198
rect 407546 149940 407574 150198
rect 408190 149940 408218 150198
rect 408834 149940 408862 150198
rect 409478 149940 409506 150198
rect 410122 149940 410150 150198
rect 410766 149940 410794 150198
rect 411410 149940 411438 150198
rect 412054 149940 412082 150198
rect 412698 149940 412726 150198
rect 412824 150204 412876 150210
rect 413296 150198 413370 150226
rect 412824 150146 412876 150152
rect 413342 149940 413370 150198
rect 413974 150204 414026 150210
rect 414492 150198 414658 150226
rect 415228 150198 415302 150226
rect 415872 150198 415946 150226
rect 416516 150198 416590 150226
rect 417160 150198 417234 150226
rect 417804 150198 417878 150226
rect 418448 150198 418522 150226
rect 419092 150198 419166 150226
rect 419736 150198 419810 150226
rect 420380 150198 420454 150226
rect 413974 150146 414026 150152
rect 413986 149940 414014 150146
rect 414630 149940 414658 150198
rect 415274 149940 415302 150198
rect 415918 149940 415946 150198
rect 416562 149940 416590 150198
rect 417206 149940 417234 150198
rect 417850 149940 417878 150198
rect 418494 149940 418522 150198
rect 419138 149940 419166 150198
rect 419782 149940 419810 150198
rect 420426 149940 420454 150198
rect 421070 150198 421144 150226
rect 421668 150226 421696 152662
rect 422312 150226 422340 155314
rect 422588 154222 422616 163200
rect 423416 157010 423444 163200
rect 424232 159520 424284 159526
rect 424232 159462 424284 159468
rect 423404 157004 423456 157010
rect 423404 156946 423456 156952
rect 423772 156868 423824 156874
rect 423772 156810 423824 156816
rect 422576 154216 422628 154222
rect 422576 154158 422628 154164
rect 422944 154080 422996 154086
rect 422944 154022 422996 154028
rect 422956 150226 422984 154022
rect 423588 152584 423640 152590
rect 423588 152526 423640 152532
rect 423600 150226 423628 152526
rect 421668 150198 421742 150226
rect 422312 150198 422386 150226
rect 422956 150198 423030 150226
rect 423600 150198 423674 150226
rect 423784 150210 423812 156810
rect 424244 150226 424272 159462
rect 424336 155378 424364 163200
rect 425164 161474 425192 163200
rect 425164 161446 425284 161474
rect 425152 156800 425204 156806
rect 425152 156742 425204 156748
rect 424324 155372 424376 155378
rect 424324 155314 424376 155320
rect 425164 151814 425192 156742
rect 425256 154018 425284 161446
rect 425992 160070 426020 163200
rect 425980 160064 426032 160070
rect 425980 160006 426032 160012
rect 426440 160064 426492 160070
rect 426440 160006 426492 160012
rect 426164 159792 426216 159798
rect 426164 159734 426216 159740
rect 425244 154012 425296 154018
rect 425244 153954 425296 153960
rect 425164 151786 425560 151814
rect 425532 150226 425560 151786
rect 426176 150226 426204 159734
rect 426452 158302 426480 160006
rect 426820 159118 426848 163200
rect 426808 159112 426860 159118
rect 426808 159054 426860 159060
rect 426440 158296 426492 158302
rect 426440 158238 426492 158244
rect 427360 158160 427412 158166
rect 427360 158102 427412 158108
rect 426808 152856 426860 152862
rect 426808 152798 426860 152804
rect 426820 150226 426848 152798
rect 427372 150226 427400 158102
rect 427648 156806 427676 163200
rect 428004 158228 428056 158234
rect 428004 158170 428056 158176
rect 427636 156800 427688 156806
rect 427636 156742 427688 156748
rect 428016 150226 428044 158170
rect 428476 158166 428504 163200
rect 428464 158160 428516 158166
rect 428464 158102 428516 158108
rect 429304 155446 429332 163200
rect 429384 159860 429436 159866
rect 429384 159802 429436 159808
rect 429292 155440 429344 155446
rect 429292 155382 429344 155388
rect 428648 152652 428700 152658
rect 428648 152594 428700 152600
rect 428660 150226 428688 152594
rect 429396 150226 429424 159802
rect 430224 158778 430252 163200
rect 430212 158772 430264 158778
rect 430212 158714 430264 158720
rect 430580 155508 430632 155514
rect 430580 155450 430632 155456
rect 429936 154148 429988 154154
rect 429936 154090 429988 154096
rect 421070 149940 421098 150198
rect 421714 149940 421742 150198
rect 422358 149940 422386 150198
rect 423002 149940 423030 150198
rect 423646 149940 423674 150198
rect 423772 150204 423824 150210
rect 424244 150198 424318 150226
rect 423772 150146 423824 150152
rect 424290 149940 424318 150198
rect 424922 150204 424974 150210
rect 425532 150198 425606 150226
rect 426176 150198 426250 150226
rect 426820 150198 426894 150226
rect 427372 150198 427446 150226
rect 428016 150198 428090 150226
rect 428660 150198 428734 150226
rect 424922 150146 424974 150152
rect 424934 149940 424962 150146
rect 425578 149940 425606 150198
rect 426222 149940 426250 150198
rect 426866 149940 426894 150198
rect 427418 149940 427446 150198
rect 428062 149940 428090 150198
rect 428706 149940 428734 150198
rect 429350 150198 429424 150226
rect 429948 150226 429976 154090
rect 430592 150226 430620 155450
rect 431052 154154 431080 163200
rect 431224 159996 431276 160002
rect 431224 159938 431276 159944
rect 431040 154148 431092 154154
rect 431040 154090 431092 154096
rect 431236 150226 431264 159938
rect 431880 159594 431908 163200
rect 431868 159588 431920 159594
rect 431868 159530 431920 159536
rect 432708 159458 432736 163200
rect 433536 159526 433564 163200
rect 433524 159520 433576 159526
rect 433524 159462 433576 159468
rect 432696 159452 432748 159458
rect 432696 159394 432748 159400
rect 434364 159390 434392 163200
rect 434444 159724 434496 159730
rect 434444 159666 434496 159672
rect 434352 159384 434404 159390
rect 434352 159326 434404 159332
rect 433064 159112 433116 159118
rect 433064 159054 433116 159060
rect 433076 155514 433104 159054
rect 433248 158772 433300 158778
rect 433248 158714 433300 158720
rect 433156 156936 433208 156942
rect 433156 156878 433208 156884
rect 433064 155508 433116 155514
rect 433064 155450 433116 155456
rect 432052 155236 432104 155242
rect 432052 155178 432104 155184
rect 431868 153060 431920 153066
rect 431868 153002 431920 153008
rect 431880 150226 431908 153002
rect 432064 151814 432092 155178
rect 432064 151786 432552 151814
rect 432524 150226 432552 151786
rect 433168 150226 433196 156878
rect 433260 156874 433288 158714
rect 433248 156868 433300 156874
rect 433248 156810 433300 156816
rect 433800 152924 433852 152930
rect 433800 152866 433852 152872
rect 433812 150226 433840 152866
rect 434456 150226 434484 159666
rect 435192 158030 435220 163200
rect 435824 159656 435876 159662
rect 435824 159598 435876 159604
rect 434720 158024 434772 158030
rect 434720 157966 434772 157972
rect 435180 158024 435232 158030
rect 435180 157966 435232 157972
rect 429948 150198 430022 150226
rect 430592 150198 430666 150226
rect 431236 150198 431310 150226
rect 431880 150198 431954 150226
rect 432524 150198 432598 150226
rect 433168 150198 433242 150226
rect 433812 150198 433886 150226
rect 434456 150198 434530 150226
rect 434732 150210 434760 157966
rect 435088 156664 435140 156670
rect 435088 156606 435140 156612
rect 435100 150226 435128 156606
rect 435836 153202 435864 159598
rect 436112 158846 436140 163200
rect 436940 163146 436968 163200
rect 437032 163146 437060 163254
rect 436940 163118 437060 163146
rect 436560 159588 436612 159594
rect 436560 159530 436612 159536
rect 436100 158840 436152 158846
rect 436100 158782 436152 158788
rect 436572 156942 436600 159530
rect 436560 156936 436612 156942
rect 436560 156878 436612 156884
rect 435824 153196 435876 153202
rect 435824 153138 435876 153144
rect 436376 152992 436428 152998
rect 436376 152934 436428 152940
rect 436388 150226 436416 152934
rect 437020 152788 437072 152794
rect 437020 152730 437072 152736
rect 437032 150226 437060 152730
rect 437400 152522 437428 163254
rect 437754 163200 437810 164400
rect 438582 163200 438638 164400
rect 439410 163200 439466 164400
rect 440238 163200 440294 164400
rect 441066 163200 441122 164400
rect 441986 163200 442042 164400
rect 442814 163200 442870 164400
rect 443642 163200 443698 164400
rect 444470 163200 444526 164400
rect 445298 163200 445354 164400
rect 446126 163200 446182 164400
rect 446954 163200 447010 164400
rect 447874 163200 447930 164400
rect 448702 163200 448758 164400
rect 449530 163200 449586 164400
rect 450358 163200 450414 164400
rect 451186 163200 451242 164400
rect 452014 163200 452070 164400
rect 452842 163200 452898 164400
rect 453762 163200 453818 164400
rect 454590 163200 454646 164400
rect 455418 163200 455474 164400
rect 456246 163200 456302 164400
rect 457074 163200 457130 164400
rect 457902 163200 457958 164400
rect 458730 163200 458786 164400
rect 459650 163200 459706 164400
rect 460478 163200 460534 164400
rect 460584 163254 460888 163282
rect 437768 158982 437796 163200
rect 437756 158976 437808 158982
rect 437756 158918 437808 158924
rect 438308 153944 438360 153950
rect 438308 153886 438360 153892
rect 437664 153876 437716 153882
rect 437664 153818 437716 153824
rect 437388 152516 437440 152522
rect 437388 152458 437440 152464
rect 437676 150226 437704 153818
rect 438320 150226 438348 153886
rect 438596 153814 438624 163200
rect 438860 158840 438912 158846
rect 438860 158782 438912 158788
rect 438872 154222 438900 158782
rect 439424 158234 439452 163200
rect 439412 158228 439464 158234
rect 439412 158170 439464 158176
rect 438952 156732 439004 156738
rect 438952 156674 439004 156680
rect 438860 154216 438912 154222
rect 438860 154158 438912 154164
rect 438584 153808 438636 153814
rect 438584 153750 438636 153756
rect 438964 150226 438992 156674
rect 440252 153950 440280 163200
rect 441080 159662 441108 163200
rect 441068 159656 441120 159662
rect 441068 159598 441120 159604
rect 440332 158092 440384 158098
rect 440332 158034 440384 158040
rect 440240 153944 440292 153950
rect 440240 153886 440292 153892
rect 439596 153196 439648 153202
rect 439596 153138 439648 153144
rect 439608 150226 439636 153138
rect 440344 150226 440372 158034
rect 441712 155372 441764 155378
rect 441712 155314 441764 155320
rect 440884 155304 440936 155310
rect 440884 155246 440936 155252
rect 429350 149940 429378 150198
rect 429994 149940 430022 150198
rect 430638 149940 430666 150198
rect 431282 149940 431310 150198
rect 431926 149940 431954 150198
rect 432570 149940 432598 150198
rect 433214 149940 433242 150198
rect 433858 149940 433886 150198
rect 434502 149940 434530 150198
rect 434720 150204 434772 150210
rect 435100 150198 435174 150226
rect 434720 150146 434772 150152
rect 435146 149940 435174 150198
rect 435778 150204 435830 150210
rect 436388 150198 436462 150226
rect 437032 150198 437106 150226
rect 437676 150198 437750 150226
rect 438320 150198 438394 150226
rect 438964 150198 439038 150226
rect 439608 150198 439682 150226
rect 435778 150146 435830 150152
rect 435790 149940 435818 150146
rect 436434 149940 436462 150198
rect 437078 149940 437106 150198
rect 437722 149940 437750 150198
rect 438366 149940 438394 150198
rect 439010 149940 439038 150198
rect 439654 149940 439682 150198
rect 440298 150198 440372 150226
rect 440896 150226 440924 155246
rect 441436 154080 441488 154086
rect 441436 154022 441488 154028
rect 441448 151814 441476 154022
rect 441448 151786 441568 151814
rect 441540 150226 441568 151786
rect 440896 150198 440970 150226
rect 441540 150198 441614 150226
rect 441724 150210 441752 155314
rect 442000 155310 442028 163200
rect 442172 157004 442224 157010
rect 442172 156946 442224 156952
rect 441988 155304 442040 155310
rect 441988 155246 442040 155252
rect 442184 150226 442212 156946
rect 442828 155242 442856 163200
rect 443000 158296 443052 158302
rect 443000 158238 443052 158244
rect 442816 155236 442868 155242
rect 442816 155178 442868 155184
rect 440298 149940 440326 150198
rect 440942 149940 440970 150198
rect 441586 149940 441614 150198
rect 441712 150204 441764 150210
rect 442184 150198 442258 150226
rect 443012 150210 443040 158238
rect 443656 158098 443684 163200
rect 444288 158976 444340 158982
rect 444288 158918 444340 158924
rect 443644 158092 443696 158098
rect 443644 158034 443696 158040
rect 443460 154012 443512 154018
rect 443460 153954 443512 153960
rect 443472 150226 443500 153954
rect 444300 152794 444328 158918
rect 444380 156800 444432 156806
rect 444380 156742 444432 156748
rect 444288 152788 444340 152794
rect 444288 152730 444340 152736
rect 441712 150146 441764 150152
rect 442230 149940 442258 150198
rect 442862 150204 442914 150210
rect 442862 150146 442914 150152
rect 443000 150204 443052 150210
rect 443472 150198 443546 150226
rect 444392 150210 444420 156742
rect 444484 155378 444512 163200
rect 445312 156670 445340 163200
rect 445484 159656 445536 159662
rect 445484 159598 445536 159604
rect 445300 156664 445352 156670
rect 445300 156606 445352 156612
rect 444748 155508 444800 155514
rect 444748 155450 444800 155456
rect 444472 155372 444524 155378
rect 444472 155314 444524 155320
rect 444760 150226 444788 155450
rect 445496 152726 445524 159598
rect 445760 158160 445812 158166
rect 445760 158102 445812 158108
rect 445484 152720 445536 152726
rect 445484 152662 445536 152668
rect 445772 151814 445800 158102
rect 446140 156738 446168 163200
rect 446128 156732 446180 156738
rect 446128 156674 446180 156680
rect 446680 155440 446732 155446
rect 446680 155382 446732 155388
rect 445772 151786 446076 151814
rect 446048 150226 446076 151786
rect 446692 150226 446720 155382
rect 446968 152590 446996 163200
rect 447140 159452 447192 159458
rect 447140 159394 447192 159400
rect 447152 153202 447180 159394
rect 447888 158982 447916 163200
rect 447876 158976 447928 158982
rect 447876 158918 447928 158924
rect 448716 158166 448744 163200
rect 449544 158846 449572 163200
rect 449808 159520 449860 159526
rect 449808 159462 449860 159468
rect 449532 158840 449584 158846
rect 449532 158782 449584 158788
rect 448704 158160 448756 158166
rect 448704 158102 448756 158108
rect 448612 156936 448664 156942
rect 448612 156878 448664 156884
rect 447324 156868 447376 156874
rect 447324 156810 447376 156816
rect 447140 153196 447192 153202
rect 447140 153138 447192 153144
rect 446956 152584 447008 152590
rect 446956 152526 447008 152532
rect 447336 150226 447364 156810
rect 447968 154148 448020 154154
rect 447968 154090 448020 154096
rect 447980 150226 448008 154090
rect 448624 150226 448652 156878
rect 449256 153196 449308 153202
rect 449256 153138 449308 153144
rect 449268 150226 449296 153138
rect 449820 151814 449848 159462
rect 450084 159384 450136 159390
rect 450084 159326 450136 159332
rect 450096 151814 450124 159326
rect 450372 152658 450400 163200
rect 451200 159526 451228 163200
rect 451188 159520 451240 159526
rect 451188 159462 451240 159468
rect 451096 158024 451148 158030
rect 451096 157966 451148 157972
rect 450360 152652 450412 152658
rect 450360 152594 450412 152600
rect 451108 151814 451136 157966
rect 451832 154216 451884 154222
rect 451832 154158 451884 154164
rect 449820 151786 449940 151814
rect 450096 151786 450584 151814
rect 451108 151786 451228 151814
rect 449912 150226 449940 151786
rect 450556 150226 450584 151786
rect 451200 150226 451228 151786
rect 451844 150226 451872 154158
rect 452028 152454 452056 163200
rect 452476 158976 452528 158982
rect 452476 158918 452528 158924
rect 452488 153202 452516 158918
rect 452476 153196 452528 153202
rect 452476 153138 452528 153144
rect 452856 152930 452884 163200
rect 453776 159050 453804 163200
rect 453764 159044 453816 159050
rect 453764 158986 453816 158992
rect 453948 158840 454000 158846
rect 453948 158782 454000 158788
rect 453960 153882 453988 158782
rect 454408 158228 454460 158234
rect 454408 158170 454460 158176
rect 453948 153876 454000 153882
rect 453948 153818 454000 153824
rect 453764 153808 453816 153814
rect 453764 153750 453816 153756
rect 452844 152924 452896 152930
rect 452844 152866 452896 152872
rect 453120 152788 453172 152794
rect 453120 152730 453172 152736
rect 452476 152516 452528 152522
rect 452476 152458 452528 152464
rect 452016 152448 452068 152454
rect 452016 152390 452068 152396
rect 452488 150226 452516 152458
rect 453132 150226 453160 152730
rect 453776 150226 453804 153750
rect 454420 150226 454448 158170
rect 454604 152998 454632 163200
rect 455328 159520 455380 159526
rect 455328 159462 455380 159468
rect 455052 153944 455104 153950
rect 455052 153886 455104 153892
rect 454592 152992 454644 152998
rect 454592 152934 454644 152940
rect 455064 150226 455092 153886
rect 455340 153270 455368 159462
rect 455328 153264 455380 153270
rect 455328 153206 455380 153212
rect 455432 152794 455460 163200
rect 456260 155310 456288 163200
rect 456800 158092 456852 158098
rect 456800 158034 456852 158040
rect 456248 155304 456300 155310
rect 456248 155246 456300 155252
rect 456340 155236 456392 155242
rect 456340 155178 456392 155184
rect 455420 152788 455472 152794
rect 455420 152730 455472 152736
rect 455696 152720 455748 152726
rect 455696 152662 455748 152668
rect 455708 150226 455736 152662
rect 456352 150226 456380 155178
rect 443000 150146 443052 150152
rect 442874 149940 442902 150146
rect 443518 149940 443546 150198
rect 444150 150204 444202 150210
rect 444150 150146 444202 150152
rect 444380 150204 444432 150210
rect 444760 150198 444834 150226
rect 444380 150146 444432 150152
rect 444162 149940 444190 150146
rect 444806 149940 444834 150198
rect 445438 150204 445490 150210
rect 446048 150198 446122 150226
rect 446692 150198 446766 150226
rect 447336 150198 447410 150226
rect 447980 150198 448054 150226
rect 448624 150198 448698 150226
rect 449268 150198 449342 150226
rect 449912 150198 449986 150226
rect 450556 150198 450630 150226
rect 451200 150198 451274 150226
rect 451844 150198 451918 150226
rect 452488 150198 452562 150226
rect 453132 150198 453206 150226
rect 453776 150198 453850 150226
rect 454420 150198 454494 150226
rect 455064 150198 455138 150226
rect 455708 150198 455782 150226
rect 456352 150198 456426 150226
rect 456812 150210 456840 158034
rect 456984 155168 457036 155174
rect 456984 155110 457036 155116
rect 456996 150226 457024 155110
rect 457088 152930 457116 163200
rect 457916 158030 457944 163200
rect 458180 159044 458232 159050
rect 458180 158986 458232 158992
rect 457904 158024 457956 158030
rect 457904 157966 457956 157972
rect 458192 156670 458220 158986
rect 458744 158778 458772 163200
rect 458732 158772 458784 158778
rect 458732 158714 458784 158720
rect 459468 156732 459520 156738
rect 459468 156674 459520 156680
rect 458180 156664 458232 156670
rect 458180 156606 458232 156612
rect 458364 156596 458416 156602
rect 458364 156538 458416 156544
rect 458180 155372 458232 155378
rect 458180 155314 458232 155320
rect 457076 152924 457128 152930
rect 457076 152866 457128 152872
rect 458192 150226 458220 155314
rect 458376 151814 458404 156538
rect 458376 151786 458864 151814
rect 458836 150226 458864 151786
rect 459480 150226 459508 156674
rect 459664 152522 459692 163200
rect 460492 163146 460520 163200
rect 460584 163146 460612 163254
rect 460492 163118 460612 163146
rect 460664 153196 460716 153202
rect 460664 153138 460716 153144
rect 460112 152584 460164 152590
rect 460112 152526 460164 152532
rect 459652 152516 459704 152522
rect 459652 152458 459704 152464
rect 460124 150226 460152 152526
rect 460676 151814 460704 153138
rect 460860 152998 460888 163254
rect 461306 163200 461362 164400
rect 462134 163200 462190 164400
rect 462962 163200 463018 164400
rect 463790 163200 463846 164400
rect 464618 163200 464674 164400
rect 464724 163254 465028 163282
rect 461320 159390 461348 163200
rect 461308 159384 461360 159390
rect 461308 159326 461360 159332
rect 461400 158160 461452 158166
rect 461400 158102 461452 158108
rect 460848 152992 460900 152998
rect 460848 152934 460900 152940
rect 460676 151786 460796 151814
rect 460768 150226 460796 151786
rect 461412 150226 461440 158102
rect 462044 153876 462096 153882
rect 462044 153818 462096 153824
rect 462056 150226 462084 153818
rect 462148 153066 462176 163200
rect 462136 153060 462188 153066
rect 462136 153002 462188 153008
rect 462976 152658 463004 163200
rect 463804 158982 463832 163200
rect 464632 163146 464660 163200
rect 464724 163146 464752 163254
rect 464632 163118 464752 163146
rect 464896 159384 464948 159390
rect 464896 159326 464948 159332
rect 463792 158976 463844 158982
rect 463792 158918 463844 158924
rect 463332 158772 463384 158778
rect 463332 158714 463384 158720
rect 463344 154562 463372 158714
rect 464908 157010 464936 159326
rect 464896 157004 464948 157010
rect 464896 156946 464948 156952
rect 463332 154556 463384 154562
rect 463332 154498 463384 154504
rect 463332 153264 463384 153270
rect 463332 153206 463384 153212
rect 462688 152652 462740 152658
rect 462688 152594 462740 152600
rect 462964 152652 463016 152658
rect 462964 152594 463016 152600
rect 462700 150226 462728 152594
rect 463344 150226 463372 153206
rect 464620 152788 464672 152794
rect 464620 152730 464672 152736
rect 463976 152516 464028 152522
rect 463976 152458 464028 152464
rect 463988 150226 464016 152458
rect 464632 150226 464660 152730
rect 465000 152522 465028 163254
rect 465538 163200 465594 164400
rect 466366 163200 466422 164400
rect 467194 163200 467250 164400
rect 468022 163200 468078 164400
rect 468850 163200 468906 164400
rect 468956 163254 469168 163282
rect 465264 156664 465316 156670
rect 465264 156606 465316 156612
rect 464988 152516 465040 152522
rect 464988 152458 465040 152464
rect 465276 150226 465304 156606
rect 465552 153134 465580 163200
rect 466380 158098 466408 163200
rect 466368 158092 466420 158098
rect 466368 158034 466420 158040
rect 467104 155304 467156 155310
rect 467104 155246 467156 155252
rect 465540 153128 465592 153134
rect 465540 153070 465592 153076
rect 465908 152856 465960 152862
rect 465908 152798 465960 152804
rect 465920 150226 465948 152798
rect 466552 152720 466604 152726
rect 466552 152662 466604 152668
rect 466564 150226 466592 152662
rect 467116 151814 467144 155246
rect 467208 152794 467236 163200
rect 467840 152924 467892 152930
rect 467840 152866 467892 152872
rect 467196 152788 467248 152794
rect 467196 152730 467248 152736
rect 467116 151786 467236 151814
rect 467208 150226 467236 151786
rect 467852 150226 467880 152866
rect 468036 152726 468064 163200
rect 468864 163146 468892 163200
rect 468956 163146 468984 163254
rect 468864 163118 468984 163146
rect 468484 158024 468536 158030
rect 468484 157966 468536 157972
rect 468024 152720 468076 152726
rect 468024 152662 468076 152668
rect 468496 150226 468524 157966
rect 468944 154556 468996 154562
rect 468944 154498 468996 154504
rect 468956 151814 468984 154498
rect 469140 152930 469168 163254
rect 469678 163200 469734 164400
rect 470506 163200 470562 164400
rect 471426 163200 471482 164400
rect 472254 163200 472310 164400
rect 473082 163200 473138 164400
rect 473910 163200 473966 164400
rect 474738 163200 474794 164400
rect 475566 163200 475622 164400
rect 476394 163200 476450 164400
rect 477314 163200 477370 164400
rect 478142 163200 478198 164400
rect 478970 163200 479026 164400
rect 479798 163200 479854 164400
rect 480626 163200 480682 164400
rect 481454 163200 481510 164400
rect 482282 163200 482338 164400
rect 483202 163200 483258 164400
rect 484030 163200 484086 164400
rect 484858 163200 484914 164400
rect 485686 163200 485742 164400
rect 486514 163200 486570 164400
rect 487342 163200 487398 164400
rect 488170 163200 488226 164400
rect 489090 163200 489146 164400
rect 489918 163200 489974 164400
rect 490746 163200 490802 164400
rect 491574 163200 491630 164400
rect 492402 163200 492458 164400
rect 493230 163200 493286 164400
rect 494058 163200 494114 164400
rect 494978 163200 495034 164400
rect 495806 163200 495862 164400
rect 496634 163200 496690 164400
rect 497462 163200 497518 164400
rect 498290 163200 498346 164400
rect 499118 163200 499174 164400
rect 499224 163254 499528 163282
rect 469128 152924 469180 152930
rect 469128 152866 469180 152872
rect 469692 152862 469720 163200
rect 470324 152992 470376 152998
rect 470324 152934 470376 152940
rect 469680 152856 469732 152862
rect 469680 152798 469732 152804
rect 469772 152584 469824 152590
rect 469772 152526 469824 152532
rect 468956 151786 469168 151814
rect 469140 150226 469168 151786
rect 469784 150226 469812 152526
rect 470336 151814 470364 152934
rect 470520 152590 470548 163200
rect 471440 159118 471468 163200
rect 472268 159866 472296 163200
rect 472256 159860 472308 159866
rect 472256 159802 472308 159808
rect 471428 159112 471480 159118
rect 471428 159054 471480 159060
rect 473096 159050 473124 163200
rect 473084 159044 473136 159050
rect 473084 158986 473136 158992
rect 471796 158976 471848 158982
rect 471796 158918 471848 158924
rect 471060 157004 471112 157010
rect 471060 156946 471112 156952
rect 470508 152584 470560 152590
rect 470508 152526 470560 152532
rect 470336 151786 470456 151814
rect 470428 150226 470456 151786
rect 471072 150226 471100 156946
rect 471808 154562 471836 158918
rect 473924 158914 473952 163200
rect 473912 158908 473964 158914
rect 473912 158850 473964 158856
rect 474752 158846 474780 163200
rect 475580 158982 475608 163200
rect 475568 158976 475620 158982
rect 475568 158918 475620 158924
rect 474740 158840 474792 158846
rect 474740 158782 474792 158788
rect 476408 158778 476436 163200
rect 477328 159390 477356 163200
rect 478156 159662 478184 163200
rect 478984 159730 479012 163200
rect 479432 159860 479484 159866
rect 479432 159802 479484 159808
rect 478972 159724 479024 159730
rect 478972 159666 479024 159672
rect 478144 159656 478196 159662
rect 478144 159598 478196 159604
rect 477316 159384 477368 159390
rect 477316 159326 477368 159332
rect 477684 159112 477736 159118
rect 477684 159054 477736 159060
rect 476396 158772 476448 158778
rect 476396 158714 476448 158720
rect 474924 158092 474976 158098
rect 474924 158034 474976 158040
rect 471796 154556 471848 154562
rect 471796 154498 471848 154504
rect 472992 154556 473044 154562
rect 472992 154498 473044 154504
rect 471704 153060 471756 153066
rect 471704 153002 471756 153008
rect 471716 150226 471744 153002
rect 472348 152652 472400 152658
rect 472348 152594 472400 152600
rect 472360 150226 472388 152594
rect 473004 150226 473032 154498
rect 474280 153128 474332 153134
rect 474280 153070 474332 153076
rect 473636 152516 473688 152522
rect 473636 152458 473688 152464
rect 473648 150226 473676 152458
rect 474292 150226 474320 153070
rect 474936 150226 474964 158034
rect 476856 152924 476908 152930
rect 476856 152866 476908 152872
rect 475568 152788 475620 152794
rect 475568 152730 475620 152736
rect 475580 150226 475608 152730
rect 476212 152720 476264 152726
rect 476212 152662 476264 152668
rect 476224 150226 476252 152662
rect 476868 150226 476896 152866
rect 477500 152856 477552 152862
rect 477500 152798 477552 152804
rect 477512 150226 477540 152798
rect 445438 150146 445490 150152
rect 445450 149940 445478 150146
rect 446094 149940 446122 150198
rect 446738 149940 446766 150198
rect 447382 149940 447410 150198
rect 448026 149940 448054 150198
rect 448670 149940 448698 150198
rect 449314 149940 449342 150198
rect 449958 149940 449986 150198
rect 450602 149940 450630 150198
rect 451246 149940 451274 150198
rect 451890 149940 451918 150198
rect 452534 149940 452562 150198
rect 453178 149940 453206 150198
rect 453822 149940 453850 150198
rect 454466 149940 454494 150198
rect 455110 149940 455138 150198
rect 455754 149940 455782 150198
rect 456398 149940 456426 150198
rect 456800 150204 456852 150210
rect 456996 150198 457070 150226
rect 456800 150146 456852 150152
rect 457042 149940 457070 150198
rect 457674 150204 457726 150210
rect 458192 150198 458266 150226
rect 458836 150198 458910 150226
rect 459480 150198 459554 150226
rect 460124 150198 460198 150226
rect 460768 150198 460842 150226
rect 461412 150198 461486 150226
rect 462056 150198 462130 150226
rect 462700 150198 462774 150226
rect 463344 150198 463418 150226
rect 463988 150198 464062 150226
rect 464632 150198 464706 150226
rect 465276 150198 465350 150226
rect 465920 150198 465994 150226
rect 466564 150198 466638 150226
rect 467208 150198 467282 150226
rect 467852 150198 467926 150226
rect 468496 150198 468570 150226
rect 469140 150198 469214 150226
rect 469784 150198 469858 150226
rect 470428 150198 470502 150226
rect 471072 150198 471146 150226
rect 471716 150198 471790 150226
rect 472360 150198 472434 150226
rect 473004 150198 473078 150226
rect 473648 150198 473722 150226
rect 474292 150198 474366 150226
rect 474936 150198 475010 150226
rect 475580 150198 475654 150226
rect 476224 150198 476298 150226
rect 476868 150198 476942 150226
rect 477512 150198 477586 150226
rect 477696 150210 477724 159054
rect 478972 159044 479024 159050
rect 478972 158986 479024 158992
rect 478144 152584 478196 152590
rect 478144 152526 478196 152532
rect 478156 150226 478184 152526
rect 457674 150146 457726 150152
rect 457686 149940 457714 150146
rect 458238 149940 458266 150198
rect 458882 149940 458910 150198
rect 459526 149940 459554 150198
rect 460170 149940 460198 150198
rect 460814 149940 460842 150198
rect 461458 149940 461486 150198
rect 462102 149940 462130 150198
rect 462746 149940 462774 150198
rect 463390 149940 463418 150198
rect 464034 149940 464062 150198
rect 464678 149940 464706 150198
rect 465322 149940 465350 150198
rect 465966 149940 465994 150198
rect 466610 149940 466638 150198
rect 467254 149940 467282 150198
rect 467898 149940 467926 150198
rect 468542 149940 468570 150198
rect 469186 149940 469214 150198
rect 469830 149940 469858 150198
rect 470474 149940 470502 150198
rect 471118 149940 471146 150198
rect 471762 149940 471790 150198
rect 472406 149940 472434 150198
rect 473050 149940 473078 150198
rect 473694 149940 473722 150198
rect 474338 149940 474366 150198
rect 474982 149940 475010 150198
rect 475626 149940 475654 150198
rect 476270 149940 476298 150198
rect 476914 149940 476942 150198
rect 477558 149940 477586 150198
rect 477684 150204 477736 150210
rect 478156 150198 478230 150226
rect 478984 150210 479012 158986
rect 479444 150226 479472 159802
rect 479812 159458 479840 163200
rect 479800 159452 479852 159458
rect 479800 159394 479852 159400
rect 480640 159322 480668 163200
rect 481468 159798 481496 163200
rect 481456 159792 481508 159798
rect 481456 159734 481508 159740
rect 480628 159316 480680 159322
rect 480628 159258 480680 159264
rect 481640 158976 481692 158982
rect 481640 158918 481692 158924
rect 480260 158908 480312 158914
rect 480260 158850 480312 158856
rect 480272 151814 480300 158850
rect 481364 158840 481416 158846
rect 481364 158782 481416 158788
rect 480272 151786 480760 151814
rect 480732 150226 480760 151786
rect 481376 150226 481404 158782
rect 481652 151814 481680 158918
rect 482296 158914 482324 163200
rect 483020 159656 483072 159662
rect 483020 159598 483072 159604
rect 482284 158908 482336 158914
rect 482284 158850 482336 158856
rect 482652 158772 482704 158778
rect 482652 158714 482704 158720
rect 481652 151786 482048 151814
rect 482020 150226 482048 151786
rect 482664 150226 482692 158714
rect 477684 150146 477736 150152
rect 478202 149940 478230 150198
rect 478834 150204 478886 150210
rect 478834 150146 478886 150152
rect 478972 150204 479024 150210
rect 479444 150198 479518 150226
rect 478972 150146 479024 150152
rect 478846 149940 478874 150146
rect 479490 149940 479518 150198
rect 480122 150204 480174 150210
rect 480732 150198 480806 150226
rect 481376 150198 481450 150226
rect 482020 150198 482094 150226
rect 482664 150198 482738 150226
rect 483032 150210 483060 159598
rect 483216 158846 483244 163200
rect 483296 159384 483348 159390
rect 483296 159326 483348 159332
rect 483204 158840 483256 158846
rect 483204 158782 483256 158788
rect 483308 150226 483336 159326
rect 484044 159118 484072 163200
rect 484872 160002 484900 163200
rect 484860 159996 484912 160002
rect 484860 159938 484912 159944
rect 484400 159724 484452 159730
rect 484400 159666 484452 159672
rect 484032 159112 484084 159118
rect 484032 159054 484084 159060
rect 484412 151814 484440 159666
rect 485228 159452 485280 159458
rect 485228 159394 485280 159400
rect 484412 151786 484624 151814
rect 484596 150226 484624 151786
rect 485240 150226 485268 159394
rect 485700 158778 485728 163200
rect 485780 159792 485832 159798
rect 485780 159734 485832 159740
rect 485688 158772 485740 158778
rect 485688 158714 485740 158720
rect 480122 150146 480174 150152
rect 480134 149940 480162 150146
rect 480778 149940 480806 150198
rect 481422 149940 481450 150198
rect 482066 149940 482094 150198
rect 482710 149940 482738 150198
rect 483020 150204 483072 150210
rect 483308 150198 483382 150226
rect 483020 150146 483072 150152
rect 483354 149940 483382 150198
rect 483986 150204 484038 150210
rect 484596 150198 484670 150226
rect 485240 150198 485314 150226
rect 485792 150210 485820 159734
rect 485872 159316 485924 159322
rect 485872 159258 485924 159264
rect 485884 150226 485912 159258
rect 486528 159050 486556 163200
rect 486516 159044 486568 159050
rect 486516 158986 486568 158992
rect 487356 158982 487384 163200
rect 487344 158976 487396 158982
rect 487344 158918 487396 158924
rect 487160 158908 487212 158914
rect 487160 158850 487212 158856
rect 487172 150226 487200 158850
rect 488184 158846 488212 163200
rect 489000 159996 489052 160002
rect 489000 159938 489052 159944
rect 488448 159112 488500 159118
rect 488448 159054 488500 159060
rect 487528 158840 487580 158846
rect 487528 158782 487580 158788
rect 488172 158840 488224 158846
rect 488172 158782 488224 158788
rect 487540 151814 487568 158782
rect 487540 151786 487844 151814
rect 487816 150226 487844 151786
rect 488460 150226 488488 159054
rect 488632 158772 488684 158778
rect 488632 158714 488684 158720
rect 483986 150146 484038 150152
rect 483998 149940 484026 150146
rect 484642 149940 484670 150198
rect 485286 149940 485314 150198
rect 485780 150204 485832 150210
rect 485884 150198 485958 150226
rect 485780 150146 485832 150152
rect 485930 149940 485958 150198
rect 486562 150204 486614 150210
rect 487172 150198 487246 150226
rect 487816 150198 487890 150226
rect 488460 150198 488534 150226
rect 488644 150210 488672 158714
rect 489012 150226 489040 159938
rect 489104 158914 489132 163200
rect 489932 159254 489960 163200
rect 489920 159248 489972 159254
rect 489920 159190 489972 159196
rect 490288 159044 490340 159050
rect 490288 158986 490340 158992
rect 489920 158976 489972 158982
rect 489920 158918 489972 158924
rect 489092 158908 489144 158914
rect 489092 158850 489144 158856
rect 486562 150146 486614 150152
rect 486574 149940 486602 150146
rect 487218 149940 487246 150198
rect 487862 149940 487890 150198
rect 488506 149940 488534 150198
rect 488632 150204 488684 150210
rect 489012 150198 489086 150226
rect 489932 150210 489960 158918
rect 490300 150226 490328 158986
rect 490760 158778 490788 163200
rect 491588 158982 491616 163200
rect 492416 159798 492444 163200
rect 492404 159792 492456 159798
rect 492404 159734 492456 159740
rect 492680 159248 492732 159254
rect 492680 159190 492732 159196
rect 491576 158976 491628 158982
rect 491576 158918 491628 158924
rect 491300 158908 491352 158914
rect 491300 158850 491352 158856
rect 490748 158772 490800 158778
rect 490748 158714 490800 158720
rect 488632 150146 488684 150152
rect 489058 149940 489086 150198
rect 489690 150204 489742 150210
rect 489690 150146 489742 150152
rect 489920 150204 489972 150210
rect 490300 150198 490374 150226
rect 491312 150210 491340 158850
rect 491576 158840 491628 158846
rect 491576 158782 491628 158788
rect 491588 150226 491616 158782
rect 492692 151814 492720 159190
rect 493244 159186 493272 163200
rect 493232 159180 493284 159186
rect 493232 159122 493284 159128
rect 494072 158778 494100 163200
rect 494796 159792 494848 159798
rect 494796 159734 494848 159740
rect 494152 158976 494204 158982
rect 494152 158918 494204 158924
rect 493508 158772 493560 158778
rect 493508 158714 493560 158720
rect 494060 158772 494112 158778
rect 494060 158714 494112 158720
rect 492692 151786 492904 151814
rect 492876 150226 492904 151786
rect 493520 150226 493548 158714
rect 494164 150226 494192 158918
rect 494808 150226 494836 159734
rect 494992 159322 495020 163200
rect 494980 159316 495032 159322
rect 494980 159258 495032 159264
rect 495440 159180 495492 159186
rect 495440 159122 495492 159128
rect 495452 150226 495480 159122
rect 495820 158778 495848 163200
rect 496648 159458 496676 163200
rect 496636 159452 496688 159458
rect 496636 159394 496688 159400
rect 497476 159390 497504 163200
rect 498016 159452 498068 159458
rect 498016 159394 498068 159400
rect 497464 159384 497516 159390
rect 497464 159326 497516 159332
rect 496728 159316 496780 159322
rect 496728 159258 496780 159264
rect 495716 158772 495768 158778
rect 495716 158714 495768 158720
rect 495808 158772 495860 158778
rect 495808 158714 495860 158720
rect 495728 151814 495756 158714
rect 495728 151786 496124 151814
rect 496096 150226 496124 151786
rect 496740 150226 496768 159258
rect 497004 158772 497056 158778
rect 497004 158714 497056 158720
rect 497016 151814 497044 158714
rect 497016 151786 497412 151814
rect 497384 150226 497412 151786
rect 498028 150226 498056 159394
rect 498304 153202 498332 163200
rect 499132 163146 499160 163200
rect 499224 163146 499252 163254
rect 499132 163118 499252 163146
rect 498660 159384 498712 159390
rect 498660 159326 498712 159332
rect 498292 153196 498344 153202
rect 498292 153138 498344 153144
rect 498672 150226 498700 159326
rect 499500 158930 499528 163254
rect 499684 163254 499896 163282
rect 499500 158902 499620 158930
rect 499304 153196 499356 153202
rect 499304 153138 499356 153144
rect 499316 150226 499344 153138
rect 499592 151814 499620 158902
rect 499684 158778 499712 163254
rect 499868 163146 499896 163254
rect 499946 163200 500002 164400
rect 500866 163200 500922 164400
rect 501694 163200 501750 164400
rect 502522 163200 502578 164400
rect 503350 163200 503406 164400
rect 503824 163254 504128 163282
rect 499960 163146 499988 163200
rect 499868 163118 499988 163146
rect 500880 158794 500908 163200
rect 501708 161474 501736 163200
rect 501708 161446 501920 161474
rect 499672 158772 499724 158778
rect 499672 158714 499724 158720
rect 500592 158772 500644 158778
rect 500880 158766 501000 158794
rect 500592 158714 500644 158720
rect 499592 151786 499988 151814
rect 499960 150226 499988 151786
rect 500604 150226 500632 158714
rect 500972 151814 501000 158766
rect 500972 151786 501276 151814
rect 501248 150226 501276 151786
rect 501892 150226 501920 161446
rect 502536 150226 502564 163200
rect 503364 151814 503392 163200
rect 503272 151786 503392 151814
rect 503272 150226 503300 151786
rect 489920 150146 489972 150152
rect 489702 149940 489730 150146
rect 490346 149940 490374 150198
rect 490978 150204 491030 150210
rect 490978 150146 491030 150152
rect 491300 150204 491352 150210
rect 491588 150198 491662 150226
rect 491300 150146 491352 150152
rect 490990 149940 491018 150146
rect 491634 149940 491662 150198
rect 492266 150204 492318 150210
rect 492876 150198 492950 150226
rect 493520 150198 493594 150226
rect 494164 150198 494238 150226
rect 494808 150198 494882 150226
rect 495452 150198 495526 150226
rect 496096 150198 496170 150226
rect 496740 150198 496814 150226
rect 497384 150198 497458 150226
rect 498028 150198 498102 150226
rect 498672 150198 498746 150226
rect 499316 150198 499390 150226
rect 499960 150198 500034 150226
rect 500604 150198 500678 150226
rect 501248 150198 501322 150226
rect 501892 150198 501966 150226
rect 502536 150198 502610 150226
rect 492266 150146 492318 150152
rect 492278 149940 492306 150146
rect 492922 149940 492950 150198
rect 493566 149940 493594 150198
rect 494210 149940 494238 150198
rect 494854 149940 494882 150198
rect 495498 149940 495526 150198
rect 496142 149940 496170 150198
rect 496786 149940 496814 150198
rect 497430 149940 497458 150198
rect 498074 149940 498102 150198
rect 498718 149940 498746 150198
rect 499362 149940 499390 150198
rect 500006 149940 500034 150198
rect 500650 149940 500678 150198
rect 501294 149940 501322 150198
rect 501938 149940 501966 150198
rect 502582 149940 502610 150198
rect 503226 150198 503300 150226
rect 503824 150226 503852 163254
rect 504100 163146 504128 163254
rect 504178 163200 504234 164400
rect 505006 163200 505062 164400
rect 505112 163254 505784 163282
rect 504192 163146 504220 163200
rect 504100 163118 504220 163146
rect 505020 158778 505048 163200
rect 504456 158772 504508 158778
rect 504456 158714 504508 158720
rect 505008 158772 505060 158778
rect 505008 158714 505060 158720
rect 504468 150226 504496 158714
rect 505112 150226 505140 163254
rect 505756 163146 505784 163254
rect 505834 163200 505890 164400
rect 506754 163200 506810 164400
rect 507582 163200 507638 164400
rect 507872 163254 508360 163282
rect 505848 163146 505876 163200
rect 505756 163118 505876 163146
rect 506768 153202 506796 163200
rect 505836 153196 505888 153202
rect 505836 153138 505888 153144
rect 506756 153196 506808 153202
rect 506756 153138 506808 153144
rect 505848 150226 505876 153138
rect 507596 153134 507624 163200
rect 506388 153128 506440 153134
rect 506388 153070 506440 153076
rect 507584 153128 507636 153134
rect 507584 153070 507636 153076
rect 503824 150198 503898 150226
rect 504468 150198 504542 150226
rect 505112 150198 505186 150226
rect 503226 149940 503254 150198
rect 503870 149940 503898 150198
rect 504514 149940 504542 150198
rect 505158 149940 505186 150198
rect 505802 150198 505876 150226
rect 506400 150226 506428 153070
rect 507872 152386 507900 163254
rect 508332 163146 508360 163254
rect 508410 163200 508466 164400
rect 509238 163200 509294 164400
rect 510066 163200 510122 164400
rect 510894 163200 510950 164400
rect 511722 163200 511778 164400
rect 512012 163254 512592 163282
rect 508424 163146 508452 163200
rect 508332 163118 508452 163146
rect 507124 152380 507176 152386
rect 507124 152322 507176 152328
rect 507860 152380 507912 152386
rect 507860 152322 507912 152328
rect 507136 150226 507164 152322
rect 509252 151978 509280 163200
rect 509700 153196 509752 153202
rect 509700 153138 509752 153144
rect 507768 151972 507820 151978
rect 507768 151914 507820 151920
rect 509240 151972 509292 151978
rect 509240 151914 509292 151920
rect 507780 150226 507808 151914
rect 508412 151904 508464 151910
rect 508412 151846 508464 151852
rect 508424 150226 508452 151846
rect 509056 151836 509108 151842
rect 509056 151778 509108 151784
rect 509068 150226 509096 151778
rect 509712 150226 509740 153138
rect 510080 151910 510108 163200
rect 510344 152856 510396 152862
rect 510344 152798 510396 152804
rect 510068 151904 510120 151910
rect 510068 151846 510120 151852
rect 510356 150226 510384 152798
rect 510908 151842 510936 163200
rect 511736 153202 511764 163200
rect 511724 153196 511776 153202
rect 511724 153138 511776 153144
rect 510988 153128 511040 153134
rect 510988 153070 511040 153076
rect 510896 151836 510948 151842
rect 510896 151778 510948 151784
rect 511000 150226 511028 153070
rect 512012 152862 512040 163254
rect 512564 163146 512592 163254
rect 512642 163200 512698 164400
rect 513470 163200 513526 164400
rect 513576 163254 514248 163282
rect 512656 163146 512684 163200
rect 512564 163118 512684 163146
rect 512276 153196 512328 153202
rect 512276 153138 512328 153144
rect 512000 152856 512052 152862
rect 512000 152798 512052 152804
rect 511632 152380 511684 152386
rect 511632 152322 511684 152328
rect 511644 150226 511672 152322
rect 512288 150226 512316 153138
rect 513484 153134 513512 163200
rect 513472 153128 513524 153134
rect 513472 153070 513524 153076
rect 512920 153060 512972 153066
rect 512920 153002 512972 153008
rect 512932 150226 512960 153002
rect 513576 152386 513604 163254
rect 514220 163146 514248 163254
rect 514298 163200 514354 164400
rect 514864 163254 515076 163282
rect 514312 163146 514340 163200
rect 514220 163118 514340 163146
rect 514864 153202 514892 163254
rect 515048 163146 515076 163254
rect 515126 163200 515182 164400
rect 515954 163200 516010 164400
rect 516152 163254 516732 163282
rect 515140 163146 515168 163200
rect 515048 163118 515168 163146
rect 514852 153196 514904 153202
rect 514852 153138 514904 153144
rect 514208 153128 514260 153134
rect 514208 153070 514260 153076
rect 513564 152380 513616 152386
rect 513564 152322 513616 152328
rect 513564 152244 513616 152250
rect 513564 152186 513616 152192
rect 513576 150226 513604 152186
rect 514220 150226 514248 153070
rect 515968 153066 515996 163200
rect 515956 153060 516008 153066
rect 515956 153002 516008 153008
rect 514852 152992 514904 152998
rect 514852 152934 514904 152940
rect 514864 150226 514892 152934
rect 516152 152250 516180 163254
rect 516704 163146 516732 163254
rect 516782 163200 516838 164400
rect 517610 163200 517666 164400
rect 518530 163200 518586 164400
rect 519004 163254 519308 163282
rect 516796 163146 516824 163200
rect 516704 163118 516824 163146
rect 517624 153134 517652 163200
rect 517612 153128 517664 153134
rect 517612 153070 517664 153076
rect 518544 152998 518572 163200
rect 518532 152992 518584 152998
rect 518532 152934 518584 152940
rect 518072 152856 518124 152862
rect 518072 152798 518124 152804
rect 517428 152516 517480 152522
rect 517428 152458 517480 152464
rect 516140 152244 516192 152250
rect 516140 152186 516192 152192
rect 515496 152040 515548 152046
rect 515496 151982 515548 151988
rect 515508 150226 515536 151982
rect 516784 151972 516836 151978
rect 516784 151914 516836 151920
rect 516048 151836 516100 151842
rect 516048 151778 516100 151784
rect 506400 150198 506474 150226
rect 505802 149940 505830 150198
rect 506446 149940 506474 150198
rect 507090 150198 507164 150226
rect 507734 150198 507808 150226
rect 508378 150198 508452 150226
rect 509022 150198 509096 150226
rect 509666 150198 509740 150226
rect 510310 150198 510384 150226
rect 510954 150198 511028 150226
rect 511598 150198 511672 150226
rect 512242 150198 512316 150226
rect 512886 150198 512960 150226
rect 513530 150198 513604 150226
rect 514174 150198 514248 150226
rect 514818 150198 514892 150226
rect 515462 150198 515536 150226
rect 516060 150226 516088 151778
rect 516796 150226 516824 151914
rect 517440 150226 517468 152458
rect 518084 150226 518112 152798
rect 518808 152652 518860 152658
rect 518808 152594 518860 152600
rect 516060 150198 516134 150226
rect 507090 149940 507118 150198
rect 507734 149940 507762 150198
rect 508378 149940 508406 150198
rect 509022 149940 509050 150198
rect 509666 149940 509694 150198
rect 510310 149940 510338 150198
rect 510954 149940 510982 150198
rect 511598 149940 511626 150198
rect 512242 149940 512270 150198
rect 512886 149940 512914 150198
rect 513530 149940 513558 150198
rect 514174 149940 514202 150198
rect 514818 149940 514846 150198
rect 515462 149940 515490 150198
rect 516106 149940 516134 150198
rect 516750 150198 516824 150226
rect 517394 150198 517468 150226
rect 518038 150198 518112 150226
rect 516750 149940 516778 150198
rect 517394 149940 517422 150198
rect 518038 149940 518066 150198
rect 518820 149954 518848 152594
rect 519004 152046 519032 163254
rect 519280 163146 519308 163254
rect 519358 163200 519414 164400
rect 520186 163200 520242 164400
rect 520292 163254 520964 163282
rect 519372 163146 519400 163200
rect 519280 163118 519400 163146
rect 519542 161664 519598 161673
rect 519542 161599 519598 161608
rect 518992 152040 519044 152046
rect 518992 151982 519044 151988
rect 518696 149926 518848 149954
rect 117136 149796 117188 149802
rect 117136 149738 117188 149744
rect 117042 135552 117098 135561
rect 117042 135487 117098 135496
rect 117044 134564 117096 134570
rect 117044 134506 117096 134512
rect 116950 106856 117006 106865
rect 116950 106791 117006 106800
rect 117056 102921 117084 134506
rect 117148 127945 117176 149738
rect 519556 147937 519584 161599
rect 519634 160168 519690 160177
rect 519634 160103 519690 160112
rect 519542 147928 519598 147937
rect 519542 147863 519598 147872
rect 519648 146577 519676 160103
rect 520200 151842 520228 163200
rect 520292 151978 520320 163254
rect 520936 163146 520964 163254
rect 521014 163200 521070 164400
rect 521842 163200 521898 164400
rect 522670 163200 522726 164400
rect 523498 163200 523554 164400
rect 521028 163146 521056 163200
rect 520936 163118 521056 163146
rect 520922 163024 520978 163033
rect 520922 162959 520978 162968
rect 520280 151972 520332 151978
rect 520280 151914 520332 151920
rect 520188 151836 520240 151842
rect 520188 151778 520240 151784
rect 520936 149297 520964 162959
rect 521566 158672 521622 158681
rect 521566 158607 521622 158616
rect 521014 157176 521070 157185
rect 521014 157111 521070 157120
rect 520922 149288 520978 149297
rect 520922 149223 520978 149232
rect 520922 148064 520978 148073
rect 520922 147999 520978 148008
rect 519634 146568 519690 146577
rect 519634 146503 519690 146512
rect 519818 146568 519874 146577
rect 519818 146503 519874 146512
rect 519542 144936 519598 144945
rect 519542 144871 519598 144880
rect 519556 132977 519584 144871
rect 519832 134337 519860 146503
rect 520738 143440 520794 143449
rect 520738 143375 520794 143384
rect 519818 134328 519874 134337
rect 519818 134263 519874 134272
rect 519542 132968 519598 132977
rect 519542 132903 519598 132912
rect 520752 131481 520780 143375
rect 520830 141944 520886 141953
rect 520830 141879 520886 141888
rect 520738 131472 520794 131481
rect 520738 131407 520794 131416
rect 520844 130121 520872 141879
rect 520936 135697 520964 147999
rect 521028 143857 521056 157111
rect 521290 155680 521346 155689
rect 521290 155615 521346 155624
rect 521198 151056 521254 151065
rect 521198 150991 521254 151000
rect 521106 149560 521162 149569
rect 521106 149495 521162 149504
rect 521014 143848 521070 143857
rect 521014 143783 521070 143792
rect 521120 137057 521148 149495
rect 521212 138417 521240 150991
rect 521304 142497 521332 155615
rect 521474 154048 521530 154057
rect 521474 153983 521530 153992
rect 521382 152552 521438 152561
rect 521382 152487 521438 152496
rect 521290 142488 521346 142497
rect 521290 142423 521346 142432
rect 521396 139777 521424 152487
rect 521488 141137 521516 153983
rect 521580 145217 521608 158607
rect 521856 152522 521884 163200
rect 522684 152862 522712 163200
rect 522672 152856 522724 152862
rect 522672 152798 522724 152804
rect 523512 152658 523540 163200
rect 523500 152652 523552 152658
rect 523500 152594 523552 152600
rect 521844 152516 521896 152522
rect 521844 152458 521896 152464
rect 521566 145208 521622 145217
rect 521566 145143 521622 145152
rect 521474 141128 521530 141137
rect 521474 141063 521530 141072
rect 521566 140448 521622 140457
rect 521566 140383 521622 140392
rect 521382 139768 521438 139777
rect 521382 139703 521438 139712
rect 521382 138952 521438 138961
rect 521382 138887 521438 138896
rect 521198 138408 521254 138417
rect 521198 138343 521254 138352
rect 521106 137048 521162 137057
rect 521106 136983 521162 136992
rect 521290 135824 521346 135833
rect 521290 135759 521346 135768
rect 520922 135688 520978 135697
rect 520922 135623 520978 135632
rect 521198 134328 521254 134337
rect 521198 134263 521254 134272
rect 521106 132832 521162 132841
rect 521106 132767 521162 132776
rect 520922 131336 520978 131345
rect 520922 131271 520978 131280
rect 520830 130112 520886 130121
rect 520830 130047 520886 130056
rect 520830 128344 520886 128353
rect 520830 128279 520886 128288
rect 117134 127936 117190 127945
rect 117134 127871 117190 127880
rect 520738 126712 520794 126721
rect 520738 126647 520794 126656
rect 520752 116521 520780 126647
rect 520844 117881 520872 128279
rect 520936 120601 520964 131271
rect 521014 129840 521070 129849
rect 521014 129775 521070 129784
rect 520922 120592 520978 120601
rect 520922 120527 520978 120536
rect 521028 119241 521056 129775
rect 521120 121961 521148 132767
rect 521212 123321 521240 134263
rect 521304 124681 521332 135759
rect 521396 127401 521424 138887
rect 521474 137456 521530 137465
rect 521474 137391 521530 137400
rect 521382 127392 521438 127401
rect 521382 127327 521438 127336
rect 521488 126041 521516 137391
rect 521580 128761 521608 140383
rect 521566 128752 521622 128761
rect 521566 128687 521622 128696
rect 521474 126032 521530 126041
rect 521474 125967 521530 125976
rect 521474 125216 521530 125225
rect 521474 125151 521530 125160
rect 521290 124672 521346 124681
rect 521290 124607 521346 124616
rect 521382 123720 521438 123729
rect 521382 123655 521438 123664
rect 521198 123312 521254 123321
rect 521198 123247 521254 123256
rect 521290 122224 521346 122233
rect 521290 122159 521346 122168
rect 521106 121952 521162 121961
rect 521106 121887 521162 121896
rect 521014 119232 521070 119241
rect 521014 119167 521070 119176
rect 521198 119232 521254 119241
rect 521198 119167 521254 119176
rect 520830 117872 520886 117881
rect 520830 117807 520886 117816
rect 521014 117600 521070 117609
rect 521014 117535 521070 117544
rect 520738 116512 520794 116521
rect 520738 116447 520794 116456
rect 520922 116104 520978 116113
rect 520922 116039 520978 116048
rect 520738 113112 520794 113121
rect 520738 113047 520794 113056
rect 520278 105496 520334 105505
rect 520278 105431 520334 105440
rect 117042 102912 117098 102921
rect 117042 102847 117098 102856
rect 116858 101008 116914 101017
rect 116858 100943 116914 100952
rect 116766 99104 116822 99113
rect 116766 99039 116822 99048
rect 520292 97345 520320 105431
rect 520752 104145 520780 113047
rect 520830 111616 520886 111625
rect 520830 111551 520886 111560
rect 520738 104136 520794 104145
rect 520738 104071 520794 104080
rect 520844 102785 520872 111551
rect 520936 106865 520964 116039
rect 521028 108225 521056 117535
rect 521106 114608 521162 114617
rect 521106 114543 521162 114552
rect 521014 108216 521070 108225
rect 521014 108151 521070 108160
rect 520922 106856 520978 106865
rect 520922 106791 520978 106800
rect 521120 105641 521148 114543
rect 521212 109585 521240 119167
rect 521304 112305 521332 122159
rect 521396 113801 521424 123655
rect 521488 115161 521516 125151
rect 521566 120728 521622 120737
rect 521566 120663 521622 120672
rect 521474 115152 521530 115161
rect 521474 115087 521530 115096
rect 521382 113792 521438 113801
rect 521382 113727 521438 113736
rect 521290 112296 521346 112305
rect 521290 112231 521346 112240
rect 521580 110945 521608 120663
rect 521566 110936 521622 110945
rect 521566 110871 521622 110880
rect 521566 110120 521622 110129
rect 521566 110055 521622 110064
rect 521198 109576 521254 109585
rect 521198 109511 521254 109520
rect 521198 108488 521254 108497
rect 521198 108423 521254 108432
rect 521106 105632 521162 105641
rect 521106 105567 521162 105576
rect 521106 104000 521162 104009
rect 521106 103935 521162 103944
rect 520830 102776 520886 102785
rect 520830 102711 520886 102720
rect 521014 102504 521070 102513
rect 521014 102439 521070 102448
rect 520922 101008 520978 101017
rect 520922 100943 520978 100952
rect 520830 97880 520886 97889
rect 520830 97815 520886 97824
rect 520278 97336 520334 97345
rect 520278 97271 520334 97280
rect 116768 96892 116820 96898
rect 116768 96834 116820 96840
rect 116674 95296 116730 95305
rect 116674 95231 116730 95240
rect 116492 93628 116544 93634
rect 116492 93570 116544 93576
rect 116504 93401 116532 93570
rect 116490 93392 116546 93401
rect 116490 93327 116546 93336
rect 116124 92472 116176 92478
rect 116124 92414 116176 92420
rect 116136 91361 116164 92414
rect 116122 91352 116178 91361
rect 116122 91287 116178 91296
rect 116676 87236 116728 87242
rect 116676 87178 116728 87184
rect 116216 86964 116268 86970
rect 116216 86906 116268 86912
rect 116228 85649 116256 86906
rect 116214 85640 116270 85649
rect 116214 85575 116270 85584
rect 115386 81832 115442 81841
rect 115386 81767 115442 81776
rect 116688 78033 116716 87178
rect 116780 79937 116808 96834
rect 520370 96384 520426 96393
rect 520370 96319 520426 96328
rect 520278 94888 520334 94897
rect 520278 94823 520334 94832
rect 116860 91656 116912 91662
rect 116860 91598 116912 91604
rect 116872 87553 116900 91598
rect 520292 87689 520320 94823
rect 520384 89049 520412 96319
rect 520738 93392 520794 93401
rect 520738 93327 520794 93336
rect 520370 89040 520426 89049
rect 520370 88975 520426 88984
rect 520278 87680 520334 87689
rect 520278 87615 520334 87624
rect 116858 87544 116914 87553
rect 116858 87479 116914 87488
rect 520752 86329 520780 93327
rect 520844 90409 520872 97815
rect 520936 93129 520964 100943
rect 521028 94489 521056 102439
rect 521120 95985 521148 103935
rect 521212 100065 521240 108423
rect 521382 106992 521438 107001
rect 521382 106927 521438 106936
rect 521198 100056 521254 100065
rect 521198 99991 521254 100000
rect 521198 99376 521254 99385
rect 521198 99311 521254 99320
rect 521106 95976 521162 95985
rect 521106 95911 521162 95920
rect 521014 94480 521070 94489
rect 521014 94415 521070 94424
rect 520922 93120 520978 93129
rect 520922 93055 520978 93064
rect 521014 91896 521070 91905
rect 521014 91831 521070 91840
rect 520830 90400 520886 90409
rect 520830 90335 520886 90344
rect 520738 86320 520794 86329
rect 520738 86255 520794 86264
rect 520370 85776 520426 85785
rect 520370 85711 520426 85720
rect 520278 84280 520334 84289
rect 520278 84215 520334 84224
rect 116766 79928 116822 79937
rect 116766 79863 116822 79872
rect 520292 78169 520320 84215
rect 520384 79529 520412 85711
rect 521028 84969 521056 91831
rect 521212 91769 521240 99311
rect 521396 98705 521424 106927
rect 521580 101425 521608 110055
rect 521566 101416 521622 101425
rect 521566 101351 521622 101360
rect 521382 98696 521438 98705
rect 521382 98631 521438 98640
rect 521198 91760 521254 91769
rect 521198 91695 521254 91704
rect 521198 90264 521254 90273
rect 521198 90199 521254 90208
rect 521106 87272 521162 87281
rect 521106 87207 521162 87216
rect 521014 84960 521070 84969
rect 521014 84895 521070 84904
rect 520738 82784 520794 82793
rect 520738 82719 520794 82728
rect 520370 79520 520426 79529
rect 520370 79455 520426 79464
rect 520278 78160 520334 78169
rect 520278 78095 520334 78104
rect 116674 78024 116730 78033
rect 116674 77959 116730 77968
rect 520752 76809 520780 82719
rect 521014 81152 521070 81161
rect 521014 81087 521070 81096
rect 520738 76800 520794 76809
rect 520738 76735 520794 76744
rect 520462 76664 520518 76673
rect 520462 76599 520518 76608
rect 520278 75168 520334 75177
rect 520278 75103 520334 75112
rect 116582 74080 116638 74089
rect 116582 74015 116638 74024
rect 116398 72176 116454 72185
rect 116398 72111 116454 72120
rect 116412 71806 116440 72111
rect 113824 71800 113876 71806
rect 113824 71742 113876 71748
rect 116400 71800 116452 71806
rect 116400 71742 116452 71748
rect 112444 62144 112496 62150
rect 112444 62086 112496 62092
rect 111064 59424 111116 59430
rect 111064 59366 111116 59372
rect 109684 37324 109736 37330
rect 109684 37266 109736 37272
rect 109592 4548 109644 4554
rect 109592 4490 109644 4496
rect 2504 2848 2556 2854
rect 2504 2790 2556 2796
rect 2516 2666 2544 2790
rect 109604 2666 109632 4490
rect 2516 2638 2714 2666
rect 106030 2650 106228 2666
rect 32772 2644 32824 2650
rect 32772 2586 32824 2592
rect 98276 2644 98328 2650
rect 106030 2644 106240 2650
rect 106030 2638 106188 2644
rect 98276 2586 98328 2592
rect 109342 2638 109632 2666
rect 106188 2586 106240 2592
rect 29550 2136 29606 2145
rect 6012 1601 6040 2108
rect 5998 1592 6054 1601
rect 5998 1527 6054 1536
rect 9324 1426 9352 2108
rect 12636 1494 12664 2108
rect 15948 1873 15976 2108
rect 15934 1864 15990 1873
rect 15934 1799 15990 1808
rect 19352 1737 19380 2108
rect 19338 1728 19394 1737
rect 19338 1663 19394 1672
rect 12624 1488 12676 1494
rect 12624 1430 12676 1436
rect 9312 1420 9364 1426
rect 9312 1362 9364 1368
rect 22664 814 22692 2108
rect 25990 2094 26096 2122
rect 29302 2094 29550 2122
rect 26068 2009 26096 2094
rect 29550 2071 29606 2080
rect 26054 2000 26110 2009
rect 26054 1935 26110 1944
rect 32692 1562 32720 2108
rect 32680 1556 32732 1562
rect 32680 1498 32732 1504
rect 22652 808 22704 814
rect 32784 800 32812 2586
rect 42706 2272 42762 2281
rect 42642 2230 42706 2258
rect 42706 2207 42762 2216
rect 93032 2168 93084 2174
rect 36004 1290 36032 2108
rect 35992 1284 36044 1290
rect 35992 1226 36044 1232
rect 39316 1222 39344 2108
rect 46032 1698 46060 2108
rect 46020 1692 46072 1698
rect 46020 1634 46072 1640
rect 49344 1630 49372 2108
rect 52656 1766 52684 2108
rect 52644 1760 52696 1766
rect 52644 1702 52696 1708
rect 49332 1624 49384 1630
rect 49332 1566 49384 1572
rect 55968 1465 55996 2108
rect 59372 1834 59400 2108
rect 59360 1828 59412 1834
rect 59360 1770 59412 1776
rect 55954 1456 56010 1465
rect 55954 1391 56010 1400
rect 39304 1216 39356 1222
rect 39304 1158 39356 1164
rect 62684 1154 62712 2108
rect 65996 1902 66024 2108
rect 65984 1896 66036 1902
rect 65984 1838 66036 1844
rect 62672 1148 62724 1154
rect 62672 1090 62724 1096
rect 69308 1086 69336 2108
rect 72712 1970 72740 2108
rect 72700 1964 72752 1970
rect 72700 1906 72752 1912
rect 69296 1080 69348 1086
rect 69296 1022 69348 1028
rect 76024 1018 76052 2108
rect 79350 2094 79640 2122
rect 79612 2038 79640 2094
rect 79600 2032 79652 2038
rect 79600 1974 79652 1980
rect 76012 1012 76064 1018
rect 76012 954 76064 960
rect 82648 950 82676 2108
rect 86066 2106 86448 2122
rect 92690 2116 93032 2122
rect 92690 2110 93084 2116
rect 86066 2100 86460 2106
rect 86066 2094 86408 2100
rect 86408 2042 86460 2048
rect 82636 944 82688 950
rect 82636 886 82688 892
rect 89364 882 89392 2108
rect 92690 2094 93072 2110
rect 95988 1358 96016 2108
rect 98000 1488 98052 1494
rect 98000 1430 98052 1436
rect 95976 1352 96028 1358
rect 98012 1329 98040 1430
rect 95976 1294 96028 1300
rect 97998 1320 98054 1329
rect 97998 1255 98054 1264
rect 89352 876 89404 882
rect 89352 818 89404 824
rect 98288 800 98316 2586
rect 99392 1494 99420 2108
rect 99380 1488 99432 1494
rect 99380 1430 99432 1436
rect 102704 1426 102732 2108
rect 109696 1902 109724 37266
rect 109776 33176 109828 33182
rect 109776 33118 109828 33124
rect 109684 1896 109736 1902
rect 109684 1838 109736 1844
rect 109788 1834 109816 33118
rect 109868 4888 109920 4894
rect 109868 4830 109920 4836
rect 109880 1970 109908 4830
rect 109960 4820 110012 4826
rect 109960 4762 110012 4768
rect 109868 1964 109920 1970
rect 109868 1906 109920 1912
rect 109972 1873 110000 4762
rect 111076 2650 111104 59366
rect 111248 22840 111300 22846
rect 111248 22782 111300 22788
rect 111156 22772 111208 22778
rect 111156 22714 111208 22720
rect 111064 2644 111116 2650
rect 111064 2586 111116 2592
rect 109958 1864 110014 1873
rect 109776 1828 109828 1834
rect 109958 1799 110014 1808
rect 109776 1770 109828 1776
rect 111168 1494 111196 22714
rect 111156 1488 111208 1494
rect 111156 1430 111208 1436
rect 111260 1426 111288 22782
rect 111340 19372 111392 19378
rect 111340 19314 111392 19320
rect 111352 1562 111380 19314
rect 111432 18012 111484 18018
rect 111432 17954 111484 17960
rect 111444 2145 111472 17954
rect 111616 15224 111668 15230
rect 111616 15166 111668 15172
rect 111524 3052 111576 3058
rect 111524 2994 111576 3000
rect 111430 2136 111486 2145
rect 111430 2071 111486 2080
rect 111340 1556 111392 1562
rect 111340 1498 111392 1504
rect 111536 1426 111564 2994
rect 111628 2009 111656 15166
rect 112456 4554 112484 62086
rect 113836 53145 113864 71742
rect 116306 70272 116362 70281
rect 116306 70207 116362 70216
rect 116320 69086 116348 70207
rect 114100 69080 114152 69086
rect 114100 69022 114152 69028
rect 116308 69080 116360 69086
rect 116308 69022 116360 69028
rect 113822 53136 113878 53145
rect 113822 53071 113878 53080
rect 113824 51128 113876 51134
rect 113824 51070 113876 51076
rect 112536 27668 112588 27674
rect 112536 27610 112588 27616
rect 112444 4548 112496 4554
rect 112444 4490 112496 4496
rect 111614 2000 111670 2009
rect 111614 1935 111670 1944
rect 112548 1698 112576 27610
rect 112628 23520 112680 23526
rect 112628 23462 112680 23468
rect 112536 1692 112588 1698
rect 112536 1634 112588 1640
rect 100760 1420 100812 1426
rect 100760 1362 100812 1368
rect 102692 1420 102744 1426
rect 102692 1362 102744 1368
rect 111248 1420 111300 1426
rect 111248 1362 111300 1368
rect 111524 1420 111576 1426
rect 111524 1362 111576 1368
rect 100772 1193 100800 1362
rect 112640 1222 112668 23462
rect 112720 22160 112772 22166
rect 112720 22102 112772 22108
rect 112732 1290 112760 22102
rect 112720 1284 112772 1290
rect 112720 1226 112772 1232
rect 112628 1216 112680 1222
rect 100758 1184 100814 1193
rect 112628 1158 112680 1164
rect 100758 1119 100814 1128
rect 113836 882 113864 51070
rect 113916 46980 113968 46986
rect 113916 46922 113968 46928
rect 113928 950 113956 46922
rect 114008 42832 114060 42838
rect 114008 42774 114060 42780
rect 114020 1018 114048 42774
rect 114112 41857 114140 69022
rect 116214 68368 116270 68377
rect 116214 68303 116270 68312
rect 116228 67658 116256 68303
rect 114192 67652 114244 67658
rect 114192 67594 114244 67600
rect 116216 67652 116268 67658
rect 116216 67594 116268 67600
rect 114098 41848 114154 41857
rect 114098 41783 114154 41792
rect 114100 38684 114152 38690
rect 114100 38626 114152 38632
rect 114112 1086 114140 38626
rect 114204 30433 114232 67594
rect 116596 64734 116624 74015
rect 520292 69873 520320 75103
rect 520476 71233 520504 76599
rect 521028 75313 521056 81087
rect 521120 80889 521148 87207
rect 521212 83609 521240 90199
rect 521290 88768 521346 88777
rect 521290 88703 521346 88712
rect 521198 83600 521254 83609
rect 521198 83535 521254 83544
rect 521304 82249 521332 88703
rect 521290 82240 521346 82249
rect 521290 82175 521346 82184
rect 521106 80880 521162 80889
rect 521106 80815 521162 80824
rect 521382 79656 521438 79665
rect 521382 79591 521438 79600
rect 521106 78160 521162 78169
rect 521106 78095 521162 78104
rect 521014 75304 521070 75313
rect 521014 75239 521070 75248
rect 520738 73672 520794 73681
rect 520738 73607 520794 73616
rect 520462 71224 520518 71233
rect 520462 71159 520518 71168
rect 520278 69864 520334 69873
rect 520278 69799 520334 69808
rect 520752 68513 520780 73607
rect 521120 72593 521148 78095
rect 521396 73953 521424 79591
rect 521382 73944 521438 73953
rect 521382 73879 521438 73888
rect 521106 72584 521162 72593
rect 521106 72519 521162 72528
rect 521014 72040 521070 72049
rect 521014 71975 521070 71984
rect 520738 68504 520794 68513
rect 520738 68439 520794 68448
rect 520462 67552 520518 67561
rect 520462 67487 520518 67496
rect 116858 66464 116914 66473
rect 116858 66399 116914 66408
rect 114468 64728 114520 64734
rect 114468 64670 114520 64676
rect 116584 64728 116636 64734
rect 116584 64670 116636 64676
rect 114480 64569 114508 64670
rect 114466 64560 114522 64569
rect 114466 64495 114522 64504
rect 115202 64560 115258 64569
rect 115202 64495 115258 64504
rect 114284 48272 114336 48278
rect 114284 48214 114336 48220
rect 114190 30424 114246 30433
rect 114190 30359 114246 30368
rect 114296 19009 114324 48214
rect 114282 19000 114338 19009
rect 114282 18935 114338 18944
rect 114284 13864 114336 13870
rect 114284 13806 114336 13812
rect 114192 8016 114244 8022
rect 114192 7958 114244 7964
rect 114204 7721 114232 7958
rect 114190 7712 114246 7721
rect 114190 7647 114246 7656
rect 114296 6914 114324 13806
rect 115216 8022 115244 64495
rect 116122 62656 116178 62665
rect 116122 62591 116178 62600
rect 116136 62150 116164 62591
rect 116124 62144 116176 62150
rect 116124 62086 116176 62092
rect 116122 60616 116178 60625
rect 116122 60551 116178 60560
rect 116136 59430 116164 60551
rect 116124 59424 116176 59430
rect 116124 59366 116176 59372
rect 116582 54904 116638 54913
rect 116582 54839 116638 54848
rect 115940 51128 115992 51134
rect 115938 51096 115940 51105
rect 115992 51096 115994 51105
rect 115938 51031 115994 51040
rect 116030 47152 116086 47161
rect 116030 47087 116086 47096
rect 116044 46986 116072 47087
rect 116032 46980 116084 46986
rect 116032 46922 116084 46928
rect 116398 43344 116454 43353
rect 116398 43279 116454 43288
rect 116412 42838 116440 43279
rect 116400 42832 116452 42838
rect 116400 42774 116452 42780
rect 115938 39536 115994 39545
rect 115938 39471 115994 39480
rect 115952 38690 115980 39471
rect 115940 38684 115992 38690
rect 115940 38626 115992 38632
rect 116122 37632 116178 37641
rect 116122 37567 116178 37576
rect 116136 37330 116164 37567
rect 116124 37324 116176 37330
rect 116124 37266 116176 37272
rect 116122 33824 116178 33833
rect 116122 33759 116178 33768
rect 116136 33182 116164 33759
rect 116124 33176 116176 33182
rect 116124 33118 116176 33124
rect 116490 31784 116546 31793
rect 116490 31719 116546 31728
rect 116308 31068 116360 31074
rect 116308 31010 116360 31016
rect 116122 27976 116178 27985
rect 116122 27911 116178 27920
rect 116136 27674 116164 27911
rect 116124 27668 116176 27674
rect 116124 27610 116176 27616
rect 116122 24168 116178 24177
rect 116122 24103 116178 24112
rect 116136 23526 116164 24103
rect 116124 23520 116176 23526
rect 116124 23462 116176 23468
rect 116320 22778 116348 31010
rect 116398 29880 116454 29889
rect 116398 29815 116454 29824
rect 116308 22772 116360 22778
rect 116308 22714 116360 22720
rect 116122 22264 116178 22273
rect 116122 22199 116178 22208
rect 116136 22166 116164 22199
rect 116124 22160 116176 22166
rect 116124 22102 116176 22108
rect 116122 20360 116178 20369
rect 116122 20295 116178 20304
rect 116136 19378 116164 20295
rect 116124 19372 116176 19378
rect 116124 19314 116176 19320
rect 116122 18456 116178 18465
rect 116122 18391 116178 18400
rect 116136 18018 116164 18391
rect 116124 18012 116176 18018
rect 116124 17954 116176 17960
rect 116122 16416 116178 16425
rect 116122 16351 116178 16360
rect 116136 15230 116164 16351
rect 116124 15224 116176 15230
rect 116124 15166 116176 15172
rect 115938 14512 115994 14521
rect 115938 14447 115994 14456
rect 115952 13870 115980 14447
rect 115940 13864 115992 13870
rect 115940 13806 115992 13812
rect 115204 8016 115256 8022
rect 115204 7958 115256 7964
rect 114204 6886 114324 6914
rect 114100 1080 114152 1086
rect 114100 1022 114152 1028
rect 114008 1012 114060 1018
rect 114008 954 114060 960
rect 113916 944 113968 950
rect 113916 886 113968 892
rect 113824 876 113876 882
rect 113824 818 113876 824
rect 114204 814 114232 6886
rect 116030 4992 116086 5001
rect 116030 4927 116086 4936
rect 116044 1601 116072 4927
rect 116122 3088 116178 3097
rect 116122 3023 116178 3032
rect 116136 2854 116164 3023
rect 116124 2848 116176 2854
rect 116124 2790 116176 2796
rect 116412 1630 116440 29815
rect 116504 1766 116532 31719
rect 116492 1760 116544 1766
rect 116492 1702 116544 1708
rect 116400 1624 116452 1630
rect 116030 1592 116086 1601
rect 116400 1566 116452 1572
rect 116030 1527 116086 1536
rect 116596 1358 116624 54839
rect 116674 53000 116730 53009
rect 116674 52935 116730 52944
rect 116688 2174 116716 52935
rect 116766 49192 116822 49201
rect 116766 49127 116822 49136
rect 116676 2168 116728 2174
rect 116676 2110 116728 2116
rect 116780 2106 116808 49127
rect 116872 48278 116900 66399
rect 520370 66056 520426 66065
rect 520370 65991 520426 66000
rect 520384 61713 520412 65991
rect 520476 63073 520504 67487
rect 521028 67153 521056 71975
rect 521106 70544 521162 70553
rect 521106 70479 521162 70488
rect 521014 67144 521070 67153
rect 521014 67079 521070 67088
rect 521120 65793 521148 70479
rect 521290 69048 521346 69057
rect 521290 68983 521346 68992
rect 521106 65784 521162 65793
rect 521106 65719 521162 65728
rect 520738 64560 520794 64569
rect 520738 64495 520794 64504
rect 520462 63064 520518 63073
rect 520462 62999 520518 63008
rect 520370 61704 520426 61713
rect 520370 61639 520426 61648
rect 520752 60353 520780 64495
rect 521304 64433 521332 68983
rect 521290 64424 521346 64433
rect 521290 64359 521346 64368
rect 521106 62928 521162 62937
rect 521106 62863 521162 62872
rect 521014 61432 521070 61441
rect 521014 61367 521070 61376
rect 520738 60344 520794 60353
rect 520738 60279 520794 60288
rect 520738 59936 520794 59945
rect 520738 59871 520794 59880
rect 117042 58712 117098 58721
rect 117042 58647 117098 58656
rect 116860 48272 116912 48278
rect 116860 48214 116912 48220
rect 116858 45248 116914 45257
rect 116858 45183 116914 45192
rect 116768 2100 116820 2106
rect 116768 2042 116820 2048
rect 116872 2038 116900 45183
rect 116950 41440 117006 41449
rect 116950 41375 117006 41384
rect 116964 4894 116992 41375
rect 117056 22846 117084 58647
rect 520370 56944 520426 56953
rect 520370 56879 520426 56888
rect 117134 56808 117190 56817
rect 117134 56743 117190 56752
rect 117148 55214 117176 56743
rect 520278 55448 520334 55457
rect 520278 55383 520334 55392
rect 117148 55186 117268 55214
rect 117134 35728 117190 35737
rect 117134 35663 117190 35672
rect 117044 22840 117096 22846
rect 117044 22782 117096 22788
rect 117042 12608 117098 12617
rect 117042 12543 117098 12552
rect 116952 4888 117004 4894
rect 116952 4830 117004 4836
rect 116860 2032 116912 2038
rect 116860 1974 116912 1980
rect 117056 1737 117084 12543
rect 117042 1728 117098 1737
rect 117042 1663 117098 1672
rect 116584 1352 116636 1358
rect 116584 1294 116636 1300
rect 117148 1154 117176 35663
rect 117240 31074 117268 55186
rect 520292 52057 520320 55383
rect 520384 53417 520412 56879
rect 520752 56137 520780 59871
rect 521028 57497 521056 61367
rect 521120 58993 521148 62863
rect 521106 58984 521162 58993
rect 521106 58919 521162 58928
rect 521106 58440 521162 58449
rect 521106 58375 521162 58384
rect 521014 57488 521070 57497
rect 521014 57423 521070 57432
rect 520738 56128 520794 56137
rect 520738 56063 520794 56072
rect 521120 54777 521148 58375
rect 521106 54768 521162 54777
rect 521106 54703 521162 54712
rect 521106 53816 521162 53825
rect 521106 53751 521162 53760
rect 520370 53408 520426 53417
rect 520370 53343 520426 53352
rect 520922 52320 520978 52329
rect 520922 52255 520978 52264
rect 520278 52048 520334 52057
rect 520278 51983 520334 51992
rect 520370 50824 520426 50833
rect 520370 50759 520426 50768
rect 520384 47977 520412 50759
rect 520936 49337 520964 52255
rect 521120 50697 521148 53751
rect 521106 50688 521162 50697
rect 521106 50623 521162 50632
rect 520922 49328 520978 49337
rect 520922 49263 520978 49272
rect 521106 49328 521162 49337
rect 521106 49263 521162 49272
rect 520370 47968 520426 47977
rect 520370 47903 520426 47912
rect 520278 47832 520334 47841
rect 520278 47767 520334 47776
rect 520292 45257 520320 47767
rect 521120 46617 521148 49263
rect 521106 46608 521162 46617
rect 521106 46543 521162 46552
rect 520370 46336 520426 46345
rect 520370 46271 520426 46280
rect 520278 45248 520334 45257
rect 520278 45183 520334 45192
rect 520384 43897 520412 46271
rect 521014 44704 521070 44713
rect 521014 44639 521070 44648
rect 520370 43888 520426 43897
rect 520370 43823 520426 43832
rect 521028 42537 521056 44639
rect 521106 43208 521162 43217
rect 521106 43143 521162 43152
rect 521014 42528 521070 42537
rect 521014 42463 521070 42472
rect 521014 41712 521070 41721
rect 521014 41647 521070 41656
rect 521028 39817 521056 41647
rect 521120 41177 521148 43143
rect 521106 41168 521162 41177
rect 521106 41103 521162 41112
rect 521106 40216 521162 40225
rect 521106 40151 521162 40160
rect 521014 39808 521070 39817
rect 521014 39743 521070 39752
rect 520922 38720 520978 38729
rect 520922 38655 520978 38664
rect 520936 36961 520964 38655
rect 521120 38321 521148 40151
rect 521106 38312 521162 38321
rect 521106 38247 521162 38256
rect 521106 37224 521162 37233
rect 521106 37159 521162 37168
rect 520922 36952 520978 36961
rect 520922 36887 520978 36896
rect 521120 36009 521148 37159
rect 521106 36000 521162 36009
rect 521106 35935 521162 35944
rect 520922 35592 520978 35601
rect 520922 35527 520978 35536
rect 520936 34649 520964 35527
rect 520922 34640 520978 34649
rect 520922 34575 520978 34584
rect 520830 34096 520886 34105
rect 520830 34031 520886 34040
rect 520844 33289 520872 34031
rect 520830 33280 520886 33289
rect 520830 33215 520886 33224
rect 521106 32600 521162 32609
rect 521106 32535 521162 32544
rect 521120 31793 521148 32535
rect 521106 31784 521162 31793
rect 521106 31719 521162 31728
rect 521106 31104 521162 31113
rect 117228 31068 117280 31074
rect 521106 31039 521162 31048
rect 117228 31010 117280 31016
rect 521120 30433 521148 31039
rect 521106 30424 521162 30433
rect 521106 30359 521162 30368
rect 521106 29608 521162 29617
rect 521106 29543 521162 29552
rect 521120 28801 521148 29543
rect 521106 28792 521162 28801
rect 521106 28727 521162 28736
rect 521106 20496 521162 20505
rect 521106 20431 521162 20440
rect 521120 19825 521148 20431
rect 521106 19816 521162 19825
rect 521106 19751 521162 19760
rect 521106 15056 521162 15065
rect 521106 14991 521162 15000
rect 521120 14385 521148 14991
rect 521106 14376 521162 14385
rect 521106 14311 521162 14320
rect 521106 13696 521162 13705
rect 521106 13631 521162 13640
rect 521120 12889 521148 13631
rect 521106 12880 521162 12889
rect 521106 12815 521162 12824
rect 519634 12336 519690 12345
rect 519634 12271 519690 12280
rect 519648 11393 519676 12271
rect 519634 11384 519690 11393
rect 519634 11319 519690 11328
rect 521106 10976 521162 10985
rect 521106 10911 521162 10920
rect 117226 10704 117282 10713
rect 117226 10639 117282 10648
rect 117240 4826 117268 10639
rect 521120 9897 521148 10911
rect 521106 9888 521162 9897
rect 521106 9823 521162 9832
rect 521106 9616 521162 9625
rect 521106 9551 521162 9560
rect 521120 8265 521148 9551
rect 520370 8256 520426 8265
rect 520370 8191 520426 8200
rect 521106 8256 521162 8265
rect 521106 8191 521162 8200
rect 520384 6769 520412 8191
rect 521106 6896 521162 6905
rect 521106 6831 521162 6840
rect 520370 6760 520426 6769
rect 520370 6695 520426 6704
rect 521014 5536 521070 5545
rect 521014 5471 521070 5480
rect 117228 4820 117280 4826
rect 117228 4762 117280 4768
rect 520922 4176 520978 4185
rect 520922 4111 520978 4120
rect 118700 2984 118752 2990
rect 118700 2926 118752 2932
rect 118712 1494 118740 2926
rect 520936 2281 520964 4111
rect 521028 3777 521056 5471
rect 521120 5273 521148 6831
rect 521106 5264 521162 5273
rect 521106 5199 521162 5208
rect 521014 3768 521070 3777
rect 521014 3703 521070 3712
rect 521106 2816 521162 2825
rect 521106 2751 521162 2760
rect 520922 2272 520978 2281
rect 520922 2207 520978 2216
rect 143644 2094 143980 2122
rect 193600 2094 193936 2122
rect 243648 2094 243984 2122
rect 293604 2094 293940 2122
rect 143644 1494 143672 2094
rect 118700 1488 118752 1494
rect 118700 1430 118752 1436
rect 143632 1488 143684 1494
rect 143632 1430 143684 1436
rect 193600 1426 193628 2094
rect 243648 1426 243676 2094
rect 293604 1426 293632 2094
rect 343974 1873 344002 2108
rect 393944 2094 394280 2122
rect 443992 2094 444328 2122
rect 343960 1864 344016 1873
rect 343960 1799 344016 1808
rect 394252 1494 394280 2094
rect 444300 1494 444328 2094
rect 493612 2094 493948 2122
rect 394240 1488 394292 1494
rect 294786 1456 294842 1465
rect 193588 1420 193640 1426
rect 193588 1362 193640 1368
rect 193680 1420 193732 1426
rect 193680 1362 193732 1368
rect 243636 1420 243688 1426
rect 243636 1362 243688 1368
rect 243728 1420 243780 1426
rect 243728 1362 243780 1368
rect 293592 1420 293644 1426
rect 294786 1391 294842 1400
rect 295338 1456 295394 1465
rect 394240 1430 394292 1436
rect 425796 1488 425848 1494
rect 425796 1430 425848 1436
rect 444288 1488 444340 1494
rect 444288 1430 444340 1436
rect 491300 1488 491352 1494
rect 491300 1430 491352 1436
rect 295338 1391 295340 1400
rect 293592 1362 293644 1368
rect 117136 1148 117188 1154
rect 117136 1090 117188 1096
rect 193692 1057 193720 1362
rect 243740 1057 243768 1362
rect 163778 1048 163834 1057
rect 163778 983 163834 992
rect 193678 1048 193734 1057
rect 193678 983 193734 992
rect 229282 1048 229338 1057
rect 229282 983 229338 992
rect 243726 1048 243782 1057
rect 243726 983 243782 992
rect 114192 808 114244 814
rect 22652 750 22704 756
rect 32770 -400 32826 800
rect 98274 -400 98330 800
rect 163792 800 163820 983
rect 229296 800 229324 983
rect 294800 800 294828 1391
rect 295392 1391 295394 1400
rect 295340 1362 295392 1368
rect 360290 1048 360346 1057
rect 360290 983 360346 992
rect 360304 800 360332 983
rect 425808 800 425836 1430
rect 491312 800 491340 1430
rect 493612 1426 493640 2094
rect 493600 1420 493652 1426
rect 493600 1362 493652 1368
rect 114192 750 114244 756
rect 163778 -400 163834 800
rect 229282 -400 229338 800
rect 294786 -400 294842 800
rect 360290 -400 360346 800
rect 425794 -400 425850 800
rect 491298 -400 491354 800
rect 521120 785 521148 2751
rect 521106 776 521162 785
rect 521106 711 521162 720
<< via2 >>
rect 5354 155216 5410 155272
rect 7930 156576 7986 156632
rect 7102 153720 7158 153776
rect 12162 157936 12218 157992
rect 10414 153856 10470 153912
rect 19706 159296 19762 159352
rect 21362 156712 21418 156768
rect 27250 155352 27306 155408
rect 16302 152496 16358 152552
rect 9586 152360 9642 152416
rect 12990 152088 13046 152144
rect 9494 151952 9550 152008
rect 2686 151816 2742 151872
rect 2042 151000 2098 151056
rect 33138 159432 33194 159488
rect 30654 155488 30710 155544
rect 35714 158072 35770 158128
rect 38474 153992 38530 154048
rect 28906 151136 28962 151192
rect 30194 150456 30250 150512
rect 44086 151272 44142 151328
rect 55770 152768 55826 152824
rect 37002 150592 37058 150648
rect 60094 159568 60150 159624
rect 74354 160656 74410 160712
rect 71686 151408 71742 151464
rect 79414 158208 79470 158264
rect 82818 156848 82874 156904
rect 84106 152632 84162 152688
rect 87786 160792 87842 160848
rect 85486 151544 85542 151600
rect 6366 149368 6422 149424
rect 16486 149368 16542 149424
rect 20166 149368 20222 149424
rect 116306 152088 116362 152144
rect 113822 151952 113878 152008
rect 113730 144200 113786 144256
rect 113546 110064 113602 110120
rect 114282 150592 114338 150648
rect 113914 149096 113970 149152
rect 114098 150456 114154 150512
rect 114006 132776 114062 132832
rect 114190 121352 114246 121408
rect 120170 155624 120226 155680
rect 116122 148996 116124 149016
rect 116124 148996 116176 149016
rect 116176 148996 116178 149016
rect 116122 148960 116178 148996
rect 116030 147056 116086 147112
rect 116122 145152 116178 145208
rect 114466 98640 114522 98696
rect 115938 143248 115994 143304
rect 115938 141344 115994 141400
rect 115938 139440 115994 139496
rect 116122 131688 116178 131744
rect 115938 129784 115994 129840
rect 116122 125976 116178 126032
rect 116122 124108 116124 124128
rect 116124 124108 116176 124128
rect 116176 124108 116178 124128
rect 116122 124072 116178 124108
rect 115938 122168 115994 122224
rect 115938 120128 115994 120184
rect 114466 87236 114522 87272
rect 114466 87216 114468 87236
rect 114468 87216 114520 87236
rect 114520 87216 114522 87236
rect 116398 137536 116454 137592
rect 116582 149232 116638 149288
rect 116490 133592 116546 133648
rect 116214 118224 116270 118280
rect 116030 116320 116086 116376
rect 116122 114452 116124 114472
rect 116124 114452 116176 114472
rect 116176 114452 116178 114472
rect 116122 114416 116178 114452
rect 116122 112512 116178 112568
rect 116122 110608 116178 110664
rect 115294 83680 115350 83736
rect 116398 108704 116454 108760
rect 115938 104796 115940 104816
rect 115940 104796 115992 104816
rect 115992 104796 115994 104816
rect 115938 104760 115994 104796
rect 116582 97144 116638 97200
rect 118974 151000 119030 151056
rect 116766 149368 116822 149424
rect 123022 155216 123078 155272
rect 124770 156576 124826 156632
rect 124310 153720 124366 153776
rect 125506 153720 125562 153776
rect 127622 159296 127678 159352
rect 127070 157936 127126 157992
rect 126886 153856 126942 153912
rect 126334 152360 126390 152416
rect 131394 152496 131450 152552
rect 133418 159568 133474 159624
rect 135258 156712 135314 156768
rect 137466 159568 137522 159624
rect 138018 159432 138074 159488
rect 142342 155488 142398 155544
rect 139766 155352 139822 155408
rect 141698 152768 141754 152824
rect 141054 151136 141110 151192
rect 142526 155216 142582 155272
rect 145102 158072 145158 158128
rect 148138 153992 148194 154048
rect 152554 151272 152610 151328
rect 154210 155624 154266 155680
rect 156050 157936 156106 157992
rect 159362 159296 159418 159352
rect 162674 156576 162730 156632
rect 175462 160656 175518 160712
rect 173162 151408 173218 151464
rect 179418 157936 179474 157992
rect 179418 157800 179474 157856
rect 178682 153856 178738 153912
rect 179602 158208 179658 158264
rect 180982 156848 181038 156904
rect 182914 156712 182970 156768
rect 182730 152632 182786 152688
rect 182362 152496 182418 152552
rect 183374 151544 183430 151600
rect 184846 158072 184902 158128
rect 185950 160792 186006 160848
rect 187698 152360 187754 152416
rect 189630 155352 189686 155408
rect 201314 159568 201370 159624
rect 203338 157936 203394 157992
rect 204718 159432 204774 159488
rect 207294 157936 207350 157992
rect 209962 158072 210018 158128
rect 209778 153720 209834 153776
rect 213550 152360 213606 152416
rect 222106 152360 222162 152416
rect 223486 153720 223542 153776
rect 227718 155216 227774 155272
rect 227902 155216 227958 155272
rect 235906 158072 235962 158128
rect 236734 152496 236790 152552
rect 237470 159296 237526 159352
rect 243082 156576 243138 156632
rect 247038 156576 247094 156632
rect 255318 153856 255374 153912
rect 255502 153856 255558 153912
rect 258538 156712 258594 156768
rect 263690 155352 263746 155408
rect 265070 159432 265126 159488
rect 263874 155352 263930 155408
rect 276018 157936 276074 157992
rect 277766 152360 277822 152416
rect 284850 153720 284906 153776
rect 287426 155216 287482 155272
rect 292578 156576 292634 156632
rect 298650 158072 298706 158128
rect 297730 153856 297786 153912
rect 302882 155352 302938 155408
rect 519542 161608 519598 161664
rect 117042 135496 117098 135552
rect 116950 106800 117006 106856
rect 519634 160112 519690 160168
rect 519542 147872 519598 147928
rect 520922 162968 520978 163024
rect 521566 158616 521622 158672
rect 521014 157120 521070 157176
rect 520922 149232 520978 149288
rect 520922 148008 520978 148064
rect 519634 146512 519690 146568
rect 519818 146512 519874 146568
rect 519542 144880 519598 144936
rect 520738 143384 520794 143440
rect 519818 134272 519874 134328
rect 519542 132912 519598 132968
rect 520830 141888 520886 141944
rect 520738 131416 520794 131472
rect 521290 155624 521346 155680
rect 521198 151000 521254 151056
rect 521106 149504 521162 149560
rect 521014 143792 521070 143848
rect 521474 153992 521530 154048
rect 521382 152496 521438 152552
rect 521290 142432 521346 142488
rect 521566 145152 521622 145208
rect 521474 141072 521530 141128
rect 521566 140392 521622 140448
rect 521382 139712 521438 139768
rect 521382 138896 521438 138952
rect 521198 138352 521254 138408
rect 521106 136992 521162 137048
rect 521290 135768 521346 135824
rect 520922 135632 520978 135688
rect 521198 134272 521254 134328
rect 521106 132776 521162 132832
rect 520922 131280 520978 131336
rect 520830 130056 520886 130112
rect 520830 128288 520886 128344
rect 117134 127880 117190 127936
rect 520738 126656 520794 126712
rect 521014 129784 521070 129840
rect 520922 120536 520978 120592
rect 521474 137400 521530 137456
rect 521382 127336 521438 127392
rect 521566 128696 521622 128752
rect 521474 125976 521530 126032
rect 521474 125160 521530 125216
rect 521290 124616 521346 124672
rect 521382 123664 521438 123720
rect 521198 123256 521254 123312
rect 521290 122168 521346 122224
rect 521106 121896 521162 121952
rect 521014 119176 521070 119232
rect 521198 119176 521254 119232
rect 520830 117816 520886 117872
rect 521014 117544 521070 117600
rect 520738 116456 520794 116512
rect 520922 116048 520978 116104
rect 520738 113056 520794 113112
rect 520278 105440 520334 105496
rect 117042 102856 117098 102912
rect 116858 100952 116914 101008
rect 116766 99048 116822 99104
rect 520830 111560 520886 111616
rect 520738 104080 520794 104136
rect 521106 114552 521162 114608
rect 521014 108160 521070 108216
rect 520922 106800 520978 106856
rect 521566 120672 521622 120728
rect 521474 115096 521530 115152
rect 521382 113736 521438 113792
rect 521290 112240 521346 112296
rect 521566 110880 521622 110936
rect 521566 110064 521622 110120
rect 521198 109520 521254 109576
rect 521198 108432 521254 108488
rect 521106 105576 521162 105632
rect 521106 103944 521162 104000
rect 520830 102720 520886 102776
rect 521014 102448 521070 102504
rect 520922 100952 520978 101008
rect 520830 97824 520886 97880
rect 520278 97280 520334 97336
rect 116674 95240 116730 95296
rect 116490 93336 116546 93392
rect 116122 91296 116178 91352
rect 116214 85584 116270 85640
rect 115386 81776 115442 81832
rect 520370 96328 520426 96384
rect 520278 94832 520334 94888
rect 520738 93336 520794 93392
rect 520370 88984 520426 89040
rect 520278 87624 520334 87680
rect 116858 87488 116914 87544
rect 521382 106936 521438 106992
rect 521198 100000 521254 100056
rect 521198 99320 521254 99376
rect 521106 95920 521162 95976
rect 521014 94424 521070 94480
rect 520922 93064 520978 93120
rect 521014 91840 521070 91896
rect 520830 90344 520886 90400
rect 520738 86264 520794 86320
rect 520370 85720 520426 85776
rect 520278 84224 520334 84280
rect 116766 79872 116822 79928
rect 521566 101360 521622 101416
rect 521382 98640 521438 98696
rect 521198 91704 521254 91760
rect 521198 90208 521254 90264
rect 521106 87216 521162 87272
rect 521014 84904 521070 84960
rect 520738 82728 520794 82784
rect 520370 79464 520426 79520
rect 520278 78104 520334 78160
rect 116674 77968 116730 78024
rect 521014 81096 521070 81152
rect 520738 76744 520794 76800
rect 520462 76608 520518 76664
rect 520278 75112 520334 75168
rect 116582 74024 116638 74080
rect 116398 72120 116454 72176
rect 5998 1536 6054 1592
rect 15934 1808 15990 1864
rect 19338 1672 19394 1728
rect 29550 2080 29606 2136
rect 26054 1944 26110 2000
rect 42706 2216 42762 2272
rect 55954 1400 56010 1456
rect 97998 1264 98054 1320
rect 109958 1808 110014 1864
rect 111430 2080 111486 2136
rect 116306 70216 116362 70272
rect 113822 53080 113878 53136
rect 111614 1944 111670 2000
rect 100758 1128 100814 1184
rect 116214 68312 116270 68368
rect 114098 41792 114154 41848
rect 521290 88712 521346 88768
rect 521198 83544 521254 83600
rect 521290 82184 521346 82240
rect 521106 80824 521162 80880
rect 521382 79600 521438 79656
rect 521106 78104 521162 78160
rect 521014 75248 521070 75304
rect 520738 73616 520794 73672
rect 520462 71168 520518 71224
rect 520278 69808 520334 69864
rect 521382 73888 521438 73944
rect 521106 72528 521162 72584
rect 521014 71984 521070 72040
rect 520738 68448 520794 68504
rect 520462 67496 520518 67552
rect 116858 66408 116914 66464
rect 114466 64504 114522 64560
rect 115202 64504 115258 64560
rect 114190 30368 114246 30424
rect 114282 18944 114338 19000
rect 114190 7656 114246 7712
rect 116122 62600 116178 62656
rect 116122 60560 116178 60616
rect 116582 54848 116638 54904
rect 115938 51076 115940 51096
rect 115940 51076 115992 51096
rect 115992 51076 115994 51096
rect 115938 51040 115994 51076
rect 116030 47096 116086 47152
rect 116398 43288 116454 43344
rect 115938 39480 115994 39536
rect 116122 37576 116178 37632
rect 116122 33768 116178 33824
rect 116490 31728 116546 31784
rect 116122 27920 116178 27976
rect 116122 24112 116178 24168
rect 116398 29824 116454 29880
rect 116122 22208 116178 22264
rect 116122 20304 116178 20360
rect 116122 18400 116178 18456
rect 116122 16360 116178 16416
rect 115938 14456 115994 14512
rect 116030 4936 116086 4992
rect 116122 3032 116178 3088
rect 116030 1536 116086 1592
rect 116674 52944 116730 53000
rect 116766 49136 116822 49192
rect 520370 66000 520426 66056
rect 521106 70488 521162 70544
rect 521014 67088 521070 67144
rect 521290 68992 521346 69048
rect 521106 65728 521162 65784
rect 520738 64504 520794 64560
rect 520462 63008 520518 63064
rect 520370 61648 520426 61704
rect 521290 64368 521346 64424
rect 521106 62872 521162 62928
rect 521014 61376 521070 61432
rect 520738 60288 520794 60344
rect 520738 59880 520794 59936
rect 117042 58656 117098 58712
rect 116858 45192 116914 45248
rect 116950 41384 117006 41440
rect 520370 56888 520426 56944
rect 117134 56752 117190 56808
rect 520278 55392 520334 55448
rect 117134 35672 117190 35728
rect 117042 12552 117098 12608
rect 117042 1672 117098 1728
rect 521106 58928 521162 58984
rect 521106 58384 521162 58440
rect 521014 57432 521070 57488
rect 520738 56072 520794 56128
rect 521106 54712 521162 54768
rect 521106 53760 521162 53816
rect 520370 53352 520426 53408
rect 520922 52264 520978 52320
rect 520278 51992 520334 52048
rect 520370 50768 520426 50824
rect 521106 50632 521162 50688
rect 520922 49272 520978 49328
rect 521106 49272 521162 49328
rect 520370 47912 520426 47968
rect 520278 47776 520334 47832
rect 521106 46552 521162 46608
rect 520370 46280 520426 46336
rect 520278 45192 520334 45248
rect 521014 44648 521070 44704
rect 520370 43832 520426 43888
rect 521106 43152 521162 43208
rect 521014 42472 521070 42528
rect 521014 41656 521070 41712
rect 521106 41112 521162 41168
rect 521106 40160 521162 40216
rect 521014 39752 521070 39808
rect 520922 38664 520978 38720
rect 521106 38256 521162 38312
rect 521106 37168 521162 37224
rect 520922 36896 520978 36952
rect 521106 35944 521162 36000
rect 520922 35536 520978 35592
rect 520922 34584 520978 34640
rect 520830 34040 520886 34096
rect 520830 33224 520886 33280
rect 521106 32544 521162 32600
rect 521106 31728 521162 31784
rect 521106 31048 521162 31104
rect 521106 30368 521162 30424
rect 521106 29552 521162 29608
rect 521106 28736 521162 28792
rect 521106 20440 521162 20496
rect 521106 19760 521162 19816
rect 521106 15000 521162 15056
rect 521106 14320 521162 14376
rect 521106 13640 521162 13696
rect 521106 12824 521162 12880
rect 519634 12280 519690 12336
rect 519634 11328 519690 11384
rect 521106 10920 521162 10976
rect 117226 10648 117282 10704
rect 521106 9832 521162 9888
rect 521106 9560 521162 9616
rect 520370 8200 520426 8256
rect 521106 8200 521162 8256
rect 521106 6840 521162 6896
rect 520370 6704 520426 6760
rect 521014 5480 521070 5536
rect 520922 4120 520978 4176
rect 521106 5208 521162 5264
rect 521014 3712 521070 3768
rect 521106 2760 521162 2816
rect 520922 2216 520978 2272
rect 343960 1808 344016 1864
rect 294786 1400 294842 1456
rect 295338 1420 295394 1456
rect 295338 1400 295340 1420
rect 295340 1400 295392 1420
rect 295392 1400 295394 1420
rect 163778 992 163834 1048
rect 193678 992 193734 1048
rect 229282 992 229338 1048
rect 243726 992 243782 1048
rect 360290 992 360346 1048
rect 521106 720 521162 776
<< metal3 >>
rect 523200 163162 524400 163192
rect 520966 163102 524400 163162
rect 520966 163029 521026 163102
rect 523200 163072 524400 163102
rect 520917 163024 521026 163029
rect 520917 162968 520922 163024
rect 520978 162968 521026 163024
rect 520917 162966 521026 162968
rect 520917 162963 520983 162966
rect 519537 161666 519603 161669
rect 523200 161666 524400 161696
rect 519537 161664 524400 161666
rect 519537 161608 519542 161664
rect 519598 161608 524400 161664
rect 519537 161606 524400 161608
rect 519537 161603 519603 161606
rect 523200 161576 524400 161606
rect 87781 160850 87847 160853
rect 185945 160850 186011 160853
rect 87781 160848 186011 160850
rect 87781 160792 87786 160848
rect 87842 160792 185950 160848
rect 186006 160792 186011 160848
rect 87781 160790 186011 160792
rect 87781 160787 87847 160790
rect 185945 160787 186011 160790
rect 74349 160714 74415 160717
rect 175457 160714 175523 160717
rect 74349 160712 175523 160714
rect 74349 160656 74354 160712
rect 74410 160656 175462 160712
rect 175518 160656 175523 160712
rect 74349 160654 175523 160656
rect 74349 160651 74415 160654
rect 175457 160651 175523 160654
rect 519629 160170 519695 160173
rect 523200 160170 524400 160200
rect 519629 160168 524400 160170
rect 519629 160112 519634 160168
rect 519690 160112 524400 160168
rect 519629 160110 524400 160112
rect 519629 160107 519695 160110
rect 523200 160080 524400 160110
rect 60089 159626 60155 159629
rect 133413 159626 133479 159629
rect 60089 159624 133479 159626
rect 60089 159568 60094 159624
rect 60150 159568 133418 159624
rect 133474 159568 133479 159624
rect 60089 159566 133479 159568
rect 60089 159563 60155 159566
rect 133413 159563 133479 159566
rect 137461 159626 137527 159629
rect 201309 159626 201375 159629
rect 137461 159624 201375 159626
rect 137461 159568 137466 159624
rect 137522 159568 201314 159624
rect 201370 159568 201375 159624
rect 137461 159566 201375 159568
rect 137461 159563 137527 159566
rect 201309 159563 201375 159566
rect 33133 159490 33199 159493
rect 138013 159490 138079 159493
rect 33133 159488 138079 159490
rect 33133 159432 33138 159488
rect 33194 159432 138018 159488
rect 138074 159432 138079 159488
rect 33133 159430 138079 159432
rect 33133 159427 33199 159430
rect 138013 159427 138079 159430
rect 204713 159490 204779 159493
rect 265065 159490 265131 159493
rect 204713 159488 265131 159490
rect 204713 159432 204718 159488
rect 204774 159432 265070 159488
rect 265126 159432 265131 159488
rect 204713 159430 265131 159432
rect 204713 159427 204779 159430
rect 265065 159427 265131 159430
rect 19701 159354 19767 159357
rect 127617 159354 127683 159357
rect 19701 159352 127683 159354
rect 19701 159296 19706 159352
rect 19762 159296 127622 159352
rect 127678 159296 127683 159352
rect 19701 159294 127683 159296
rect 19701 159291 19767 159294
rect 127617 159291 127683 159294
rect 159357 159354 159423 159357
rect 237465 159354 237531 159357
rect 159357 159352 237531 159354
rect 159357 159296 159362 159352
rect 159418 159296 237470 159352
rect 237526 159296 237531 159352
rect 159357 159294 237531 159296
rect 159357 159291 159423 159294
rect 237465 159291 237531 159294
rect 521561 158674 521627 158677
rect 523200 158674 524400 158704
rect 521561 158672 524400 158674
rect 521561 158616 521566 158672
rect 521622 158616 524400 158672
rect 521561 158614 524400 158616
rect 521561 158611 521627 158614
rect 523200 158584 524400 158614
rect 79409 158266 79475 158269
rect 179597 158266 179663 158269
rect 79409 158264 179663 158266
rect 79409 158208 79414 158264
rect 79470 158208 179602 158264
rect 179658 158208 179663 158264
rect 79409 158206 179663 158208
rect 79409 158203 79475 158206
rect 179597 158203 179663 158206
rect 35709 158130 35775 158133
rect 145097 158130 145163 158133
rect 35709 158128 145163 158130
rect 35709 158072 35714 158128
rect 35770 158072 145102 158128
rect 145158 158072 145163 158128
rect 35709 158070 145163 158072
rect 35709 158067 35775 158070
rect 145097 158067 145163 158070
rect 184841 158130 184907 158133
rect 209957 158130 210023 158133
rect 184841 158128 210023 158130
rect 184841 158072 184846 158128
rect 184902 158072 209962 158128
rect 210018 158072 210023 158128
rect 184841 158070 210023 158072
rect 184841 158067 184907 158070
rect 209957 158067 210023 158070
rect 235901 158130 235967 158133
rect 298645 158130 298711 158133
rect 235901 158128 298711 158130
rect 235901 158072 235906 158128
rect 235962 158072 298650 158128
rect 298706 158072 298711 158128
rect 235901 158070 298711 158072
rect 235901 158067 235967 158070
rect 298645 158067 298711 158070
rect 12157 157994 12223 157997
rect 127065 157994 127131 157997
rect 12157 157992 127131 157994
rect 12157 157936 12162 157992
rect 12218 157936 127070 157992
rect 127126 157936 127131 157992
rect 12157 157934 127131 157936
rect 12157 157931 12223 157934
rect 127065 157931 127131 157934
rect 156045 157994 156111 157997
rect 179413 157994 179479 157997
rect 203333 157994 203399 157997
rect 156045 157992 161490 157994
rect 156045 157936 156050 157992
rect 156106 157936 161490 157992
rect 156045 157934 161490 157936
rect 156045 157931 156111 157934
rect 161430 157858 161490 157934
rect 179413 157992 203399 157994
rect 179413 157936 179418 157992
rect 179474 157936 203338 157992
rect 203394 157936 203399 157992
rect 179413 157934 203399 157936
rect 179413 157931 179479 157934
rect 203333 157931 203399 157934
rect 207289 157994 207355 157997
rect 276013 157994 276079 157997
rect 207289 157992 276079 157994
rect 207289 157936 207294 157992
rect 207350 157936 276018 157992
rect 276074 157936 276079 157992
rect 207289 157934 276079 157936
rect 207289 157931 207355 157934
rect 276013 157931 276079 157934
rect 179413 157858 179479 157861
rect 161430 157856 179479 157858
rect 161430 157800 179418 157856
rect 179474 157800 179479 157856
rect 161430 157798 179479 157800
rect 179413 157795 179479 157798
rect 521009 157178 521075 157181
rect 523200 157178 524400 157208
rect 521009 157176 524400 157178
rect 521009 157120 521014 157176
rect 521070 157120 524400 157176
rect 521009 157118 524400 157120
rect 521009 157115 521075 157118
rect 523200 157088 524400 157118
rect 82813 156906 82879 156909
rect 180977 156906 181043 156909
rect 82813 156904 181043 156906
rect 82813 156848 82818 156904
rect 82874 156848 180982 156904
rect 181038 156848 181043 156904
rect 82813 156846 181043 156848
rect 82813 156843 82879 156846
rect 180977 156843 181043 156846
rect 21357 156770 21423 156773
rect 135253 156770 135319 156773
rect 21357 156768 135319 156770
rect 21357 156712 21362 156768
rect 21418 156712 135258 156768
rect 135314 156712 135319 156768
rect 21357 156710 135319 156712
rect 21357 156707 21423 156710
rect 135253 156707 135319 156710
rect 182909 156770 182975 156773
rect 258533 156770 258599 156773
rect 182909 156768 258599 156770
rect 182909 156712 182914 156768
rect 182970 156712 258538 156768
rect 258594 156712 258599 156768
rect 182909 156710 258599 156712
rect 182909 156707 182975 156710
rect 258533 156707 258599 156710
rect 7925 156634 7991 156637
rect 124765 156634 124831 156637
rect 7925 156632 124831 156634
rect 7925 156576 7930 156632
rect 7986 156576 124770 156632
rect 124826 156576 124831 156632
rect 7925 156574 124831 156576
rect 7925 156571 7991 156574
rect 124765 156571 124831 156574
rect 162669 156634 162735 156637
rect 243077 156634 243143 156637
rect 162669 156632 243143 156634
rect 162669 156576 162674 156632
rect 162730 156576 243082 156632
rect 243138 156576 243143 156632
rect 162669 156574 243143 156576
rect 162669 156571 162735 156574
rect 243077 156571 243143 156574
rect 247033 156634 247099 156637
rect 292573 156634 292639 156637
rect 247033 156632 292639 156634
rect 247033 156576 247038 156632
rect 247094 156576 292578 156632
rect 292634 156576 292639 156632
rect 247033 156574 292639 156576
rect 247033 156571 247099 156574
rect 292573 156571 292639 156574
rect 120165 155682 120231 155685
rect 154205 155682 154271 155685
rect 120165 155680 154271 155682
rect 120165 155624 120170 155680
rect 120226 155624 154210 155680
rect 154266 155624 154271 155680
rect 120165 155622 154271 155624
rect 120165 155619 120231 155622
rect 154205 155619 154271 155622
rect 521285 155682 521351 155685
rect 523200 155682 524400 155712
rect 521285 155680 524400 155682
rect 521285 155624 521290 155680
rect 521346 155624 524400 155680
rect 521285 155622 524400 155624
rect 521285 155619 521351 155622
rect 523200 155592 524400 155622
rect 30649 155546 30715 155549
rect 142337 155546 142403 155549
rect 30649 155544 142403 155546
rect 30649 155488 30654 155544
rect 30710 155488 142342 155544
rect 142398 155488 142403 155544
rect 30649 155486 142403 155488
rect 30649 155483 30715 155486
rect 142337 155483 142403 155486
rect 27245 155410 27311 155413
rect 139761 155410 139827 155413
rect 27245 155408 139827 155410
rect 27245 155352 27250 155408
rect 27306 155352 139766 155408
rect 139822 155352 139827 155408
rect 27245 155350 139827 155352
rect 27245 155347 27311 155350
rect 139761 155347 139827 155350
rect 189625 155410 189691 155413
rect 263685 155410 263751 155413
rect 189625 155408 263751 155410
rect 189625 155352 189630 155408
rect 189686 155352 263690 155408
rect 263746 155352 263751 155408
rect 189625 155350 263751 155352
rect 189625 155347 189691 155350
rect 263685 155347 263751 155350
rect 263869 155410 263935 155413
rect 302877 155410 302943 155413
rect 263869 155408 302943 155410
rect 263869 155352 263874 155408
rect 263930 155352 302882 155408
rect 302938 155352 302943 155408
rect 263869 155350 302943 155352
rect 263869 155347 263935 155350
rect 302877 155347 302943 155350
rect 5349 155274 5415 155277
rect 123017 155274 123083 155277
rect 5349 155272 123083 155274
rect 5349 155216 5354 155272
rect 5410 155216 123022 155272
rect 123078 155216 123083 155272
rect 5349 155214 123083 155216
rect 5349 155211 5415 155214
rect 123017 155211 123083 155214
rect 142521 155274 142587 155277
rect 227713 155274 227779 155277
rect 142521 155272 227779 155274
rect 142521 155216 142526 155272
rect 142582 155216 227718 155272
rect 227774 155216 227779 155272
rect 142521 155214 227779 155216
rect 142521 155211 142587 155214
rect 227713 155211 227779 155214
rect 227897 155274 227963 155277
rect 287421 155274 287487 155277
rect 227897 155272 287487 155274
rect 227897 155216 227902 155272
rect 227958 155216 287426 155272
rect 287482 155216 287487 155272
rect 227897 155214 287487 155216
rect 227897 155211 227963 155214
rect 287421 155211 287487 155214
rect 38469 154050 38535 154053
rect 148133 154050 148199 154053
rect 38469 154048 148199 154050
rect 38469 153992 38474 154048
rect 38530 153992 148138 154048
rect 148194 153992 148199 154048
rect 38469 153990 148199 153992
rect 38469 153987 38535 153990
rect 148133 153987 148199 153990
rect 521469 154050 521535 154053
rect 523200 154050 524400 154080
rect 521469 154048 524400 154050
rect 521469 153992 521474 154048
rect 521530 153992 524400 154048
rect 521469 153990 524400 153992
rect 521469 153987 521535 153990
rect 523200 153960 524400 153990
rect 10409 153914 10475 153917
rect 126881 153914 126947 153917
rect 10409 153912 126947 153914
rect 10409 153856 10414 153912
rect 10470 153856 126886 153912
rect 126942 153856 126947 153912
rect 10409 153854 126947 153856
rect 10409 153851 10475 153854
rect 126881 153851 126947 153854
rect 178677 153914 178743 153917
rect 255313 153914 255379 153917
rect 178677 153912 255379 153914
rect 178677 153856 178682 153912
rect 178738 153856 255318 153912
rect 255374 153856 255379 153912
rect 178677 153854 255379 153856
rect 178677 153851 178743 153854
rect 255313 153851 255379 153854
rect 255497 153914 255563 153917
rect 297725 153914 297791 153917
rect 255497 153912 297791 153914
rect 255497 153856 255502 153912
rect 255558 153856 297730 153912
rect 297786 153856 297791 153912
rect 255497 153854 297791 153856
rect 255497 153851 255563 153854
rect 297725 153851 297791 153854
rect 7097 153778 7163 153781
rect 124305 153778 124371 153781
rect 7097 153776 124371 153778
rect 7097 153720 7102 153776
rect 7158 153720 124310 153776
rect 124366 153720 124371 153776
rect 7097 153718 124371 153720
rect 7097 153715 7163 153718
rect 124305 153715 124371 153718
rect 125501 153778 125567 153781
rect 209773 153778 209839 153781
rect 125501 153776 209839 153778
rect 125501 153720 125506 153776
rect 125562 153720 209778 153776
rect 209834 153720 209839 153776
rect 125501 153718 209839 153720
rect 125501 153715 125567 153718
rect 209773 153715 209839 153718
rect 223481 153778 223547 153781
rect 284845 153778 284911 153781
rect 223481 153776 284911 153778
rect 223481 153720 223486 153776
rect 223542 153720 284850 153776
rect 284906 153720 284911 153776
rect 223481 153718 284911 153720
rect 223481 153715 223547 153718
rect 284845 153715 284911 153718
rect 55765 152826 55831 152829
rect 141693 152826 141759 152829
rect 55765 152824 141759 152826
rect 55765 152768 55770 152824
rect 55826 152768 141698 152824
rect 141754 152768 141759 152824
rect 55765 152766 141759 152768
rect 55765 152763 55831 152766
rect 141693 152763 141759 152766
rect 84101 152690 84167 152693
rect 182725 152690 182791 152693
rect 84101 152688 182791 152690
rect 84101 152632 84106 152688
rect 84162 152632 182730 152688
rect 182786 152632 182791 152688
rect 84101 152630 182791 152632
rect 84101 152627 84167 152630
rect 182725 152627 182791 152630
rect 16297 152554 16363 152557
rect 131389 152554 131455 152557
rect 16297 152552 131455 152554
rect 16297 152496 16302 152552
rect 16358 152496 131394 152552
rect 131450 152496 131455 152552
rect 16297 152494 131455 152496
rect 16297 152491 16363 152494
rect 131389 152491 131455 152494
rect 182357 152554 182423 152557
rect 236729 152554 236795 152557
rect 182357 152552 236795 152554
rect 182357 152496 182362 152552
rect 182418 152496 236734 152552
rect 236790 152496 236795 152552
rect 182357 152494 236795 152496
rect 182357 152491 182423 152494
rect 236729 152491 236795 152494
rect 521377 152554 521443 152557
rect 523200 152554 524400 152584
rect 521377 152552 524400 152554
rect 521377 152496 521382 152552
rect 521438 152496 524400 152552
rect 521377 152494 524400 152496
rect 521377 152491 521443 152494
rect 523200 152464 524400 152494
rect 9581 152418 9647 152421
rect 126329 152418 126395 152421
rect 9581 152416 126395 152418
rect 9581 152360 9586 152416
rect 9642 152360 126334 152416
rect 126390 152360 126395 152416
rect 9581 152358 126395 152360
rect 9581 152355 9647 152358
rect 126329 152355 126395 152358
rect 187693 152418 187759 152421
rect 213545 152418 213611 152421
rect 187693 152416 213611 152418
rect 187693 152360 187698 152416
rect 187754 152360 213550 152416
rect 213606 152360 213611 152416
rect 187693 152358 213611 152360
rect 187693 152355 187759 152358
rect 213545 152355 213611 152358
rect 222101 152418 222167 152421
rect 277761 152418 277827 152421
rect 222101 152416 277827 152418
rect 222101 152360 222106 152416
rect 222162 152360 277766 152416
rect 277822 152360 277827 152416
rect 222101 152358 277827 152360
rect 222101 152355 222167 152358
rect 277761 152355 277827 152358
rect 12985 152146 13051 152149
rect 116301 152146 116367 152149
rect 12985 152144 116367 152146
rect 12985 152088 12990 152144
rect 13046 152088 116306 152144
rect 116362 152088 116367 152144
rect 12985 152086 116367 152088
rect 12985 152083 13051 152086
rect 116301 152083 116367 152086
rect 9489 152010 9555 152013
rect 113817 152010 113883 152013
rect 9489 152008 113883 152010
rect 9489 151952 9494 152008
rect 9550 151952 113822 152008
rect 113878 151952 113883 152008
rect 9489 151950 113883 151952
rect 9489 151947 9555 151950
rect 113817 151947 113883 151950
rect 2681 151874 2747 151877
rect 116526 151874 116532 151876
rect 2681 151872 116532 151874
rect 2681 151816 2686 151872
rect 2742 151816 116532 151872
rect 2681 151814 116532 151816
rect 2681 151811 2747 151814
rect 116526 151812 116532 151814
rect 116596 151812 116602 151876
rect 85481 151602 85547 151605
rect 183369 151602 183435 151605
rect 85481 151600 183435 151602
rect 85481 151544 85486 151600
rect 85542 151544 183374 151600
rect 183430 151544 183435 151600
rect 85481 151542 183435 151544
rect 85481 151539 85547 151542
rect 183369 151539 183435 151542
rect 71681 151466 71747 151469
rect 173157 151466 173223 151469
rect 71681 151464 173223 151466
rect 71681 151408 71686 151464
rect 71742 151408 173162 151464
rect 173218 151408 173223 151464
rect 71681 151406 173223 151408
rect 71681 151403 71747 151406
rect 173157 151403 173223 151406
rect 44081 151330 44147 151333
rect 152549 151330 152615 151333
rect 44081 151328 152615 151330
rect 44081 151272 44086 151328
rect 44142 151272 152554 151328
rect 152610 151272 152615 151328
rect 44081 151270 152615 151272
rect 44081 151267 44147 151270
rect 152549 151267 152615 151270
rect 28901 151194 28967 151197
rect 141049 151194 141115 151197
rect 28901 151192 141115 151194
rect 28901 151136 28906 151192
rect 28962 151136 141054 151192
rect 141110 151136 141115 151192
rect 28901 151134 141115 151136
rect 28901 151131 28967 151134
rect 141049 151131 141115 151134
rect 2037 151058 2103 151061
rect 118969 151058 119035 151061
rect 2037 151056 119035 151058
rect 2037 151000 2042 151056
rect 2098 151000 118974 151056
rect 119030 151000 119035 151056
rect 2037 150998 119035 151000
rect 2037 150995 2103 150998
rect 118969 150995 119035 150998
rect 521193 151058 521259 151061
rect 523200 151058 524400 151088
rect 521193 151056 524400 151058
rect 521193 151000 521198 151056
rect 521254 151000 524400 151056
rect 521193 150998 524400 151000
rect 521193 150995 521259 150998
rect 523200 150968 524400 150998
rect 36997 150650 37063 150653
rect 114277 150650 114343 150653
rect 36997 150648 114343 150650
rect 36997 150592 37002 150648
rect 37058 150592 114282 150648
rect 114338 150592 114343 150648
rect 36997 150590 114343 150592
rect 36997 150587 37063 150590
rect 114277 150587 114343 150590
rect 30189 150514 30255 150517
rect 114093 150514 114159 150517
rect 30189 150512 114159 150514
rect 30189 150456 30194 150512
rect 30250 150456 114098 150512
rect 114154 150456 114159 150512
rect 30189 150454 114159 150456
rect 30189 150451 30255 150454
rect 114093 150451 114159 150454
rect 521101 149562 521167 149565
rect 523200 149562 524400 149592
rect 521101 149560 524400 149562
rect 521101 149504 521106 149560
rect 521162 149504 524400 149560
rect 521101 149502 524400 149504
rect 521101 149499 521167 149502
rect 523200 149472 524400 149502
rect 6361 149426 6427 149429
rect 16481 149426 16547 149429
rect 20161 149426 20227 149429
rect 116761 149426 116827 149429
rect 6361 149424 6930 149426
rect 6361 149368 6366 149424
rect 6422 149368 6930 149424
rect 6361 149366 6930 149368
rect 6361 149363 6427 149366
rect 6870 149154 6930 149366
rect 16481 149424 16590 149426
rect 16481 149368 16486 149424
rect 16542 149368 16590 149424
rect 16481 149363 16590 149368
rect 20161 149424 116827 149426
rect 20161 149368 20166 149424
rect 20222 149368 116766 149424
rect 116822 149368 116827 149424
rect 20161 149366 116827 149368
rect 20161 149363 20227 149366
rect 116761 149363 116827 149366
rect 16530 149290 16590 149363
rect 116577 149290 116643 149293
rect 520917 149290 520983 149293
rect 16530 149288 116643 149290
rect 16530 149232 116582 149288
rect 116638 149232 116643 149288
rect 16530 149230 116643 149232
rect 518788 149288 520983 149290
rect 518788 149232 520922 149288
rect 520978 149232 520983 149288
rect 518788 149230 520983 149232
rect 116577 149227 116643 149230
rect 520917 149227 520983 149230
rect 113909 149154 113975 149157
rect 6870 149152 113975 149154
rect 6870 149096 113914 149152
rect 113970 149096 113975 149152
rect 6870 149094 113975 149096
rect 113909 149091 113975 149094
rect 116117 149018 116183 149021
rect 116117 149016 119140 149018
rect 116117 148960 116122 149016
rect 116178 148960 119140 149016
rect 116117 148958 119140 148960
rect 116117 148955 116183 148958
rect 520917 148066 520983 148069
rect 523200 148066 524400 148096
rect 520917 148064 524400 148066
rect 520917 148008 520922 148064
rect 520978 148008 524400 148064
rect 520917 148006 524400 148008
rect 520917 148003 520983 148006
rect 523200 147976 524400 148006
rect 519537 147930 519603 147933
rect 518788 147928 519603 147930
rect 518788 147872 519542 147928
rect 519598 147872 519603 147928
rect 518788 147870 519603 147872
rect 519537 147867 519603 147870
rect 116025 147114 116091 147117
rect 116025 147112 119140 147114
rect 116025 147056 116030 147112
rect 116086 147056 119140 147112
rect 116025 147054 119140 147056
rect 116025 147051 116091 147054
rect 519629 146570 519695 146573
rect 518788 146568 519695 146570
rect 518788 146512 519634 146568
rect 519690 146512 519695 146568
rect 518788 146510 519695 146512
rect 519629 146507 519695 146510
rect 519813 146570 519879 146573
rect 523200 146570 524400 146600
rect 519813 146568 524400 146570
rect 519813 146512 519818 146568
rect 519874 146512 524400 146568
rect 519813 146510 524400 146512
rect 519813 146507 519879 146510
rect 523200 146480 524400 146510
rect 116117 145210 116183 145213
rect 521561 145210 521627 145213
rect 116117 145208 119140 145210
rect 116117 145152 116122 145208
rect 116178 145152 119140 145208
rect 116117 145150 119140 145152
rect 518788 145208 521627 145210
rect 518788 145152 521566 145208
rect 521622 145152 521627 145208
rect 518788 145150 521627 145152
rect 116117 145147 116183 145150
rect 521561 145147 521627 145150
rect 519537 144938 519603 144941
rect 523200 144938 524400 144968
rect 519537 144936 524400 144938
rect 519537 144880 519542 144936
rect 519598 144880 524400 144936
rect 519537 144878 524400 144880
rect 519537 144875 519603 144878
rect 523200 144848 524400 144878
rect 113725 144258 113791 144261
rect 110860 144256 113791 144258
rect 110860 144200 113730 144256
rect 113786 144200 113791 144256
rect 110860 144198 113791 144200
rect 113725 144195 113791 144198
rect 521009 143850 521075 143853
rect 518788 143848 521075 143850
rect 518788 143792 521014 143848
rect 521070 143792 521075 143848
rect 518788 143790 521075 143792
rect 521009 143787 521075 143790
rect 520733 143442 520799 143445
rect 523200 143442 524400 143472
rect 520733 143440 524400 143442
rect 520733 143384 520738 143440
rect 520794 143384 524400 143440
rect 520733 143382 524400 143384
rect 520733 143379 520799 143382
rect 523200 143352 524400 143382
rect 115933 143306 115999 143309
rect 115933 143304 119140 143306
rect 115933 143248 115938 143304
rect 115994 143248 119140 143304
rect 115933 143246 119140 143248
rect 115933 143243 115999 143246
rect 521285 142490 521351 142493
rect 518788 142488 521351 142490
rect 518788 142432 521290 142488
rect 521346 142432 521351 142488
rect 518788 142430 521351 142432
rect 521285 142427 521351 142430
rect 520825 141946 520891 141949
rect 523200 141946 524400 141976
rect 520825 141944 524400 141946
rect 520825 141888 520830 141944
rect 520886 141888 524400 141944
rect 520825 141886 524400 141888
rect 520825 141883 520891 141886
rect 523200 141856 524400 141886
rect 115933 141402 115999 141405
rect 115933 141400 119140 141402
rect 115933 141344 115938 141400
rect 115994 141344 119140 141400
rect 115933 141342 119140 141344
rect 115933 141339 115999 141342
rect 521469 141130 521535 141133
rect 518788 141128 521535 141130
rect 518788 141072 521474 141128
rect 521530 141072 521535 141128
rect 518788 141070 521535 141072
rect 521469 141067 521535 141070
rect 521561 140450 521627 140453
rect 523200 140450 524400 140480
rect 521561 140448 524400 140450
rect 521561 140392 521566 140448
rect 521622 140392 524400 140448
rect 521561 140390 524400 140392
rect 521561 140387 521627 140390
rect 523200 140360 524400 140390
rect 521377 139770 521443 139773
rect 518788 139768 521443 139770
rect 518788 139712 521382 139768
rect 521438 139712 521443 139768
rect 518788 139710 521443 139712
rect 521377 139707 521443 139710
rect 115933 139498 115999 139501
rect 115933 139496 119140 139498
rect 115933 139440 115938 139496
rect 115994 139440 119140 139496
rect 115933 139438 119140 139440
rect 115933 139435 115999 139438
rect 521377 138954 521443 138957
rect 523200 138954 524400 138984
rect 521377 138952 524400 138954
rect 521377 138896 521382 138952
rect 521438 138896 524400 138952
rect 521377 138894 524400 138896
rect 521377 138891 521443 138894
rect 523200 138864 524400 138894
rect 521193 138410 521259 138413
rect 518788 138408 521259 138410
rect 518788 138352 521198 138408
rect 521254 138352 521259 138408
rect 518788 138350 521259 138352
rect 521193 138347 521259 138350
rect 116393 137594 116459 137597
rect 116393 137592 119140 137594
rect 116393 137536 116398 137592
rect 116454 137536 119140 137592
rect 116393 137534 119140 137536
rect 116393 137531 116459 137534
rect 521469 137458 521535 137461
rect 523200 137458 524400 137488
rect 521469 137456 524400 137458
rect 521469 137400 521474 137456
rect 521530 137400 524400 137456
rect 521469 137398 524400 137400
rect 521469 137395 521535 137398
rect 523200 137368 524400 137398
rect 521101 137050 521167 137053
rect 518788 137048 521167 137050
rect 518788 136992 521106 137048
rect 521162 136992 521167 137048
rect 518788 136990 521167 136992
rect 521101 136987 521167 136990
rect 521285 135826 521351 135829
rect 523200 135826 524400 135856
rect 521285 135824 524400 135826
rect 521285 135768 521290 135824
rect 521346 135768 524400 135824
rect 521285 135766 524400 135768
rect 521285 135763 521351 135766
rect 523200 135736 524400 135766
rect 520917 135690 520983 135693
rect 518788 135688 520983 135690
rect 518788 135632 520922 135688
rect 520978 135632 520983 135688
rect 518788 135630 520983 135632
rect 520917 135627 520983 135630
rect 117037 135554 117103 135557
rect 117037 135552 119140 135554
rect 117037 135496 117042 135552
rect 117098 135496 119140 135552
rect 117037 135494 119140 135496
rect 117037 135491 117103 135494
rect 519813 134330 519879 134333
rect 518788 134328 519879 134330
rect 518788 134272 519818 134328
rect 519874 134272 519879 134328
rect 518788 134270 519879 134272
rect 519813 134267 519879 134270
rect 521193 134330 521259 134333
rect 523200 134330 524400 134360
rect 521193 134328 524400 134330
rect 521193 134272 521198 134328
rect 521254 134272 524400 134328
rect 521193 134270 524400 134272
rect 521193 134267 521259 134270
rect 523200 134240 524400 134270
rect 116485 133650 116551 133653
rect 116485 133648 119140 133650
rect 116485 133592 116490 133648
rect 116546 133592 119140 133648
rect 116485 133590 119140 133592
rect 116485 133587 116551 133590
rect 519537 132970 519603 132973
rect 518788 132968 519603 132970
rect 518788 132912 519542 132968
rect 519598 132912 519603 132968
rect 518788 132910 519603 132912
rect 519537 132907 519603 132910
rect 114001 132834 114067 132837
rect 110860 132832 114067 132834
rect 110860 132776 114006 132832
rect 114062 132776 114067 132832
rect 110860 132774 114067 132776
rect 114001 132771 114067 132774
rect 521101 132834 521167 132837
rect 523200 132834 524400 132864
rect 521101 132832 524400 132834
rect 521101 132776 521106 132832
rect 521162 132776 524400 132832
rect 521101 132774 524400 132776
rect 521101 132771 521167 132774
rect 523200 132744 524400 132774
rect 116117 131746 116183 131749
rect 116117 131744 119140 131746
rect 116117 131688 116122 131744
rect 116178 131688 119140 131744
rect 116117 131686 119140 131688
rect 116117 131683 116183 131686
rect 520733 131474 520799 131477
rect 518788 131472 520799 131474
rect 518788 131416 520738 131472
rect 520794 131416 520799 131472
rect 518788 131414 520799 131416
rect 520733 131411 520799 131414
rect 520917 131338 520983 131341
rect 523200 131338 524400 131368
rect 520917 131336 524400 131338
rect 520917 131280 520922 131336
rect 520978 131280 524400 131336
rect 520917 131278 524400 131280
rect 520917 131275 520983 131278
rect 523200 131248 524400 131278
rect 520825 130114 520891 130117
rect 518788 130112 520891 130114
rect 518788 130056 520830 130112
rect 520886 130056 520891 130112
rect 518788 130054 520891 130056
rect 520825 130051 520891 130054
rect 115933 129842 115999 129845
rect 521009 129842 521075 129845
rect 523200 129842 524400 129872
rect 115933 129840 119140 129842
rect 115933 129784 115938 129840
rect 115994 129784 119140 129840
rect 115933 129782 119140 129784
rect 521009 129840 524400 129842
rect 521009 129784 521014 129840
rect 521070 129784 524400 129840
rect 521009 129782 524400 129784
rect 115933 129779 115999 129782
rect 521009 129779 521075 129782
rect 523200 129752 524400 129782
rect 521561 128754 521627 128757
rect 518788 128752 521627 128754
rect 518788 128696 521566 128752
rect 521622 128696 521627 128752
rect 518788 128694 521627 128696
rect 521561 128691 521627 128694
rect 520825 128346 520891 128349
rect 523200 128346 524400 128376
rect 520825 128344 524400 128346
rect 520825 128288 520830 128344
rect 520886 128288 524400 128344
rect 520825 128286 524400 128288
rect 520825 128283 520891 128286
rect 523200 128256 524400 128286
rect 117129 127938 117195 127941
rect 117129 127936 119140 127938
rect 117129 127880 117134 127936
rect 117190 127880 119140 127936
rect 117129 127878 119140 127880
rect 117129 127875 117195 127878
rect 521377 127394 521443 127397
rect 518788 127392 521443 127394
rect 518788 127336 521382 127392
rect 521438 127336 521443 127392
rect 518788 127334 521443 127336
rect 521377 127331 521443 127334
rect 520733 126714 520799 126717
rect 523200 126714 524400 126744
rect 520733 126712 524400 126714
rect 520733 126656 520738 126712
rect 520794 126656 524400 126712
rect 520733 126654 524400 126656
rect 520733 126651 520799 126654
rect 523200 126624 524400 126654
rect 116117 126034 116183 126037
rect 521469 126034 521535 126037
rect 116117 126032 119140 126034
rect 116117 125976 116122 126032
rect 116178 125976 119140 126032
rect 116117 125974 119140 125976
rect 518788 126032 521535 126034
rect 518788 125976 521474 126032
rect 521530 125976 521535 126032
rect 518788 125974 521535 125976
rect 116117 125971 116183 125974
rect 521469 125971 521535 125974
rect 521469 125218 521535 125221
rect 523200 125218 524400 125248
rect 521469 125216 524400 125218
rect 521469 125160 521474 125216
rect 521530 125160 524400 125216
rect 521469 125158 524400 125160
rect 521469 125155 521535 125158
rect 523200 125128 524400 125158
rect 521285 124674 521351 124677
rect 518788 124672 521351 124674
rect 518788 124616 521290 124672
rect 521346 124616 521351 124672
rect 518788 124614 521351 124616
rect 521285 124611 521351 124614
rect 116117 124130 116183 124133
rect 116117 124128 119140 124130
rect 116117 124072 116122 124128
rect 116178 124072 119140 124128
rect 116117 124070 119140 124072
rect 116117 124067 116183 124070
rect 521377 123722 521443 123725
rect 523200 123722 524400 123752
rect 521377 123720 524400 123722
rect 521377 123664 521382 123720
rect 521438 123664 524400 123720
rect 521377 123662 524400 123664
rect 521377 123659 521443 123662
rect 523200 123632 524400 123662
rect 521193 123314 521259 123317
rect 518788 123312 521259 123314
rect 518788 123256 521198 123312
rect 521254 123256 521259 123312
rect 518788 123254 521259 123256
rect 521193 123251 521259 123254
rect 115933 122226 115999 122229
rect 521285 122226 521351 122229
rect 523200 122226 524400 122256
rect 115933 122224 119140 122226
rect 115933 122168 115938 122224
rect 115994 122168 119140 122224
rect 115933 122166 119140 122168
rect 521285 122224 524400 122226
rect 521285 122168 521290 122224
rect 521346 122168 524400 122224
rect 521285 122166 524400 122168
rect 115933 122163 115999 122166
rect 521285 122163 521351 122166
rect 523200 122136 524400 122166
rect 521101 121954 521167 121957
rect 518788 121952 521167 121954
rect 518788 121896 521106 121952
rect 521162 121896 521167 121952
rect 518788 121894 521167 121896
rect 521101 121891 521167 121894
rect 114185 121410 114251 121413
rect 110860 121408 114251 121410
rect 110860 121352 114190 121408
rect 114246 121352 114251 121408
rect 110860 121350 114251 121352
rect 114185 121347 114251 121350
rect 521561 120730 521627 120733
rect 523200 120730 524400 120760
rect 521561 120728 524400 120730
rect 521561 120672 521566 120728
rect 521622 120672 524400 120728
rect 521561 120670 524400 120672
rect 521561 120667 521627 120670
rect 523200 120640 524400 120670
rect 520917 120594 520983 120597
rect 518788 120592 520983 120594
rect 518788 120536 520922 120592
rect 520978 120536 520983 120592
rect 518788 120534 520983 120536
rect 520917 120531 520983 120534
rect 115933 120186 115999 120189
rect 115933 120184 119140 120186
rect 115933 120128 115938 120184
rect 115994 120128 119140 120184
rect 115933 120126 119140 120128
rect 115933 120123 115999 120126
rect 521009 119234 521075 119237
rect 518788 119232 521075 119234
rect 518788 119176 521014 119232
rect 521070 119176 521075 119232
rect 518788 119174 521075 119176
rect 521009 119171 521075 119174
rect 521193 119234 521259 119237
rect 523200 119234 524400 119264
rect 521193 119232 524400 119234
rect 521193 119176 521198 119232
rect 521254 119176 524400 119232
rect 521193 119174 524400 119176
rect 521193 119171 521259 119174
rect 523200 119144 524400 119174
rect 116209 118282 116275 118285
rect 116209 118280 119140 118282
rect 116209 118224 116214 118280
rect 116270 118224 119140 118280
rect 116209 118222 119140 118224
rect 116209 118219 116275 118222
rect 520825 117874 520891 117877
rect 518788 117872 520891 117874
rect 518788 117816 520830 117872
rect 520886 117816 520891 117872
rect 518788 117814 520891 117816
rect 520825 117811 520891 117814
rect 521009 117602 521075 117605
rect 523200 117602 524400 117632
rect 521009 117600 524400 117602
rect 521009 117544 521014 117600
rect 521070 117544 524400 117600
rect 521009 117542 524400 117544
rect 521009 117539 521075 117542
rect 523200 117512 524400 117542
rect 520733 116514 520799 116517
rect 518788 116512 520799 116514
rect 518788 116456 520738 116512
rect 520794 116456 520799 116512
rect 518788 116454 520799 116456
rect 520733 116451 520799 116454
rect 116025 116378 116091 116381
rect 116025 116376 119140 116378
rect 116025 116320 116030 116376
rect 116086 116320 119140 116376
rect 116025 116318 119140 116320
rect 116025 116315 116091 116318
rect 520917 116106 520983 116109
rect 523200 116106 524400 116136
rect 520917 116104 524400 116106
rect 520917 116048 520922 116104
rect 520978 116048 524400 116104
rect 520917 116046 524400 116048
rect 520917 116043 520983 116046
rect 523200 116016 524400 116046
rect 521469 115154 521535 115157
rect 518788 115152 521535 115154
rect 518788 115096 521474 115152
rect 521530 115096 521535 115152
rect 518788 115094 521535 115096
rect 521469 115091 521535 115094
rect 521101 114610 521167 114613
rect 523200 114610 524400 114640
rect 521101 114608 524400 114610
rect 521101 114552 521106 114608
rect 521162 114552 524400 114608
rect 521101 114550 524400 114552
rect 521101 114547 521167 114550
rect 523200 114520 524400 114550
rect 116117 114474 116183 114477
rect 116117 114472 119140 114474
rect 116117 114416 116122 114472
rect 116178 114416 119140 114472
rect 116117 114414 119140 114416
rect 116117 114411 116183 114414
rect 521377 113794 521443 113797
rect 518788 113792 521443 113794
rect 518788 113736 521382 113792
rect 521438 113736 521443 113792
rect 518788 113734 521443 113736
rect 521377 113731 521443 113734
rect 520733 113114 520799 113117
rect 523200 113114 524400 113144
rect 520733 113112 524400 113114
rect 520733 113056 520738 113112
rect 520794 113056 524400 113112
rect 520733 113054 524400 113056
rect 520733 113051 520799 113054
rect 523200 113024 524400 113054
rect 116117 112570 116183 112573
rect 116117 112568 119140 112570
rect 116117 112512 116122 112568
rect 116178 112512 119140 112568
rect 116117 112510 119140 112512
rect 116117 112507 116183 112510
rect 521285 112298 521351 112301
rect 518788 112296 521351 112298
rect 518788 112240 521290 112296
rect 521346 112240 521351 112296
rect 518788 112238 521351 112240
rect 521285 112235 521351 112238
rect 520825 111618 520891 111621
rect 523200 111618 524400 111648
rect 520825 111616 524400 111618
rect 520825 111560 520830 111616
rect 520886 111560 524400 111616
rect 520825 111558 524400 111560
rect 520825 111555 520891 111558
rect 523200 111528 524400 111558
rect 521561 110938 521627 110941
rect 518788 110936 521627 110938
rect 518788 110880 521566 110936
rect 521622 110880 521627 110936
rect 518788 110878 521627 110880
rect 521561 110875 521627 110878
rect 116117 110666 116183 110669
rect 116117 110664 119140 110666
rect 116117 110608 116122 110664
rect 116178 110608 119140 110664
rect 116117 110606 119140 110608
rect 116117 110603 116183 110606
rect 113541 110122 113607 110125
rect 110860 110120 113607 110122
rect 110860 110064 113546 110120
rect 113602 110064 113607 110120
rect 110860 110062 113607 110064
rect 113541 110059 113607 110062
rect 521561 110122 521627 110125
rect 523200 110122 524400 110152
rect 521561 110120 524400 110122
rect 521561 110064 521566 110120
rect 521622 110064 524400 110120
rect 521561 110062 524400 110064
rect 521561 110059 521627 110062
rect 523200 110032 524400 110062
rect 521193 109578 521259 109581
rect 518788 109576 521259 109578
rect 518788 109520 521198 109576
rect 521254 109520 521259 109576
rect 518788 109518 521259 109520
rect 521193 109515 521259 109518
rect 116393 108762 116459 108765
rect 116393 108760 119140 108762
rect 116393 108704 116398 108760
rect 116454 108704 119140 108760
rect 116393 108702 119140 108704
rect 116393 108699 116459 108702
rect 521193 108490 521259 108493
rect 523200 108490 524400 108520
rect 521193 108488 524400 108490
rect 521193 108432 521198 108488
rect 521254 108432 524400 108488
rect 521193 108430 524400 108432
rect 521193 108427 521259 108430
rect 523200 108400 524400 108430
rect 521009 108218 521075 108221
rect 518788 108216 521075 108218
rect 518788 108160 521014 108216
rect 521070 108160 521075 108216
rect 518788 108158 521075 108160
rect 521009 108155 521075 108158
rect 521377 106994 521443 106997
rect 523200 106994 524400 107024
rect 521377 106992 524400 106994
rect 521377 106936 521382 106992
rect 521438 106936 524400 106992
rect 521377 106934 524400 106936
rect 521377 106931 521443 106934
rect 523200 106904 524400 106934
rect 116945 106858 117011 106861
rect 520917 106858 520983 106861
rect 116945 106856 119140 106858
rect 116945 106800 116950 106856
rect 117006 106800 119140 106856
rect 116945 106798 119140 106800
rect 518788 106856 520983 106858
rect 518788 106800 520922 106856
rect 520978 106800 520983 106856
rect 518788 106798 520983 106800
rect 116945 106795 117011 106798
rect 520917 106795 520983 106798
rect 521101 105634 521167 105637
rect 518758 105632 521167 105634
rect 518758 105576 521106 105632
rect 521162 105576 521167 105632
rect 518758 105574 521167 105576
rect 518758 105468 518818 105574
rect 521101 105571 521167 105574
rect 520273 105498 520339 105501
rect 523200 105498 524400 105528
rect 520273 105496 524400 105498
rect 520273 105440 520278 105496
rect 520334 105440 524400 105496
rect 520273 105438 524400 105440
rect 520273 105435 520339 105438
rect 523200 105408 524400 105438
rect 115933 104818 115999 104821
rect 115933 104816 119140 104818
rect 115933 104760 115938 104816
rect 115994 104760 119140 104816
rect 115933 104758 119140 104760
rect 115933 104755 115999 104758
rect 520733 104138 520799 104141
rect 518788 104136 520799 104138
rect 518788 104080 520738 104136
rect 520794 104080 520799 104136
rect 518788 104078 520799 104080
rect 520733 104075 520799 104078
rect 521101 104002 521167 104005
rect 523200 104002 524400 104032
rect 521101 104000 524400 104002
rect 521101 103944 521106 104000
rect 521162 103944 524400 104000
rect 521101 103942 524400 103944
rect 521101 103939 521167 103942
rect 523200 103912 524400 103942
rect 117037 102914 117103 102917
rect 117037 102912 119140 102914
rect 117037 102856 117042 102912
rect 117098 102856 119140 102912
rect 117037 102854 119140 102856
rect 117037 102851 117103 102854
rect 520825 102778 520891 102781
rect 518788 102776 520891 102778
rect 518788 102720 520830 102776
rect 520886 102720 520891 102776
rect 518788 102718 520891 102720
rect 520825 102715 520891 102718
rect 521009 102506 521075 102509
rect 523200 102506 524400 102536
rect 521009 102504 524400 102506
rect 521009 102448 521014 102504
rect 521070 102448 524400 102504
rect 521009 102446 524400 102448
rect 521009 102443 521075 102446
rect 523200 102416 524400 102446
rect 521561 101418 521627 101421
rect 518788 101416 521627 101418
rect 518788 101360 521566 101416
rect 521622 101360 521627 101416
rect 518788 101358 521627 101360
rect 521561 101355 521627 101358
rect 116853 101010 116919 101013
rect 520917 101010 520983 101013
rect 523200 101010 524400 101040
rect 116853 101008 119140 101010
rect 116853 100952 116858 101008
rect 116914 100952 119140 101008
rect 116853 100950 119140 100952
rect 520917 101008 524400 101010
rect 520917 100952 520922 101008
rect 520978 100952 524400 101008
rect 520917 100950 524400 100952
rect 116853 100947 116919 100950
rect 520917 100947 520983 100950
rect 523200 100920 524400 100950
rect 521193 100058 521259 100061
rect 518788 100056 521259 100058
rect 518788 100000 521198 100056
rect 521254 100000 521259 100056
rect 518788 99998 521259 100000
rect 521193 99995 521259 99998
rect 521193 99378 521259 99381
rect 523200 99378 524400 99408
rect 521193 99376 524400 99378
rect 521193 99320 521198 99376
rect 521254 99320 524400 99376
rect 521193 99318 524400 99320
rect 521193 99315 521259 99318
rect 523200 99288 524400 99318
rect 116761 99106 116827 99109
rect 116761 99104 119140 99106
rect 116761 99048 116766 99104
rect 116822 99048 119140 99104
rect 116761 99046 119140 99048
rect 116761 99043 116827 99046
rect 114461 98698 114527 98701
rect 521377 98698 521443 98701
rect 110860 98696 114527 98698
rect 110860 98640 114466 98696
rect 114522 98640 114527 98696
rect 110860 98638 114527 98640
rect 518788 98696 521443 98698
rect 518788 98640 521382 98696
rect 521438 98640 521443 98696
rect 518788 98638 521443 98640
rect 114461 98635 114527 98638
rect 521377 98635 521443 98638
rect 520825 97882 520891 97885
rect 523200 97882 524400 97912
rect 520825 97880 524400 97882
rect 520825 97824 520830 97880
rect 520886 97824 524400 97880
rect 520825 97822 524400 97824
rect 520825 97819 520891 97822
rect 523200 97792 524400 97822
rect 520273 97338 520339 97341
rect 518788 97336 520339 97338
rect 518788 97280 520278 97336
rect 520334 97280 520339 97336
rect 518788 97278 520339 97280
rect 520273 97275 520339 97278
rect 116577 97202 116643 97205
rect 116577 97200 119140 97202
rect 116577 97144 116582 97200
rect 116638 97144 119140 97200
rect 116577 97142 119140 97144
rect 116577 97139 116643 97142
rect 520365 96386 520431 96389
rect 523200 96386 524400 96416
rect 520365 96384 524400 96386
rect 520365 96328 520370 96384
rect 520426 96328 524400 96384
rect 520365 96326 524400 96328
rect 520365 96323 520431 96326
rect 523200 96296 524400 96326
rect 521101 95978 521167 95981
rect 518788 95976 521167 95978
rect 518788 95920 521106 95976
rect 521162 95920 521167 95976
rect 518788 95918 521167 95920
rect 521101 95915 521167 95918
rect 116669 95298 116735 95301
rect 116669 95296 119140 95298
rect 116669 95240 116674 95296
rect 116730 95240 119140 95296
rect 116669 95238 119140 95240
rect 116669 95235 116735 95238
rect 520273 94890 520339 94893
rect 523200 94890 524400 94920
rect 520273 94888 524400 94890
rect 520273 94832 520278 94888
rect 520334 94832 524400 94888
rect 520273 94830 524400 94832
rect 520273 94827 520339 94830
rect 523200 94800 524400 94830
rect 521009 94482 521075 94485
rect 518788 94480 521075 94482
rect 518788 94424 521014 94480
rect 521070 94424 521075 94480
rect 518788 94422 521075 94424
rect 521009 94419 521075 94422
rect 116485 93394 116551 93397
rect 520733 93394 520799 93397
rect 523200 93394 524400 93424
rect 116485 93392 119140 93394
rect 116485 93336 116490 93392
rect 116546 93336 119140 93392
rect 116485 93334 119140 93336
rect 520733 93392 524400 93394
rect 520733 93336 520738 93392
rect 520794 93336 524400 93392
rect 520733 93334 524400 93336
rect 116485 93331 116551 93334
rect 520733 93331 520799 93334
rect 523200 93304 524400 93334
rect 520917 93122 520983 93125
rect 518788 93120 520983 93122
rect 518788 93064 520922 93120
rect 520978 93064 520983 93120
rect 518788 93062 520983 93064
rect 520917 93059 520983 93062
rect 521009 91898 521075 91901
rect 523200 91898 524400 91928
rect 521009 91896 524400 91898
rect 521009 91840 521014 91896
rect 521070 91840 524400 91896
rect 521009 91838 524400 91840
rect 521009 91835 521075 91838
rect 523200 91808 524400 91838
rect 521193 91762 521259 91765
rect 518788 91760 521259 91762
rect 518788 91704 521198 91760
rect 521254 91704 521259 91760
rect 518788 91702 521259 91704
rect 521193 91699 521259 91702
rect 116117 91354 116183 91357
rect 116117 91352 119140 91354
rect 116117 91296 116122 91352
rect 116178 91296 119140 91352
rect 116117 91294 119140 91296
rect 116117 91291 116183 91294
rect 520825 90402 520891 90405
rect 518788 90400 520891 90402
rect 518788 90344 520830 90400
rect 520886 90344 520891 90400
rect 518788 90342 520891 90344
rect 520825 90339 520891 90342
rect 521193 90266 521259 90269
rect 523200 90266 524400 90296
rect 521193 90264 524400 90266
rect 521193 90208 521198 90264
rect 521254 90208 524400 90264
rect 521193 90206 524400 90208
rect 521193 90203 521259 90206
rect 523200 90176 524400 90206
rect 116526 89388 116532 89452
rect 116596 89450 116602 89452
rect 116596 89390 119140 89450
rect 116596 89388 116602 89390
rect 520365 89042 520431 89045
rect 518788 89040 520431 89042
rect 518788 88984 520370 89040
rect 520426 88984 520431 89040
rect 518788 88982 520431 88984
rect 520365 88979 520431 88982
rect 521285 88770 521351 88773
rect 523200 88770 524400 88800
rect 521285 88768 524400 88770
rect 521285 88712 521290 88768
rect 521346 88712 524400 88768
rect 521285 88710 524400 88712
rect 521285 88707 521351 88710
rect 523200 88680 524400 88710
rect 520273 87682 520339 87685
rect 518788 87680 520339 87682
rect 518788 87624 520278 87680
rect 520334 87624 520339 87680
rect 518788 87622 520339 87624
rect 520273 87619 520339 87622
rect 116853 87546 116919 87549
rect 116853 87544 119140 87546
rect 116853 87488 116858 87544
rect 116914 87488 119140 87544
rect 116853 87486 119140 87488
rect 116853 87483 116919 87486
rect 114461 87274 114527 87277
rect 110860 87272 114527 87274
rect 110860 87216 114466 87272
rect 114522 87216 114527 87272
rect 110860 87214 114527 87216
rect 114461 87211 114527 87214
rect 521101 87274 521167 87277
rect 523200 87274 524400 87304
rect 521101 87272 524400 87274
rect 521101 87216 521106 87272
rect 521162 87216 524400 87272
rect 521101 87214 524400 87216
rect 521101 87211 521167 87214
rect 523200 87184 524400 87214
rect 520733 86322 520799 86325
rect 518788 86320 520799 86322
rect 518788 86264 520738 86320
rect 520794 86264 520799 86320
rect 518788 86262 520799 86264
rect 520733 86259 520799 86262
rect 520365 85778 520431 85781
rect 523200 85778 524400 85808
rect 520365 85776 524400 85778
rect 520365 85720 520370 85776
rect 520426 85720 524400 85776
rect 520365 85718 524400 85720
rect 520365 85715 520431 85718
rect 523200 85688 524400 85718
rect 116209 85642 116275 85645
rect 116209 85640 119140 85642
rect 116209 85584 116214 85640
rect 116270 85584 119140 85640
rect 116209 85582 119140 85584
rect 116209 85579 116275 85582
rect 521009 84962 521075 84965
rect 518788 84960 521075 84962
rect 518788 84904 521014 84960
rect 521070 84904 521075 84960
rect 518788 84902 521075 84904
rect 521009 84899 521075 84902
rect 520273 84282 520339 84285
rect 523200 84282 524400 84312
rect 520273 84280 524400 84282
rect 520273 84224 520278 84280
rect 520334 84224 524400 84280
rect 520273 84222 524400 84224
rect 520273 84219 520339 84222
rect 523200 84192 524400 84222
rect 115289 83738 115355 83741
rect 115289 83736 119140 83738
rect 115289 83680 115294 83736
rect 115350 83680 119140 83736
rect 115289 83678 119140 83680
rect 115289 83675 115355 83678
rect 521193 83602 521259 83605
rect 518788 83600 521259 83602
rect 518788 83544 521198 83600
rect 521254 83544 521259 83600
rect 518788 83542 521259 83544
rect 521193 83539 521259 83542
rect 520733 82786 520799 82789
rect 523200 82786 524400 82816
rect 520733 82784 524400 82786
rect 520733 82728 520738 82784
rect 520794 82728 524400 82784
rect 520733 82726 524400 82728
rect 520733 82723 520799 82726
rect 523200 82696 524400 82726
rect 521285 82242 521351 82245
rect 518788 82240 521351 82242
rect 518788 82184 521290 82240
rect 521346 82184 521351 82240
rect 518788 82182 521351 82184
rect 521285 82179 521351 82182
rect 115381 81834 115447 81837
rect 115381 81832 119140 81834
rect 115381 81776 115386 81832
rect 115442 81776 119140 81832
rect 115381 81774 119140 81776
rect 115381 81771 115447 81774
rect 521009 81154 521075 81157
rect 523200 81154 524400 81184
rect 521009 81152 524400 81154
rect 521009 81096 521014 81152
rect 521070 81096 524400 81152
rect 521009 81094 524400 81096
rect 521009 81091 521075 81094
rect 523200 81064 524400 81094
rect 521101 80882 521167 80885
rect 518788 80880 521167 80882
rect 518788 80824 521106 80880
rect 521162 80824 521167 80880
rect 518788 80822 521167 80824
rect 521101 80819 521167 80822
rect 116761 79930 116827 79933
rect 116761 79928 119140 79930
rect 116761 79872 116766 79928
rect 116822 79872 119140 79928
rect 116761 79870 119140 79872
rect 116761 79867 116827 79870
rect 521377 79658 521443 79661
rect 523200 79658 524400 79688
rect 521377 79656 524400 79658
rect 521377 79600 521382 79656
rect 521438 79600 524400 79656
rect 521377 79598 524400 79600
rect 521377 79595 521443 79598
rect 523200 79568 524400 79598
rect 520365 79522 520431 79525
rect 518788 79520 520431 79522
rect 518788 79464 520370 79520
rect 520426 79464 520431 79520
rect 518788 79462 520431 79464
rect 520365 79459 520431 79462
rect 520273 78162 520339 78165
rect 518788 78160 520339 78162
rect 518788 78104 520278 78160
rect 520334 78104 520339 78160
rect 518788 78102 520339 78104
rect 520273 78099 520339 78102
rect 521101 78162 521167 78165
rect 523200 78162 524400 78192
rect 521101 78160 524400 78162
rect 521101 78104 521106 78160
rect 521162 78104 524400 78160
rect 521101 78102 524400 78104
rect 521101 78099 521167 78102
rect 523200 78072 524400 78102
rect 116669 78026 116735 78029
rect 116669 78024 119140 78026
rect 116669 77968 116674 78024
rect 116730 77968 119140 78024
rect 116669 77966 119140 77968
rect 116669 77963 116735 77966
rect 520733 76802 520799 76805
rect 518788 76800 520799 76802
rect 518788 76744 520738 76800
rect 520794 76744 520799 76800
rect 518788 76742 520799 76744
rect 520733 76739 520799 76742
rect 520457 76666 520523 76669
rect 523200 76666 524400 76696
rect 520457 76664 524400 76666
rect 520457 76608 520462 76664
rect 520518 76608 524400 76664
rect 520457 76606 524400 76608
rect 520457 76603 520523 76606
rect 523200 76576 524400 76606
rect 110860 75926 119140 75986
rect 521009 75306 521075 75309
rect 518788 75304 521075 75306
rect 518788 75248 521014 75304
rect 521070 75248 521075 75304
rect 518788 75246 521075 75248
rect 521009 75243 521075 75246
rect 520273 75170 520339 75173
rect 523200 75170 524400 75200
rect 520273 75168 524400 75170
rect 520273 75112 520278 75168
rect 520334 75112 524400 75168
rect 520273 75110 524400 75112
rect 520273 75107 520339 75110
rect 523200 75080 524400 75110
rect 116577 74082 116643 74085
rect 116577 74080 119140 74082
rect 116577 74024 116582 74080
rect 116638 74024 119140 74080
rect 116577 74022 119140 74024
rect 116577 74019 116643 74022
rect 521377 73946 521443 73949
rect 518788 73944 521443 73946
rect 518788 73888 521382 73944
rect 521438 73888 521443 73944
rect 518788 73886 521443 73888
rect 521377 73883 521443 73886
rect 520733 73674 520799 73677
rect 523200 73674 524400 73704
rect 520733 73672 524400 73674
rect 520733 73616 520738 73672
rect 520794 73616 524400 73672
rect 520733 73614 524400 73616
rect 520733 73611 520799 73614
rect 523200 73584 524400 73614
rect 521101 72586 521167 72589
rect 518788 72584 521167 72586
rect 518788 72528 521106 72584
rect 521162 72528 521167 72584
rect 518788 72526 521167 72528
rect 521101 72523 521167 72526
rect 116393 72178 116459 72181
rect 116393 72176 119140 72178
rect 116393 72120 116398 72176
rect 116454 72120 119140 72176
rect 116393 72118 119140 72120
rect 116393 72115 116459 72118
rect 521009 72042 521075 72045
rect 523200 72042 524400 72072
rect 521009 72040 524400 72042
rect 521009 71984 521014 72040
rect 521070 71984 524400 72040
rect 521009 71982 524400 71984
rect 521009 71979 521075 71982
rect 523200 71952 524400 71982
rect 520457 71226 520523 71229
rect 518788 71224 520523 71226
rect 518788 71168 520462 71224
rect 520518 71168 520523 71224
rect 518788 71166 520523 71168
rect 520457 71163 520523 71166
rect 521101 70546 521167 70549
rect 523200 70546 524400 70576
rect 521101 70544 524400 70546
rect 521101 70488 521106 70544
rect 521162 70488 524400 70544
rect 521101 70486 524400 70488
rect 521101 70483 521167 70486
rect 523200 70456 524400 70486
rect 116301 70274 116367 70277
rect 116301 70272 119140 70274
rect 116301 70216 116306 70272
rect 116362 70216 119140 70272
rect 116301 70214 119140 70216
rect 116301 70211 116367 70214
rect 520273 69866 520339 69869
rect 518788 69864 520339 69866
rect 518788 69808 520278 69864
rect 520334 69808 520339 69864
rect 518788 69806 520339 69808
rect 520273 69803 520339 69806
rect 521285 69050 521351 69053
rect 523200 69050 524400 69080
rect 521285 69048 524400 69050
rect 521285 68992 521290 69048
rect 521346 68992 524400 69048
rect 521285 68990 524400 68992
rect 521285 68987 521351 68990
rect 523200 68960 524400 68990
rect 520733 68506 520799 68509
rect 518788 68504 520799 68506
rect 518788 68448 520738 68504
rect 520794 68448 520799 68504
rect 518788 68446 520799 68448
rect 520733 68443 520799 68446
rect 116209 68370 116275 68373
rect 116209 68368 119140 68370
rect 116209 68312 116214 68368
rect 116270 68312 119140 68368
rect 116209 68310 119140 68312
rect 116209 68307 116275 68310
rect 520457 67554 520523 67557
rect 523200 67554 524400 67584
rect 520457 67552 524400 67554
rect 520457 67496 520462 67552
rect 520518 67496 524400 67552
rect 520457 67494 524400 67496
rect 520457 67491 520523 67494
rect 523200 67464 524400 67494
rect 521009 67146 521075 67149
rect 518788 67144 521075 67146
rect 518788 67088 521014 67144
rect 521070 67088 521075 67144
rect 518788 67086 521075 67088
rect 521009 67083 521075 67086
rect 116853 66466 116919 66469
rect 116853 66464 119140 66466
rect 116853 66408 116858 66464
rect 116914 66408 119140 66464
rect 116853 66406 119140 66408
rect 116853 66403 116919 66406
rect 520365 66058 520431 66061
rect 523200 66058 524400 66088
rect 520365 66056 524400 66058
rect 520365 66000 520370 66056
rect 520426 66000 524400 66056
rect 520365 65998 524400 66000
rect 520365 65995 520431 65998
rect 523200 65968 524400 65998
rect 521101 65786 521167 65789
rect 518788 65784 521167 65786
rect 518788 65728 521106 65784
rect 521162 65728 521167 65784
rect 518788 65726 521167 65728
rect 521101 65723 521167 65726
rect 114461 64562 114527 64565
rect 110860 64560 114527 64562
rect 110860 64504 114466 64560
rect 114522 64504 114527 64560
rect 110860 64502 114527 64504
rect 114461 64499 114527 64502
rect 115197 64562 115263 64565
rect 520733 64562 520799 64565
rect 523200 64562 524400 64592
rect 115197 64560 119140 64562
rect 115197 64504 115202 64560
rect 115258 64504 119140 64560
rect 115197 64502 119140 64504
rect 520733 64560 524400 64562
rect 520733 64504 520738 64560
rect 520794 64504 524400 64560
rect 520733 64502 524400 64504
rect 115197 64499 115263 64502
rect 520733 64499 520799 64502
rect 523200 64472 524400 64502
rect 521285 64426 521351 64429
rect 518788 64424 521351 64426
rect 518788 64368 521290 64424
rect 521346 64368 521351 64424
rect 518788 64366 521351 64368
rect 521285 64363 521351 64366
rect 520457 63066 520523 63069
rect 518788 63064 520523 63066
rect 518788 63008 520462 63064
rect 520518 63008 520523 63064
rect 518788 63006 520523 63008
rect 520457 63003 520523 63006
rect 521101 62930 521167 62933
rect 523200 62930 524400 62960
rect 521101 62928 524400 62930
rect 521101 62872 521106 62928
rect 521162 62872 524400 62928
rect 521101 62870 524400 62872
rect 521101 62867 521167 62870
rect 523200 62840 524400 62870
rect 116117 62658 116183 62661
rect 116117 62656 119140 62658
rect 116117 62600 116122 62656
rect 116178 62600 119140 62656
rect 116117 62598 119140 62600
rect 116117 62595 116183 62598
rect 520365 61706 520431 61709
rect 518788 61704 520431 61706
rect 518788 61648 520370 61704
rect 520426 61648 520431 61704
rect 518788 61646 520431 61648
rect 520365 61643 520431 61646
rect 521009 61434 521075 61437
rect 523200 61434 524400 61464
rect 521009 61432 524400 61434
rect 521009 61376 521014 61432
rect 521070 61376 524400 61432
rect 521009 61374 524400 61376
rect 521009 61371 521075 61374
rect 523200 61344 524400 61374
rect 116117 60618 116183 60621
rect 116117 60616 119140 60618
rect 116117 60560 116122 60616
rect 116178 60560 119140 60616
rect 116117 60558 119140 60560
rect 116117 60555 116183 60558
rect 520733 60346 520799 60349
rect 518788 60344 520799 60346
rect 518788 60288 520738 60344
rect 520794 60288 520799 60344
rect 518788 60286 520799 60288
rect 520733 60283 520799 60286
rect 520733 59938 520799 59941
rect 523200 59938 524400 59968
rect 520733 59936 524400 59938
rect 520733 59880 520738 59936
rect 520794 59880 524400 59936
rect 520733 59878 524400 59880
rect 520733 59875 520799 59878
rect 523200 59848 524400 59878
rect 521101 58986 521167 58989
rect 518788 58984 521167 58986
rect 518788 58928 521106 58984
rect 521162 58928 521167 58984
rect 518788 58926 521167 58928
rect 521101 58923 521167 58926
rect 117037 58714 117103 58717
rect 117037 58712 119140 58714
rect 117037 58656 117042 58712
rect 117098 58656 119140 58712
rect 117037 58654 119140 58656
rect 117037 58651 117103 58654
rect 521101 58442 521167 58445
rect 523200 58442 524400 58472
rect 521101 58440 524400 58442
rect 521101 58384 521106 58440
rect 521162 58384 524400 58440
rect 521101 58382 524400 58384
rect 521101 58379 521167 58382
rect 523200 58352 524400 58382
rect 521009 57490 521075 57493
rect 518788 57488 521075 57490
rect 518788 57432 521014 57488
rect 521070 57432 521075 57488
rect 518788 57430 521075 57432
rect 521009 57427 521075 57430
rect 520365 56946 520431 56949
rect 523200 56946 524400 56976
rect 520365 56944 524400 56946
rect 520365 56888 520370 56944
rect 520426 56888 524400 56944
rect 520365 56886 524400 56888
rect 520365 56883 520431 56886
rect 523200 56856 524400 56886
rect 117129 56810 117195 56813
rect 117129 56808 119140 56810
rect 117129 56752 117134 56808
rect 117190 56752 119140 56808
rect 117129 56750 119140 56752
rect 117129 56747 117195 56750
rect 520733 56130 520799 56133
rect 518788 56128 520799 56130
rect 518788 56072 520738 56128
rect 520794 56072 520799 56128
rect 518788 56070 520799 56072
rect 520733 56067 520799 56070
rect 520273 55450 520339 55453
rect 523200 55450 524400 55480
rect 520273 55448 524400 55450
rect 520273 55392 520278 55448
rect 520334 55392 524400 55448
rect 520273 55390 524400 55392
rect 520273 55387 520339 55390
rect 523200 55360 524400 55390
rect 116577 54906 116643 54909
rect 116577 54904 119140 54906
rect 116577 54848 116582 54904
rect 116638 54848 119140 54904
rect 116577 54846 119140 54848
rect 116577 54843 116643 54846
rect 521101 54770 521167 54773
rect 518788 54768 521167 54770
rect 518788 54712 521106 54768
rect 521162 54712 521167 54768
rect 518788 54710 521167 54712
rect 521101 54707 521167 54710
rect 521101 53818 521167 53821
rect 523200 53818 524400 53848
rect 521101 53816 524400 53818
rect 521101 53760 521106 53816
rect 521162 53760 524400 53816
rect 521101 53758 524400 53760
rect 521101 53755 521167 53758
rect 523200 53728 524400 53758
rect 520365 53410 520431 53413
rect 518788 53408 520431 53410
rect 518788 53352 520370 53408
rect 520426 53352 520431 53408
rect 518788 53350 520431 53352
rect 520365 53347 520431 53350
rect 113817 53138 113883 53141
rect 110860 53136 113883 53138
rect 110860 53080 113822 53136
rect 113878 53080 113883 53136
rect 110860 53078 113883 53080
rect 113817 53075 113883 53078
rect 116669 53002 116735 53005
rect 116669 53000 119140 53002
rect 116669 52944 116674 53000
rect 116730 52944 119140 53000
rect 116669 52942 119140 52944
rect 116669 52939 116735 52942
rect 520917 52322 520983 52325
rect 523200 52322 524400 52352
rect 520917 52320 524400 52322
rect 520917 52264 520922 52320
rect 520978 52264 524400 52320
rect 520917 52262 524400 52264
rect 520917 52259 520983 52262
rect 523200 52232 524400 52262
rect 520273 52050 520339 52053
rect 518788 52048 520339 52050
rect 518788 51992 520278 52048
rect 520334 51992 520339 52048
rect 518788 51990 520339 51992
rect 520273 51987 520339 51990
rect 115933 51098 115999 51101
rect 115933 51096 119140 51098
rect 115933 51040 115938 51096
rect 115994 51040 119140 51096
rect 115933 51038 119140 51040
rect 115933 51035 115999 51038
rect 520365 50826 520431 50829
rect 523200 50826 524400 50856
rect 520365 50824 524400 50826
rect 520365 50768 520370 50824
rect 520426 50768 524400 50824
rect 520365 50766 524400 50768
rect 520365 50763 520431 50766
rect 523200 50736 524400 50766
rect 521101 50690 521167 50693
rect 518788 50688 521167 50690
rect 518788 50632 521106 50688
rect 521162 50632 521167 50688
rect 518788 50630 521167 50632
rect 521101 50627 521167 50630
rect 520917 49330 520983 49333
rect 518788 49328 520983 49330
rect 518788 49272 520922 49328
rect 520978 49272 520983 49328
rect 518788 49270 520983 49272
rect 520917 49267 520983 49270
rect 521101 49330 521167 49333
rect 523200 49330 524400 49360
rect 521101 49328 524400 49330
rect 521101 49272 521106 49328
rect 521162 49272 524400 49328
rect 521101 49270 524400 49272
rect 521101 49267 521167 49270
rect 523200 49240 524400 49270
rect 116761 49194 116827 49197
rect 116761 49192 119140 49194
rect 116761 49136 116766 49192
rect 116822 49136 119140 49192
rect 116761 49134 119140 49136
rect 116761 49131 116827 49134
rect 520365 47970 520431 47973
rect 518788 47968 520431 47970
rect 518788 47912 520370 47968
rect 520426 47912 520431 47968
rect 518788 47910 520431 47912
rect 520365 47907 520431 47910
rect 520273 47834 520339 47837
rect 523200 47834 524400 47864
rect 520273 47832 524400 47834
rect 520273 47776 520278 47832
rect 520334 47776 524400 47832
rect 520273 47774 524400 47776
rect 520273 47771 520339 47774
rect 523200 47744 524400 47774
rect 116025 47154 116091 47157
rect 116025 47152 119140 47154
rect 116025 47096 116030 47152
rect 116086 47096 119140 47152
rect 116025 47094 119140 47096
rect 116025 47091 116091 47094
rect 521101 46610 521167 46613
rect 518788 46608 521167 46610
rect 518788 46552 521106 46608
rect 521162 46552 521167 46608
rect 518788 46550 521167 46552
rect 521101 46547 521167 46550
rect 520365 46338 520431 46341
rect 523200 46338 524400 46368
rect 520365 46336 524400 46338
rect 520365 46280 520370 46336
rect 520426 46280 524400 46336
rect 520365 46278 524400 46280
rect 520365 46275 520431 46278
rect 523200 46248 524400 46278
rect 116853 45250 116919 45253
rect 520273 45250 520339 45253
rect 116853 45248 119140 45250
rect 116853 45192 116858 45248
rect 116914 45192 119140 45248
rect 116853 45190 119140 45192
rect 518788 45248 520339 45250
rect 518788 45192 520278 45248
rect 520334 45192 520339 45248
rect 518788 45190 520339 45192
rect 116853 45187 116919 45190
rect 520273 45187 520339 45190
rect 521009 44706 521075 44709
rect 523200 44706 524400 44736
rect 521009 44704 524400 44706
rect 521009 44648 521014 44704
rect 521070 44648 524400 44704
rect 521009 44646 524400 44648
rect 521009 44643 521075 44646
rect 523200 44616 524400 44646
rect 520365 43890 520431 43893
rect 518788 43888 520431 43890
rect 518788 43832 520370 43888
rect 520426 43832 520431 43888
rect 518788 43830 520431 43832
rect 520365 43827 520431 43830
rect 116393 43346 116459 43349
rect 116393 43344 119140 43346
rect 116393 43288 116398 43344
rect 116454 43288 119140 43344
rect 116393 43286 119140 43288
rect 116393 43283 116459 43286
rect 521101 43210 521167 43213
rect 523200 43210 524400 43240
rect 521101 43208 524400 43210
rect 521101 43152 521106 43208
rect 521162 43152 524400 43208
rect 521101 43150 524400 43152
rect 521101 43147 521167 43150
rect 523200 43120 524400 43150
rect 521009 42530 521075 42533
rect 518788 42528 521075 42530
rect 518788 42472 521014 42528
rect 521070 42472 521075 42528
rect 518788 42470 521075 42472
rect 521009 42467 521075 42470
rect 114093 41850 114159 41853
rect 110860 41848 114159 41850
rect 110860 41792 114098 41848
rect 114154 41792 114159 41848
rect 110860 41790 114159 41792
rect 114093 41787 114159 41790
rect 521009 41714 521075 41717
rect 523200 41714 524400 41744
rect 521009 41712 524400 41714
rect 521009 41656 521014 41712
rect 521070 41656 524400 41712
rect 521009 41654 524400 41656
rect 521009 41651 521075 41654
rect 523200 41624 524400 41654
rect 116945 41442 117011 41445
rect 116945 41440 119140 41442
rect 116945 41384 116950 41440
rect 117006 41384 119140 41440
rect 116945 41382 119140 41384
rect 116945 41379 117011 41382
rect 521101 41170 521167 41173
rect 518788 41168 521167 41170
rect 518788 41112 521106 41168
rect 521162 41112 521167 41168
rect 518788 41110 521167 41112
rect 521101 41107 521167 41110
rect 521101 40218 521167 40221
rect 523200 40218 524400 40248
rect 521101 40216 524400 40218
rect 521101 40160 521106 40216
rect 521162 40160 524400 40216
rect 521101 40158 524400 40160
rect 521101 40155 521167 40158
rect 523200 40128 524400 40158
rect 521009 39810 521075 39813
rect 518788 39808 521075 39810
rect 518788 39752 521014 39808
rect 521070 39752 521075 39808
rect 518788 39750 521075 39752
rect 521009 39747 521075 39750
rect 115933 39538 115999 39541
rect 115933 39536 119140 39538
rect 115933 39480 115938 39536
rect 115994 39480 119140 39536
rect 115933 39478 119140 39480
rect 115933 39475 115999 39478
rect 520917 38722 520983 38725
rect 523200 38722 524400 38752
rect 520917 38720 524400 38722
rect 520917 38664 520922 38720
rect 520978 38664 524400 38720
rect 520917 38662 524400 38664
rect 520917 38659 520983 38662
rect 523200 38632 524400 38662
rect 521101 38314 521167 38317
rect 518788 38312 521167 38314
rect 518788 38256 521106 38312
rect 521162 38256 521167 38312
rect 518788 38254 521167 38256
rect 521101 38251 521167 38254
rect 116117 37634 116183 37637
rect 116117 37632 119140 37634
rect 116117 37576 116122 37632
rect 116178 37576 119140 37632
rect 116117 37574 119140 37576
rect 116117 37571 116183 37574
rect 521101 37226 521167 37229
rect 523200 37226 524400 37256
rect 521101 37224 524400 37226
rect 521101 37168 521106 37224
rect 521162 37168 524400 37224
rect 521101 37166 524400 37168
rect 521101 37163 521167 37166
rect 523200 37136 524400 37166
rect 520917 36954 520983 36957
rect 518788 36952 520983 36954
rect 518788 36896 520922 36952
rect 520978 36896 520983 36952
rect 518788 36894 520983 36896
rect 520917 36891 520983 36894
rect 521101 36002 521167 36005
rect 518758 36000 521167 36002
rect 518758 35944 521106 36000
rect 521162 35944 521167 36000
rect 518758 35942 521167 35944
rect 117129 35730 117195 35733
rect 117129 35728 119140 35730
rect 117129 35672 117134 35728
rect 117190 35672 119140 35728
rect 117129 35670 119140 35672
rect 117129 35667 117195 35670
rect 518758 35564 518818 35942
rect 521101 35939 521167 35942
rect 520917 35594 520983 35597
rect 523200 35594 524400 35624
rect 520917 35592 524400 35594
rect 520917 35536 520922 35592
rect 520978 35536 524400 35592
rect 520917 35534 524400 35536
rect 520917 35531 520983 35534
rect 523200 35504 524400 35534
rect 520917 34642 520983 34645
rect 518758 34640 520983 34642
rect 518758 34584 520922 34640
rect 520978 34584 520983 34640
rect 518758 34582 520983 34584
rect 518758 34204 518818 34582
rect 520917 34579 520983 34582
rect 520825 34098 520891 34101
rect 523200 34098 524400 34128
rect 520825 34096 524400 34098
rect 520825 34040 520830 34096
rect 520886 34040 524400 34096
rect 520825 34038 524400 34040
rect 520825 34035 520891 34038
rect 523200 34008 524400 34038
rect 116117 33826 116183 33829
rect 116117 33824 119140 33826
rect 116117 33768 116122 33824
rect 116178 33768 119140 33824
rect 116117 33766 119140 33768
rect 116117 33763 116183 33766
rect 520825 33282 520891 33285
rect 518758 33280 520891 33282
rect 518758 33224 520830 33280
rect 520886 33224 520891 33280
rect 518758 33222 520891 33224
rect 518758 32844 518818 33222
rect 520825 33219 520891 33222
rect 521101 32602 521167 32605
rect 523200 32602 524400 32632
rect 521101 32600 524400 32602
rect 521101 32544 521106 32600
rect 521162 32544 524400 32600
rect 521101 32542 524400 32544
rect 521101 32539 521167 32542
rect 523200 32512 524400 32542
rect 116485 31786 116551 31789
rect 521101 31786 521167 31789
rect 116485 31784 119140 31786
rect 116485 31728 116490 31784
rect 116546 31728 119140 31784
rect 116485 31726 119140 31728
rect 518758 31784 521167 31786
rect 518758 31728 521106 31784
rect 521162 31728 521167 31784
rect 518758 31726 521167 31728
rect 116485 31723 116551 31726
rect 518758 31484 518818 31726
rect 521101 31723 521167 31726
rect 521101 31106 521167 31109
rect 523200 31106 524400 31136
rect 521101 31104 524400 31106
rect 521101 31048 521106 31104
rect 521162 31048 524400 31104
rect 521101 31046 524400 31048
rect 521101 31043 521167 31046
rect 523200 31016 524400 31046
rect 114185 30426 114251 30429
rect 521101 30426 521167 30429
rect 110860 30424 114251 30426
rect 110860 30368 114190 30424
rect 114246 30368 114251 30424
rect 110860 30366 114251 30368
rect 114185 30363 114251 30366
rect 518758 30424 521167 30426
rect 518758 30368 521106 30424
rect 521162 30368 521167 30424
rect 518758 30366 521167 30368
rect 518758 30124 518818 30366
rect 521101 30363 521167 30366
rect 116393 29882 116459 29885
rect 116393 29880 119140 29882
rect 116393 29824 116398 29880
rect 116454 29824 119140 29880
rect 116393 29822 119140 29824
rect 116393 29819 116459 29822
rect 521101 29610 521167 29613
rect 523200 29610 524400 29640
rect 521101 29608 524400 29610
rect 521101 29552 521106 29608
rect 521162 29552 524400 29608
rect 521101 29550 524400 29552
rect 521101 29547 521167 29550
rect 523200 29520 524400 29550
rect 521101 28794 521167 28797
rect 518788 28792 521167 28794
rect 518788 28736 521106 28792
rect 521162 28736 521167 28792
rect 518788 28734 521167 28736
rect 521101 28731 521167 28734
rect 523200 28114 524400 28144
rect 518850 28054 524400 28114
rect 116117 27978 116183 27981
rect 518850 27978 518910 28054
rect 523200 28024 524400 28054
rect 116117 27976 119140 27978
rect 116117 27920 116122 27976
rect 116178 27920 119140 27976
rect 116117 27918 119140 27920
rect 518758 27918 518910 27978
rect 116117 27915 116183 27918
rect 518758 27404 518818 27918
rect 523200 26482 524400 26512
rect 518850 26422 524400 26482
rect 518850 26346 518910 26422
rect 523200 26392 524400 26422
rect 518758 26286 518910 26346
rect 116526 26012 116532 26076
rect 116596 26074 116602 26076
rect 116596 26014 119140 26074
rect 518758 26044 518818 26286
rect 116596 26012 116602 26014
rect 523200 24986 524400 25016
rect 518758 24926 524400 24986
rect 518758 24684 518818 24926
rect 523200 24896 524400 24926
rect 116117 24170 116183 24173
rect 116117 24168 119140 24170
rect 116117 24112 116122 24168
rect 116178 24112 119140 24168
rect 116117 24110 119140 24112
rect 116117 24107 116183 24110
rect 523200 23490 524400 23520
rect 518758 23430 524400 23490
rect 518758 23324 518818 23430
rect 523200 23400 524400 23430
rect 116117 22266 116183 22269
rect 116117 22264 119140 22266
rect 116117 22208 116122 22264
rect 116178 22208 119140 22264
rect 116117 22206 119140 22208
rect 116117 22203 116183 22206
rect 523200 21994 524400 22024
rect 518788 21934 524400 21994
rect 523200 21904 524400 21934
rect 521101 20498 521167 20501
rect 523200 20498 524400 20528
rect 521101 20496 524400 20498
rect 116117 20362 116183 20365
rect 116117 20360 119140 20362
rect 116117 20304 116122 20360
rect 116178 20304 119140 20360
rect 116117 20302 119140 20304
rect 116117 20299 116183 20302
rect 518758 19818 518818 20468
rect 521101 20440 521106 20496
rect 521162 20440 524400 20496
rect 521101 20438 524400 20440
rect 521101 20435 521167 20438
rect 523200 20408 524400 20438
rect 521101 19818 521167 19821
rect 518758 19816 521167 19818
rect 518758 19760 521106 19816
rect 521162 19760 521167 19816
rect 518758 19758 521167 19760
rect 521101 19755 521167 19758
rect 114277 19002 114343 19005
rect 110860 19000 114343 19002
rect 110860 18944 114282 19000
rect 114338 18944 114343 19000
rect 110860 18942 114343 18944
rect 114277 18939 114343 18942
rect 116117 18458 116183 18461
rect 518758 18458 518818 19108
rect 523200 19002 524400 19032
rect 521150 18942 524400 19002
rect 521150 18458 521210 18942
rect 523200 18912 524400 18942
rect 116117 18456 119140 18458
rect 116117 18400 116122 18456
rect 116178 18400 119140 18456
rect 116117 18398 119140 18400
rect 518758 18398 521210 18458
rect 116117 18395 116183 18398
rect 518758 17098 518818 17748
rect 523200 17370 524400 17400
rect 521150 17310 524400 17370
rect 521150 17098 521210 17310
rect 523200 17280 524400 17310
rect 518758 17038 521210 17098
rect 116117 16418 116183 16421
rect 116117 16416 119140 16418
rect 116117 16360 116122 16416
rect 116178 16360 119140 16416
rect 116117 16358 119140 16360
rect 116117 16355 116183 16358
rect 518758 15738 518818 16388
rect 523200 15874 524400 15904
rect 521104 15814 524400 15874
rect 521104 15738 521164 15814
rect 523200 15784 524400 15814
rect 518758 15678 521164 15738
rect 521101 15058 521167 15061
rect 518788 15056 521167 15058
rect 518788 15000 521106 15056
rect 521162 15000 521167 15056
rect 518788 14998 521167 15000
rect 521101 14995 521167 14998
rect 115933 14514 115999 14517
rect 115933 14512 119140 14514
rect 115933 14456 115938 14512
rect 115994 14456 119140 14512
rect 115933 14454 119140 14456
rect 115933 14451 115999 14454
rect 521101 14378 521167 14381
rect 523200 14378 524400 14408
rect 521101 14376 524400 14378
rect 521101 14320 521106 14376
rect 521162 14320 524400 14376
rect 521101 14318 524400 14320
rect 521101 14315 521167 14318
rect 523200 14288 524400 14318
rect 521101 13698 521167 13701
rect 518788 13696 521167 13698
rect 518788 13640 521106 13696
rect 521162 13640 521167 13696
rect 518788 13638 521167 13640
rect 521101 13635 521167 13638
rect 521101 12882 521167 12885
rect 523200 12882 524400 12912
rect 521101 12880 524400 12882
rect 521101 12824 521106 12880
rect 521162 12824 524400 12880
rect 521101 12822 524400 12824
rect 521101 12819 521167 12822
rect 523200 12792 524400 12822
rect 117037 12610 117103 12613
rect 117037 12608 119140 12610
rect 117037 12552 117042 12608
rect 117098 12552 119140 12608
rect 117037 12550 119140 12552
rect 117037 12547 117103 12550
rect 519629 12338 519695 12341
rect 518788 12336 519695 12338
rect 518788 12280 519634 12336
rect 519690 12280 519695 12336
rect 518788 12278 519695 12280
rect 519629 12275 519695 12278
rect 519629 11386 519695 11389
rect 523200 11386 524400 11416
rect 519629 11384 524400 11386
rect 519629 11328 519634 11384
rect 519690 11328 524400 11384
rect 519629 11326 524400 11328
rect 519629 11323 519695 11326
rect 523200 11296 524400 11326
rect 521101 10978 521167 10981
rect 518788 10976 521167 10978
rect 518788 10920 521106 10976
rect 521162 10920 521167 10976
rect 518788 10918 521167 10920
rect 521101 10915 521167 10918
rect 117221 10706 117287 10709
rect 117221 10704 119140 10706
rect 117221 10648 117226 10704
rect 117282 10648 119140 10704
rect 117221 10646 119140 10648
rect 117221 10643 117287 10646
rect 521101 9890 521167 9893
rect 523200 9890 524400 9920
rect 521101 9888 524400 9890
rect 521101 9832 521106 9888
rect 521162 9832 524400 9888
rect 521101 9830 524400 9832
rect 521101 9827 521167 9830
rect 523200 9800 524400 9830
rect 521101 9618 521167 9621
rect 518788 9616 521167 9618
rect 518788 9560 521106 9616
rect 521162 9560 521167 9616
rect 518788 9558 521167 9560
rect 521101 9555 521167 9558
rect 117078 8740 117084 8804
rect 117148 8802 117154 8804
rect 117148 8742 119140 8802
rect 117148 8740 117154 8742
rect 520365 8258 520431 8261
rect 518788 8256 520431 8258
rect 518788 8200 520370 8256
rect 520426 8200 520431 8256
rect 518788 8198 520431 8200
rect 520365 8195 520431 8198
rect 521101 8258 521167 8261
rect 523200 8258 524400 8288
rect 521101 8256 524400 8258
rect 521101 8200 521106 8256
rect 521162 8200 524400 8256
rect 521101 8198 524400 8200
rect 521101 8195 521167 8198
rect 523200 8168 524400 8198
rect 114185 7714 114251 7717
rect 110860 7712 114251 7714
rect 110860 7656 114190 7712
rect 114246 7656 114251 7712
rect 110860 7654 114251 7656
rect 114185 7651 114251 7654
rect 116158 6836 116164 6900
rect 116228 6898 116234 6900
rect 521101 6898 521167 6901
rect 116228 6838 119140 6898
rect 518788 6896 521167 6898
rect 518788 6840 521106 6896
rect 521162 6840 521167 6896
rect 518788 6838 521167 6840
rect 116228 6836 116234 6838
rect 521101 6835 521167 6838
rect 520365 6762 520431 6765
rect 523200 6762 524400 6792
rect 520365 6760 524400 6762
rect 520365 6704 520370 6760
rect 520426 6704 524400 6760
rect 520365 6702 524400 6704
rect 520365 6699 520431 6702
rect 523200 6672 524400 6702
rect 521009 5538 521075 5541
rect 518788 5536 521075 5538
rect 518788 5480 521014 5536
rect 521070 5480 521075 5536
rect 518788 5478 521075 5480
rect 521009 5475 521075 5478
rect 521101 5266 521167 5269
rect 523200 5266 524400 5296
rect 521101 5264 524400 5266
rect 521101 5208 521106 5264
rect 521162 5208 524400 5264
rect 521101 5206 524400 5208
rect 521101 5203 521167 5206
rect 523200 5176 524400 5206
rect 116025 4994 116091 4997
rect 116025 4992 119140 4994
rect 116025 4936 116030 4992
rect 116086 4936 119140 4992
rect 116025 4934 119140 4936
rect 116025 4931 116091 4934
rect 520917 4178 520983 4181
rect 518788 4176 520983 4178
rect 518788 4120 520922 4176
rect 520978 4120 520983 4176
rect 518788 4118 520983 4120
rect 520917 4115 520983 4118
rect 521009 3770 521075 3773
rect 523200 3770 524400 3800
rect 521009 3768 524400 3770
rect 521009 3712 521014 3768
rect 521070 3712 524400 3768
rect 521009 3710 524400 3712
rect 521009 3707 521075 3710
rect 523200 3680 524400 3710
rect 116117 3090 116183 3093
rect 116117 3088 119140 3090
rect 116117 3032 116122 3088
rect 116178 3032 119140 3088
rect 116117 3030 119140 3032
rect 116117 3027 116183 3030
rect 521101 2818 521167 2821
rect 518788 2816 521167 2818
rect 518788 2760 521106 2816
rect 521162 2760 521167 2816
rect 518788 2758 521167 2760
rect 521101 2755 521167 2758
rect 42701 2274 42767 2277
rect 116526 2274 116532 2276
rect 42701 2272 116532 2274
rect 42701 2216 42706 2272
rect 42762 2216 116532 2272
rect 42701 2214 116532 2216
rect 42701 2211 42767 2214
rect 116526 2212 116532 2214
rect 116596 2212 116602 2276
rect 520917 2274 520983 2277
rect 523200 2274 524400 2304
rect 520917 2272 524400 2274
rect 520917 2216 520922 2272
rect 520978 2216 524400 2272
rect 520917 2214 524400 2216
rect 520917 2211 520983 2214
rect 523200 2184 524400 2214
rect 29545 2138 29611 2141
rect 111425 2138 111491 2141
rect 29545 2136 111491 2138
rect 29545 2080 29550 2136
rect 29606 2080 111430 2136
rect 111486 2080 111491 2136
rect 29545 2078 111491 2080
rect 29545 2075 29611 2078
rect 111425 2075 111491 2078
rect 26049 2002 26115 2005
rect 111609 2002 111675 2005
rect 26049 2000 111675 2002
rect 26049 1944 26054 2000
rect 26110 1944 111614 2000
rect 111670 1944 111675 2000
rect 26049 1942 111675 1944
rect 26049 1939 26115 1942
rect 111609 1939 111675 1942
rect 15929 1866 15995 1869
rect 109953 1866 110019 1869
rect 343955 1868 344021 1869
rect 343950 1866 343956 1868
rect 15929 1864 110019 1866
rect 15929 1808 15934 1864
rect 15990 1808 109958 1864
rect 110014 1808 110019 1864
rect 15929 1806 110019 1808
rect 343864 1806 343956 1866
rect 15929 1803 15995 1806
rect 109953 1803 110019 1806
rect 343950 1804 343956 1806
rect 344020 1804 344026 1868
rect 343955 1803 344021 1804
rect 19333 1730 19399 1733
rect 117037 1730 117103 1733
rect 19333 1728 117103 1730
rect 19333 1672 19338 1728
rect 19394 1672 117042 1728
rect 117098 1672 117103 1728
rect 19333 1670 117103 1672
rect 19333 1667 19399 1670
rect 117037 1667 117103 1670
rect 5993 1594 6059 1597
rect 116025 1594 116091 1597
rect 5993 1592 116091 1594
rect 5993 1536 5998 1592
rect 6054 1536 116030 1592
rect 116086 1536 116091 1592
rect 5993 1534 116091 1536
rect 5993 1531 6059 1534
rect 116025 1531 116091 1534
rect 55949 1458 56015 1461
rect 294781 1458 294847 1461
rect 295333 1458 295399 1461
rect 55949 1456 295399 1458
rect 55949 1400 55954 1456
rect 56010 1400 294786 1456
rect 294842 1400 295338 1456
rect 295394 1400 295399 1456
rect 55949 1398 295399 1400
rect 55949 1395 56015 1398
rect 294781 1395 294847 1398
rect 295333 1395 295399 1398
rect 97993 1322 98059 1325
rect 117078 1322 117084 1324
rect 97993 1320 117084 1322
rect 97993 1264 97998 1320
rect 98054 1264 117084 1320
rect 97993 1262 117084 1264
rect 97993 1259 98059 1262
rect 117078 1260 117084 1262
rect 117148 1260 117154 1324
rect 100753 1186 100819 1189
rect 116158 1186 116164 1188
rect 100753 1184 116164 1186
rect 100753 1128 100758 1184
rect 100814 1128 116164 1184
rect 100753 1126 116164 1128
rect 100753 1123 100819 1126
rect 116158 1124 116164 1126
rect 116228 1124 116234 1188
rect 163773 1050 163839 1053
rect 193673 1052 193739 1053
rect 164182 1050 164188 1052
rect 163773 1048 164188 1050
rect 163773 992 163778 1048
rect 163834 992 164188 1048
rect 163773 990 164188 992
rect 163773 987 163839 990
rect 164182 988 164188 990
rect 164252 988 164258 1052
rect 193622 1050 193628 1052
rect 193582 990 193628 1050
rect 193692 1048 193739 1052
rect 193734 992 193739 1048
rect 193622 988 193628 990
rect 193692 988 193739 992
rect 193673 987 193739 988
rect 229277 1050 229343 1053
rect 231158 1050 231164 1052
rect 229277 1048 231164 1050
rect 229277 992 229282 1048
rect 229338 992 231164 1048
rect 229277 990 231164 992
rect 229277 987 229343 990
rect 231158 988 231164 990
rect 231228 988 231234 1052
rect 241830 988 241836 1052
rect 241900 1050 241906 1052
rect 243721 1050 243787 1053
rect 241900 1048 243787 1050
rect 241900 992 243726 1048
rect 243782 992 243787 1048
rect 241900 990 243787 992
rect 241900 988 241906 990
rect 243721 987 243787 990
rect 360142 988 360148 1052
rect 360212 1050 360218 1052
rect 360285 1050 360351 1053
rect 360212 1048 360351 1050
rect 360212 992 360290 1048
rect 360346 992 360351 1048
rect 360212 990 360351 992
rect 360212 988 360218 990
rect 360285 987 360351 990
rect 521101 778 521167 781
rect 523200 778 524400 808
rect 521101 776 524400 778
rect 521101 720 521106 776
rect 521162 720 524400 776
rect 521101 718 524400 720
rect 521101 715 521167 718
rect 523200 688 524400 718
<< via3 >>
rect 116532 151812 116596 151876
rect 116532 89388 116596 89452
rect 116532 26012 116596 26076
rect 117084 8740 117148 8804
rect 116164 6836 116228 6900
rect 116532 2212 116596 2276
rect 343956 1864 344020 1868
rect 343956 1808 343960 1864
rect 343960 1808 344016 1864
rect 344016 1808 344020 1864
rect 343956 1804 344020 1808
rect 117084 1260 117148 1324
rect 116164 1124 116228 1188
rect 164188 988 164252 1052
rect 193628 1048 193692 1052
rect 193628 992 193678 1048
rect 193678 992 193692 1048
rect 193628 988 193692 992
rect 231164 988 231228 1052
rect 241836 988 241900 1052
rect 360148 988 360212 1052
<< metal4 >>
rect 116531 151876 116597 151877
rect 116531 151812 116532 151876
rect 116596 151812 116597 151876
rect 116531 151811 116597 151812
rect 1096 148624 1332 148666
rect 1096 148346 1332 148388
rect 110616 148624 110936 148666
rect 110616 148388 110658 148624
rect 110894 148388 110936 148624
rect 110616 148346 110936 148388
rect 1664 135624 1984 135666
rect 1664 135388 1706 135624
rect 1942 135388 1984 135624
rect 1664 135346 1984 135388
rect 109956 135624 110276 135666
rect 109956 135388 109998 135624
rect 110234 135388 110276 135624
rect 109956 135346 110276 135388
rect 1096 122624 1332 122666
rect 1096 122346 1332 122388
rect 110616 122624 110936 122666
rect 110616 122388 110658 122624
rect 110894 122388 110936 122624
rect 110616 122346 110936 122388
rect 1664 109624 1984 109666
rect 1664 109388 1706 109624
rect 1942 109388 1984 109624
rect 1664 109346 1984 109388
rect 109956 109624 110276 109666
rect 109956 109388 109998 109624
rect 110234 109388 110276 109624
rect 109956 109346 110276 109388
rect 1096 96624 1332 96666
rect 1096 96346 1332 96388
rect 110616 96624 110936 96666
rect 110616 96388 110658 96624
rect 110894 96388 110936 96624
rect 110616 96346 110936 96388
rect 116534 89453 116594 151811
rect 119004 148624 119324 148666
rect 119004 148388 119046 148624
rect 119282 148388 119324 148624
rect 119004 148346 119324 148388
rect 518600 148624 518920 148666
rect 518600 148388 518642 148624
rect 518878 148388 518920 148624
rect 518600 148346 518920 148388
rect 119664 135624 119984 135666
rect 119664 135388 119706 135624
rect 119942 135388 119984 135624
rect 119664 135346 119984 135388
rect 517940 135624 518260 135666
rect 517940 135388 517982 135624
rect 518218 135388 518260 135624
rect 517940 135346 518260 135388
rect 119004 122624 119324 122666
rect 119004 122388 119046 122624
rect 119282 122388 119324 122624
rect 119004 122346 119324 122388
rect 518600 122624 518920 122666
rect 518600 122388 518642 122624
rect 518878 122388 518920 122624
rect 518600 122346 518920 122388
rect 119664 109624 119984 109666
rect 119664 109388 119706 109624
rect 119942 109388 119984 109624
rect 119664 109346 119984 109388
rect 517940 109624 518260 109666
rect 517940 109388 517982 109624
rect 518218 109388 518260 109624
rect 517940 109346 518260 109388
rect 119004 96624 119324 96666
rect 119004 96388 119046 96624
rect 119282 96388 119324 96624
rect 119004 96346 119324 96388
rect 518600 96624 518920 96666
rect 518600 96388 518642 96624
rect 518878 96388 518920 96624
rect 518600 96346 518920 96388
rect 116531 89452 116597 89453
rect 116531 89388 116532 89452
rect 116596 89388 116597 89452
rect 116531 89387 116597 89388
rect 1664 83624 1984 83666
rect 1664 83388 1706 83624
rect 1942 83388 1984 83624
rect 1664 83346 1984 83388
rect 109956 83624 110276 83666
rect 109956 83388 109998 83624
rect 110234 83388 110276 83624
rect 109956 83346 110276 83388
rect 119664 83624 119984 83666
rect 119664 83388 119706 83624
rect 119942 83388 119984 83624
rect 119664 83346 119984 83388
rect 517940 83624 518260 83666
rect 517940 83388 517982 83624
rect 518218 83388 518260 83624
rect 517940 83346 518260 83388
rect 1096 70624 1332 70666
rect 1096 70346 1332 70388
rect 110616 70624 110936 70666
rect 110616 70388 110658 70624
rect 110894 70388 110936 70624
rect 110616 70346 110936 70388
rect 119004 70624 119324 70666
rect 119004 70388 119046 70624
rect 119282 70388 119324 70624
rect 119004 70346 119324 70388
rect 518600 70624 518920 70666
rect 518600 70388 518642 70624
rect 518878 70388 518920 70624
rect 518600 70346 518920 70388
rect 1664 57624 1984 57666
rect 1664 57388 1706 57624
rect 1942 57388 1984 57624
rect 1664 57346 1984 57388
rect 109956 57624 110276 57666
rect 109956 57388 109998 57624
rect 110234 57388 110276 57624
rect 109956 57346 110276 57388
rect 119664 57624 119984 57666
rect 119664 57388 119706 57624
rect 119942 57388 119984 57624
rect 119664 57346 119984 57388
rect 517940 57624 518260 57666
rect 517940 57388 517982 57624
rect 518218 57388 518260 57624
rect 517940 57346 518260 57388
rect 1096 44624 1332 44666
rect 1096 44346 1332 44388
rect 110616 44624 110936 44666
rect 110616 44388 110658 44624
rect 110894 44388 110936 44624
rect 110616 44346 110936 44388
rect 119004 44624 119324 44666
rect 119004 44388 119046 44624
rect 119282 44388 119324 44624
rect 119004 44346 119324 44388
rect 518600 44624 518920 44666
rect 518600 44388 518642 44624
rect 518878 44388 518920 44624
rect 518600 44346 518920 44388
rect 1664 31624 1984 31666
rect 1664 31388 1706 31624
rect 1942 31388 1984 31624
rect 1664 31346 1984 31388
rect 109956 31624 110276 31666
rect 109956 31388 109998 31624
rect 110234 31388 110276 31624
rect 109956 31346 110276 31388
rect 119664 31624 119984 31666
rect 119664 31388 119706 31624
rect 119942 31388 119984 31624
rect 119664 31346 119984 31388
rect 517940 31624 518260 31666
rect 517940 31388 517982 31624
rect 518218 31388 518260 31624
rect 517940 31346 518260 31388
rect 116531 26076 116597 26077
rect 116531 26012 116532 26076
rect 116596 26012 116597 26076
rect 116531 26011 116597 26012
rect 1096 18624 1332 18666
rect 1096 18346 1332 18388
rect 110616 18624 110936 18666
rect 110616 18388 110658 18624
rect 110894 18388 110936 18624
rect 110616 18346 110936 18388
rect 116163 6900 116229 6901
rect 116163 6836 116164 6900
rect 116228 6836 116229 6900
rect 116163 6835 116229 6836
rect 1664 5624 1984 5666
rect 1664 5388 1706 5624
rect 1942 5388 1984 5624
rect 1664 5346 1984 5388
rect 109956 5624 110276 5666
rect 109956 5388 109998 5624
rect 110234 5388 110276 5624
rect 109956 5346 110276 5388
rect 116166 1189 116226 6835
rect 116534 2277 116594 26011
rect 119004 18624 119324 18666
rect 119004 18388 119046 18624
rect 119282 18388 119324 18624
rect 119004 18346 119324 18388
rect 518600 18624 518920 18666
rect 518600 18388 518642 18624
rect 518878 18388 518920 18624
rect 518600 18346 518920 18388
rect 117083 8804 117149 8805
rect 117083 8740 117084 8804
rect 117148 8740 117149 8804
rect 117083 8739 117149 8740
rect 116531 2276 116597 2277
rect 116531 2212 116532 2276
rect 116596 2212 116597 2276
rect 116531 2211 116597 2212
rect 117086 1325 117146 8739
rect 119664 5624 119984 5666
rect 119664 5388 119706 5624
rect 119942 5388 119984 5624
rect 119664 5346 119984 5388
rect 517940 5624 518260 5666
rect 517940 5388 517982 5624
rect 518218 5388 518260 5624
rect 517940 5346 518260 5388
rect 343955 1868 344021 1869
rect 343955 1804 343956 1868
rect 344020 1804 344021 1868
rect 343955 1803 344021 1804
rect 117083 1324 117149 1325
rect 117083 1260 117084 1324
rect 117148 1260 117149 1324
rect 117083 1259 117149 1260
rect 116163 1188 116229 1189
rect 116163 1124 116164 1188
rect 116228 1124 116229 1188
rect 343958 1138 344018 1803
rect 116163 1123 116229 1124
<< via4 >>
rect 1096 148388 1332 148624
rect 110658 148388 110894 148624
rect 1706 135388 1942 135624
rect 109998 135388 110234 135624
rect 1096 122388 1332 122624
rect 110658 122388 110894 122624
rect 1706 109388 1942 109624
rect 109998 109388 110234 109624
rect 1096 96388 1332 96624
rect 110658 96388 110894 96624
rect 119046 148388 119282 148624
rect 518642 148388 518878 148624
rect 119706 135388 119942 135624
rect 517982 135388 518218 135624
rect 119046 122388 119282 122624
rect 518642 122388 518878 122624
rect 119706 109388 119942 109624
rect 517982 109388 518218 109624
rect 119046 96388 119282 96624
rect 518642 96388 518878 96624
rect 1706 83388 1942 83624
rect 109998 83388 110234 83624
rect 119706 83388 119942 83624
rect 517982 83388 518218 83624
rect 1096 70388 1332 70624
rect 110658 70388 110894 70624
rect 119046 70388 119282 70624
rect 518642 70388 518878 70624
rect 1706 57388 1942 57624
rect 109998 57388 110234 57624
rect 119706 57388 119942 57624
rect 517982 57388 518218 57624
rect 1096 44388 1332 44624
rect 110658 44388 110894 44624
rect 119046 44388 119282 44624
rect 518642 44388 518878 44624
rect 1706 31388 1942 31624
rect 109998 31388 110234 31624
rect 119706 31388 119942 31624
rect 517982 31388 518218 31624
rect 1096 18388 1332 18624
rect 110658 18388 110894 18624
rect 1706 5388 1942 5624
rect 109998 5388 110234 5624
rect 119046 18388 119282 18624
rect 518642 18388 518878 18624
rect 119706 5388 119942 5624
rect 517982 5388 518218 5624
rect 164102 1052 164338 1138
rect 164102 988 164188 1052
rect 164188 988 164252 1052
rect 164252 988 164338 1052
rect 164102 902 164338 988
rect 193542 1052 193778 1138
rect 193542 988 193628 1052
rect 193628 988 193692 1052
rect 193692 988 193778 1052
rect 193542 902 193778 988
rect 231078 1052 231314 1138
rect 231078 988 231164 1052
rect 231164 988 231228 1052
rect 231228 988 231314 1052
rect 231078 902 231314 988
rect 241750 1052 241986 1138
rect 241750 988 241836 1052
rect 241836 988 241900 1052
rect 241900 988 241986 1052
rect 241750 902 241986 988
rect 343870 902 344106 1138
rect 360062 1052 360298 1138
rect 360062 988 360148 1052
rect 360148 988 360212 1052
rect 360212 988 360298 1052
rect 360062 902 360298 988
<< metal5 >>
rect 1072 148624 2200 148666
rect 1072 148388 1096 148624
rect 1332 148388 2200 148624
rect 1072 148346 2200 148388
rect 109800 148624 120200 148666
rect 109800 148388 110658 148624
rect 110894 148388 119046 148624
rect 119282 148388 120200 148624
rect 109800 148346 120200 148388
rect 517800 148624 522836 148666
rect 517800 148388 518642 148624
rect 518878 148388 522836 148624
rect 517800 148346 522836 148388
rect 1104 135624 2200 135666
rect 1104 135388 1706 135624
rect 1942 135388 2200 135624
rect 1104 135346 2200 135388
rect 109800 135624 120200 135666
rect 109800 135388 109998 135624
rect 110234 135388 119706 135624
rect 119942 135388 120200 135624
rect 109800 135346 120200 135388
rect 517800 135624 522836 135666
rect 517800 135388 517982 135624
rect 518218 135388 522836 135624
rect 517800 135346 522836 135388
rect 1072 122624 2200 122666
rect 1072 122388 1096 122624
rect 1332 122388 2200 122624
rect 1072 122346 2200 122388
rect 109800 122624 120200 122666
rect 109800 122388 110658 122624
rect 110894 122388 119046 122624
rect 119282 122388 120200 122624
rect 109800 122346 120200 122388
rect 517800 122624 522836 122666
rect 517800 122388 518642 122624
rect 518878 122388 522836 122624
rect 517800 122346 522836 122388
rect 1104 109624 2200 109666
rect 1104 109388 1706 109624
rect 1942 109388 2200 109624
rect 1104 109346 2200 109388
rect 109800 109624 120200 109666
rect 109800 109388 109998 109624
rect 110234 109388 119706 109624
rect 119942 109388 120200 109624
rect 109800 109346 120200 109388
rect 517800 109624 522836 109666
rect 517800 109388 517982 109624
rect 518218 109388 522836 109624
rect 517800 109346 522836 109388
rect 1072 96624 2200 96666
rect 1072 96388 1096 96624
rect 1332 96388 2200 96624
rect 1072 96346 2200 96388
rect 109800 96624 120200 96666
rect 109800 96388 110658 96624
rect 110894 96388 119046 96624
rect 119282 96388 120200 96624
rect 109800 96346 120200 96388
rect 517800 96624 522836 96666
rect 517800 96388 518642 96624
rect 518878 96388 522836 96624
rect 517800 96346 522836 96388
rect 1104 83624 2200 83666
rect 1104 83388 1706 83624
rect 1942 83388 2200 83624
rect 1104 83346 2200 83388
rect 109800 83624 120200 83666
rect 109800 83388 109998 83624
rect 110234 83388 119706 83624
rect 119942 83388 120200 83624
rect 109800 83346 120200 83388
rect 517800 83624 522836 83666
rect 517800 83388 517982 83624
rect 518218 83388 522836 83624
rect 517800 83346 522836 83388
rect 1072 70624 2200 70666
rect 1072 70388 1096 70624
rect 1332 70388 2200 70624
rect 1072 70346 2200 70388
rect 109800 70624 120200 70666
rect 109800 70388 110658 70624
rect 110894 70388 119046 70624
rect 119282 70388 120200 70624
rect 109800 70346 120200 70388
rect 517800 70624 522836 70666
rect 517800 70388 518642 70624
rect 518878 70388 522836 70624
rect 517800 70346 522836 70388
rect 1104 57624 2200 57666
rect 1104 57388 1706 57624
rect 1942 57388 2200 57624
rect 1104 57346 2200 57388
rect 109800 57624 120200 57666
rect 109800 57388 109998 57624
rect 110234 57388 119706 57624
rect 119942 57388 120200 57624
rect 109800 57346 120200 57388
rect 517800 57624 522836 57666
rect 517800 57388 517982 57624
rect 518218 57388 522836 57624
rect 517800 57346 522836 57388
rect 1072 44624 2200 44666
rect 1072 44388 1096 44624
rect 1332 44388 2200 44624
rect 1072 44346 2200 44388
rect 109800 44624 120200 44666
rect 109800 44388 110658 44624
rect 110894 44388 119046 44624
rect 119282 44388 120200 44624
rect 109800 44346 120200 44388
rect 517800 44624 522836 44666
rect 517800 44388 518642 44624
rect 518878 44388 522836 44624
rect 517800 44346 522836 44388
rect 1104 31624 2200 31666
rect 1104 31388 1706 31624
rect 1942 31388 2200 31624
rect 1104 31346 2200 31388
rect 109800 31624 120200 31666
rect 109800 31388 109998 31624
rect 110234 31388 119706 31624
rect 119942 31388 120200 31624
rect 109800 31346 120200 31388
rect 517800 31624 522836 31666
rect 517800 31388 517982 31624
rect 518218 31388 522836 31624
rect 517800 31346 522836 31388
rect 1072 18624 2200 18666
rect 1072 18388 1096 18624
rect 1332 18388 2200 18624
rect 1072 18346 2200 18388
rect 109800 18624 120200 18666
rect 109800 18388 110658 18624
rect 110894 18388 119046 18624
rect 119282 18388 120200 18624
rect 109800 18346 120200 18388
rect 517800 18624 522836 18666
rect 517800 18388 518642 18624
rect 518878 18388 522836 18624
rect 517800 18346 522836 18388
rect 1104 5624 2200 5666
rect 1104 5388 1706 5624
rect 1942 5388 2200 5624
rect 1104 5346 2200 5388
rect 109800 5624 120200 5666
rect 109800 5388 109998 5624
rect 110234 5388 119706 5624
rect 119942 5388 120200 5624
rect 109800 5346 120200 5388
rect 517800 5624 522836 5666
rect 517800 5388 517982 5624
rect 518218 5388 522836 5624
rect 517800 5346 522836 5388
rect 183196 1220 184252 1540
rect 183196 1180 183516 1220
rect 164060 1138 183516 1180
rect 164060 902 164102 1138
rect 164338 902 183516 1138
rect 164060 860 183516 902
rect 183932 1180 184252 1220
rect 192764 1220 193820 1540
rect 192764 1180 193084 1220
rect 183932 860 193084 1180
rect 193500 1138 193820 1220
rect 193500 902 193542 1138
rect 193778 902 193820 1138
rect 193500 860 193820 902
rect 231036 1220 232000 1540
rect 231036 1138 231356 1220
rect 231036 902 231078 1138
rect 231314 902 231356 1138
rect 231036 860 231356 902
rect 231680 1180 232000 1220
rect 240972 1220 242028 1540
rect 240972 1180 241292 1220
rect 231680 860 241292 1180
rect 241708 1138 242028 1220
rect 241708 902 241750 1138
rect 241986 902 242028 1138
rect 241708 860 242028 902
rect 343828 1138 360340 1180
rect 343828 902 343870 1138
rect 344106 902 360062 1138
rect 360298 902 360340 1138
rect 343828 860 360340 902
use mgmt_core  core
timestamp 1637253870
transform 1 0 119000 0 1 2000
box 0 0 400000 148000
use DFFRAM  DFFRAM
timestamp 1637253870
transform 1 0 1000 0 1 2000
box 4 0 110000 148000
<< labels >>
rlabel metal5 s 1104 18346 2200 18666 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 18346 120200 18666 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 18346 522836 18666 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 44346 2200 44666 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 44346 120200 44666 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 44346 522836 44666 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 70346 2200 70666 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 70346 120200 70666 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 70346 522836 70666 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 96346 2200 96666 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 96346 120200 96666 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 96346 522836 96666 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 122346 2200 122666 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 122346 120200 122666 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 122346 522836 122666 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 148346 2200 148666 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 148346 120200 148666 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 148346 522836 148666 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 5346 2200 5666 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 5346 120200 5666 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 5346 522836 5666 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 31346 2200 31666 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 31346 120200 31666 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 31346 522836 31666 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 57346 2200 57666 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 57346 120200 57666 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 57346 522836 57666 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 83346 2200 83666 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 83346 120200 83666 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 83346 522836 83666 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 109346 2200 109666 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 109346 120200 109666 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 109346 522836 109666 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 135346 2200 135666 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 135346 120200 135666 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 135346 522836 135666 6 VPWR
port 1 nsew power input
rlabel metal2 s 294786 -400 294842 800 6 core_clk
port 2 nsew signal input
rlabel metal2 s 98274 -400 98330 800 6 core_rstn
port 3 nsew signal input
rlabel metal3 s 523200 64472 524400 64592 6 debug_in
port 4 nsew signal input
rlabel metal3 s 523200 65968 524400 66088 6 debug_mode
port 5 nsew signal tristate
rlabel metal3 s 523200 67464 524400 67584 6 debug_oeb
port 6 nsew signal tristate
rlabel metal3 s 523200 68960 524400 69080 6 debug_out
port 7 nsew signal tristate
rlabel metal3 s 523200 144848 524400 144968 6 flash_clk
port 8 nsew signal tristate
rlabel metal3 s 523200 143352 524400 143472 6 flash_csb
port 9 nsew signal tristate
rlabel metal3 s 523200 146480 524400 146600 6 flash_io0_di
port 10 nsew signal input
rlabel metal3 s 523200 147976 524400 148096 6 flash_io0_do
port 11 nsew signal tristate
rlabel metal3 s 523200 149472 524400 149592 6 flash_io0_oeb
port 12 nsew signal tristate
rlabel metal3 s 523200 150968 524400 151088 6 flash_io1_di
port 13 nsew signal input
rlabel metal3 s 523200 152464 524400 152584 6 flash_io1_do
port 14 nsew signal tristate
rlabel metal3 s 523200 153960 524400 154080 6 flash_io1_oeb
port 15 nsew signal tristate
rlabel metal3 s 523200 155592 524400 155712 6 flash_io2_di
port 16 nsew signal input
rlabel metal3 s 523200 157088 524400 157208 6 flash_io2_do
port 17 nsew signal tristate
rlabel metal3 s 523200 158584 524400 158704 6 flash_io2_oeb
port 18 nsew signal tristate
rlabel metal3 s 523200 160080 524400 160200 6 flash_io3_di
port 19 nsew signal input
rlabel metal3 s 523200 161576 524400 161696 6 flash_io3_do
port 20 nsew signal tristate
rlabel metal3 s 523200 163072 524400 163192 6 flash_io3_oeb
port 21 nsew signal tristate
rlabel metal2 s 32770 -400 32826 800 6 gpio_in_pad
port 22 nsew signal input
rlabel metal2 s 163778 -400 163834 800 6 gpio_inenb_pad
port 23 nsew signal tristate
rlabel metal2 s 229282 -400 229338 800 6 gpio_mode0_pad
port 24 nsew signal tristate
rlabel metal2 s 360290 -400 360346 800 6 gpio_mode1_pad
port 25 nsew signal tristate
rlabel metal2 s 425794 -400 425850 800 6 gpio_out_pad
port 26 nsew signal tristate
rlabel metal2 s 491298 -400 491354 800 6 gpio_outenb_pad
port 27 nsew signal tristate
rlabel metal3 s 523200 91808 524400 91928 6 hk_ack_i
port 28 nsew signal input
rlabel metal3 s 523200 94800 524400 94920 6 hk_dat_i[0]
port 29 nsew signal input
rlabel metal3 s 523200 110032 524400 110152 6 hk_dat_i[10]
port 30 nsew signal input
rlabel metal3 s 523200 111528 524400 111648 6 hk_dat_i[11]
port 31 nsew signal input
rlabel metal3 s 523200 113024 524400 113144 6 hk_dat_i[12]
port 32 nsew signal input
rlabel metal3 s 523200 114520 524400 114640 6 hk_dat_i[13]
port 33 nsew signal input
rlabel metal3 s 523200 116016 524400 116136 6 hk_dat_i[14]
port 34 nsew signal input
rlabel metal3 s 523200 117512 524400 117632 6 hk_dat_i[15]
port 35 nsew signal input
rlabel metal3 s 523200 119144 524400 119264 6 hk_dat_i[16]
port 36 nsew signal input
rlabel metal3 s 523200 120640 524400 120760 6 hk_dat_i[17]
port 37 nsew signal input
rlabel metal3 s 523200 122136 524400 122256 6 hk_dat_i[18]
port 38 nsew signal input
rlabel metal3 s 523200 123632 524400 123752 6 hk_dat_i[19]
port 39 nsew signal input
rlabel metal3 s 523200 96296 524400 96416 6 hk_dat_i[1]
port 40 nsew signal input
rlabel metal3 s 523200 125128 524400 125248 6 hk_dat_i[20]
port 41 nsew signal input
rlabel metal3 s 523200 126624 524400 126744 6 hk_dat_i[21]
port 42 nsew signal input
rlabel metal3 s 523200 128256 524400 128376 6 hk_dat_i[22]
port 43 nsew signal input
rlabel metal3 s 523200 129752 524400 129872 6 hk_dat_i[23]
port 44 nsew signal input
rlabel metal3 s 523200 131248 524400 131368 6 hk_dat_i[24]
port 45 nsew signal input
rlabel metal3 s 523200 132744 524400 132864 6 hk_dat_i[25]
port 46 nsew signal input
rlabel metal3 s 523200 134240 524400 134360 6 hk_dat_i[26]
port 47 nsew signal input
rlabel metal3 s 523200 135736 524400 135856 6 hk_dat_i[27]
port 48 nsew signal input
rlabel metal3 s 523200 137368 524400 137488 6 hk_dat_i[28]
port 49 nsew signal input
rlabel metal3 s 523200 138864 524400 138984 6 hk_dat_i[29]
port 50 nsew signal input
rlabel metal3 s 523200 97792 524400 97912 6 hk_dat_i[2]
port 51 nsew signal input
rlabel metal3 s 523200 140360 524400 140480 6 hk_dat_i[30]
port 52 nsew signal input
rlabel metal3 s 523200 141856 524400 141976 6 hk_dat_i[31]
port 53 nsew signal input
rlabel metal3 s 523200 99288 524400 99408 6 hk_dat_i[3]
port 54 nsew signal input
rlabel metal3 s 523200 100920 524400 101040 6 hk_dat_i[4]
port 55 nsew signal input
rlabel metal3 s 523200 102416 524400 102536 6 hk_dat_i[5]
port 56 nsew signal input
rlabel metal3 s 523200 103912 524400 104032 6 hk_dat_i[6]
port 57 nsew signal input
rlabel metal3 s 523200 105408 524400 105528 6 hk_dat_i[7]
port 58 nsew signal input
rlabel metal3 s 523200 106904 524400 107024 6 hk_dat_i[8]
port 59 nsew signal input
rlabel metal3 s 523200 108400 524400 108520 6 hk_dat_i[9]
port 60 nsew signal input
rlabel metal3 s 523200 93304 524400 93424 6 hk_stb_o
port 61 nsew signal tristate
rlabel metal2 s 521842 163200 521898 164400 6 irq[0]
port 62 nsew signal input
rlabel metal2 s 522670 163200 522726 164400 6 irq[1]
port 63 nsew signal input
rlabel metal2 s 523498 163200 523554 164400 6 irq[2]
port 64 nsew signal input
rlabel metal3 s 523200 75080 524400 75200 6 irq[3]
port 65 nsew signal input
rlabel metal3 s 523200 73584 524400 73704 6 irq[4]
port 66 nsew signal input
rlabel metal3 s 523200 71952 524400 72072 6 irq[5]
port 67 nsew signal input
rlabel metal2 s 386 163200 442 164400 6 la_iena[0]
port 68 nsew signal tristate
rlabel metal2 s 336830 163200 336886 164400 6 la_iena[100]
port 69 nsew signal tristate
rlabel metal2 s 340142 163200 340198 164400 6 la_iena[101]
port 70 nsew signal tristate
rlabel metal2 s 343546 163200 343602 164400 6 la_iena[102]
port 71 nsew signal tristate
rlabel metal2 s 346858 163200 346914 164400 6 la_iena[103]
port 72 nsew signal tristate
rlabel metal2 s 350262 163200 350318 164400 6 la_iena[104]
port 73 nsew signal tristate
rlabel metal2 s 353666 163200 353722 164400 6 la_iena[105]
port 74 nsew signal tristate
rlabel metal2 s 356978 163200 357034 164400 6 la_iena[106]
port 75 nsew signal tristate
rlabel metal2 s 360382 163200 360438 164400 6 la_iena[107]
port 76 nsew signal tristate
rlabel metal2 s 363694 163200 363750 164400 6 la_iena[108]
port 77 nsew signal tristate
rlabel metal2 s 367098 163200 367154 164400 6 la_iena[109]
port 78 nsew signal tristate
rlabel metal2 s 33966 163200 34022 164400 6 la_iena[10]
port 79 nsew signal tristate
rlabel metal2 s 370410 163200 370466 164400 6 la_iena[110]
port 80 nsew signal tristate
rlabel metal2 s 373814 163200 373870 164400 6 la_iena[111]
port 81 nsew signal tristate
rlabel metal2 s 377218 163200 377274 164400 6 la_iena[112]
port 82 nsew signal tristate
rlabel metal2 s 380530 163200 380586 164400 6 la_iena[113]
port 83 nsew signal tristate
rlabel metal2 s 383934 163200 383990 164400 6 la_iena[114]
port 84 nsew signal tristate
rlabel metal2 s 387246 163200 387302 164400 6 la_iena[115]
port 85 nsew signal tristate
rlabel metal2 s 390650 163200 390706 164400 6 la_iena[116]
port 86 nsew signal tristate
rlabel metal2 s 393962 163200 394018 164400 6 la_iena[117]
port 87 nsew signal tristate
rlabel metal2 s 397366 163200 397422 164400 6 la_iena[118]
port 88 nsew signal tristate
rlabel metal2 s 400770 163200 400826 164400 6 la_iena[119]
port 89 nsew signal tristate
rlabel metal2 s 37370 163200 37426 164400 6 la_iena[11]
port 90 nsew signal tristate
rlabel metal2 s 404082 163200 404138 164400 6 la_iena[120]
port 91 nsew signal tristate
rlabel metal2 s 407486 163200 407542 164400 6 la_iena[121]
port 92 nsew signal tristate
rlabel metal2 s 410798 163200 410854 164400 6 la_iena[122]
port 93 nsew signal tristate
rlabel metal2 s 414202 163200 414258 164400 6 la_iena[123]
port 94 nsew signal tristate
rlabel metal2 s 417514 163200 417570 164400 6 la_iena[124]
port 95 nsew signal tristate
rlabel metal2 s 420918 163200 420974 164400 6 la_iena[125]
port 96 nsew signal tristate
rlabel metal2 s 424322 163200 424378 164400 6 la_iena[126]
port 97 nsew signal tristate
rlabel metal2 s 427634 163200 427690 164400 6 la_iena[127]
port 98 nsew signal tristate
rlabel metal2 s 40682 163200 40738 164400 6 la_iena[12]
port 99 nsew signal tristate
rlabel metal2 s 44086 163200 44142 164400 6 la_iena[13]
port 100 nsew signal tristate
rlabel metal2 s 47490 163200 47546 164400 6 la_iena[14]
port 101 nsew signal tristate
rlabel metal2 s 50802 163200 50858 164400 6 la_iena[15]
port 102 nsew signal tristate
rlabel metal2 s 54206 163200 54262 164400 6 la_iena[16]
port 103 nsew signal tristate
rlabel metal2 s 57518 163200 57574 164400 6 la_iena[17]
port 104 nsew signal tristate
rlabel metal2 s 60922 163200 60978 164400 6 la_iena[18]
port 105 nsew signal tristate
rlabel metal2 s 64234 163200 64290 164400 6 la_iena[19]
port 106 nsew signal tristate
rlabel metal2 s 3698 163200 3754 164400 6 la_iena[1]
port 107 nsew signal tristate
rlabel metal2 s 67638 163200 67694 164400 6 la_iena[20]
port 108 nsew signal tristate
rlabel metal2 s 71042 163200 71098 164400 6 la_iena[21]
port 109 nsew signal tristate
rlabel metal2 s 74354 163200 74410 164400 6 la_iena[22]
port 110 nsew signal tristate
rlabel metal2 s 77758 163200 77814 164400 6 la_iena[23]
port 111 nsew signal tristate
rlabel metal2 s 81070 163200 81126 164400 6 la_iena[24]
port 112 nsew signal tristate
rlabel metal2 s 84474 163200 84530 164400 6 la_iena[25]
port 113 nsew signal tristate
rlabel metal2 s 87786 163200 87842 164400 6 la_iena[26]
port 114 nsew signal tristate
rlabel metal2 s 91190 163200 91246 164400 6 la_iena[27]
port 115 nsew signal tristate
rlabel metal2 s 94594 163200 94650 164400 6 la_iena[28]
port 116 nsew signal tristate
rlabel metal2 s 97906 163200 97962 164400 6 la_iena[29]
port 117 nsew signal tristate
rlabel metal2 s 7102 163200 7158 164400 6 la_iena[2]
port 118 nsew signal tristate
rlabel metal2 s 101310 163200 101366 164400 6 la_iena[30]
port 119 nsew signal tristate
rlabel metal2 s 104622 163200 104678 164400 6 la_iena[31]
port 120 nsew signal tristate
rlabel metal2 s 108026 163200 108082 164400 6 la_iena[32]
port 121 nsew signal tristate
rlabel metal2 s 111338 163200 111394 164400 6 la_iena[33]
port 122 nsew signal tristate
rlabel metal2 s 114742 163200 114798 164400 6 la_iena[34]
port 123 nsew signal tristate
rlabel metal2 s 118146 163200 118202 164400 6 la_iena[35]
port 124 nsew signal tristate
rlabel metal2 s 121458 163200 121514 164400 6 la_iena[36]
port 125 nsew signal tristate
rlabel metal2 s 124862 163200 124918 164400 6 la_iena[37]
port 126 nsew signal tristate
rlabel metal2 s 128174 163200 128230 164400 6 la_iena[38]
port 127 nsew signal tristate
rlabel metal2 s 131578 163200 131634 164400 6 la_iena[39]
port 128 nsew signal tristate
rlabel metal2 s 10414 163200 10470 164400 6 la_iena[3]
port 129 nsew signal tristate
rlabel metal2 s 134890 163200 134946 164400 6 la_iena[40]
port 130 nsew signal tristate
rlabel metal2 s 138294 163200 138350 164400 6 la_iena[41]
port 131 nsew signal tristate
rlabel metal2 s 141698 163200 141754 164400 6 la_iena[42]
port 132 nsew signal tristate
rlabel metal2 s 145010 163200 145066 164400 6 la_iena[43]
port 133 nsew signal tristate
rlabel metal2 s 148414 163200 148470 164400 6 la_iena[44]
port 134 nsew signal tristate
rlabel metal2 s 151726 163200 151782 164400 6 la_iena[45]
port 135 nsew signal tristate
rlabel metal2 s 155130 163200 155186 164400 6 la_iena[46]
port 136 nsew signal tristate
rlabel metal2 s 158442 163200 158498 164400 6 la_iena[47]
port 137 nsew signal tristate
rlabel metal2 s 161846 163200 161902 164400 6 la_iena[48]
port 138 nsew signal tristate
rlabel metal2 s 165250 163200 165306 164400 6 la_iena[49]
port 139 nsew signal tristate
rlabel metal2 s 13818 163200 13874 164400 6 la_iena[4]
port 140 nsew signal tristate
rlabel metal2 s 168562 163200 168618 164400 6 la_iena[50]
port 141 nsew signal tristate
rlabel metal2 s 171966 163200 172022 164400 6 la_iena[51]
port 142 nsew signal tristate
rlabel metal2 s 175278 163200 175334 164400 6 la_iena[52]
port 143 nsew signal tristate
rlabel metal2 s 178682 163200 178738 164400 6 la_iena[53]
port 144 nsew signal tristate
rlabel metal2 s 181994 163200 182050 164400 6 la_iena[54]
port 145 nsew signal tristate
rlabel metal2 s 185398 163200 185454 164400 6 la_iena[55]
port 146 nsew signal tristate
rlabel metal2 s 188802 163200 188858 164400 6 la_iena[56]
port 147 nsew signal tristate
rlabel metal2 s 192114 163200 192170 164400 6 la_iena[57]
port 148 nsew signal tristate
rlabel metal2 s 195518 163200 195574 164400 6 la_iena[58]
port 149 nsew signal tristate
rlabel metal2 s 198830 163200 198886 164400 6 la_iena[59]
port 150 nsew signal tristate
rlabel metal2 s 17130 163200 17186 164400 6 la_iena[5]
port 151 nsew signal tristate
rlabel metal2 s 202234 163200 202290 164400 6 la_iena[60]
port 152 nsew signal tristate
rlabel metal2 s 205546 163200 205602 164400 6 la_iena[61]
port 153 nsew signal tristate
rlabel metal2 s 208950 163200 209006 164400 6 la_iena[62]
port 154 nsew signal tristate
rlabel metal2 s 212354 163200 212410 164400 6 la_iena[63]
port 155 nsew signal tristate
rlabel metal2 s 215666 163200 215722 164400 6 la_iena[64]
port 156 nsew signal tristate
rlabel metal2 s 219070 163200 219126 164400 6 la_iena[65]
port 157 nsew signal tristate
rlabel metal2 s 222382 163200 222438 164400 6 la_iena[66]
port 158 nsew signal tristate
rlabel metal2 s 225786 163200 225842 164400 6 la_iena[67]
port 159 nsew signal tristate
rlabel metal2 s 229098 163200 229154 164400 6 la_iena[68]
port 160 nsew signal tristate
rlabel metal2 s 232502 163200 232558 164400 6 la_iena[69]
port 161 nsew signal tristate
rlabel metal2 s 20534 163200 20590 164400 6 la_iena[6]
port 162 nsew signal tristate
rlabel metal2 s 235906 163200 235962 164400 6 la_iena[70]
port 163 nsew signal tristate
rlabel metal2 s 239218 163200 239274 164400 6 la_iena[71]
port 164 nsew signal tristate
rlabel metal2 s 242622 163200 242678 164400 6 la_iena[72]
port 165 nsew signal tristate
rlabel metal2 s 245934 163200 245990 164400 6 la_iena[73]
port 166 nsew signal tristate
rlabel metal2 s 249338 163200 249394 164400 6 la_iena[74]
port 167 nsew signal tristate
rlabel metal2 s 252650 163200 252706 164400 6 la_iena[75]
port 168 nsew signal tristate
rlabel metal2 s 256054 163200 256110 164400 6 la_iena[76]
port 169 nsew signal tristate
rlabel metal2 s 259458 163200 259514 164400 6 la_iena[77]
port 170 nsew signal tristate
rlabel metal2 s 262770 163200 262826 164400 6 la_iena[78]
port 171 nsew signal tristate
rlabel metal2 s 266174 163200 266230 164400 6 la_iena[79]
port 172 nsew signal tristate
rlabel metal2 s 23938 163200 23994 164400 6 la_iena[7]
port 173 nsew signal tristate
rlabel metal2 s 269486 163200 269542 164400 6 la_iena[80]
port 174 nsew signal tristate
rlabel metal2 s 272890 163200 272946 164400 6 la_iena[81]
port 175 nsew signal tristate
rlabel metal2 s 276202 163200 276258 164400 6 la_iena[82]
port 176 nsew signal tristate
rlabel metal2 s 279606 163200 279662 164400 6 la_iena[83]
port 177 nsew signal tristate
rlabel metal2 s 283010 163200 283066 164400 6 la_iena[84]
port 178 nsew signal tristate
rlabel metal2 s 286322 163200 286378 164400 6 la_iena[85]
port 179 nsew signal tristate
rlabel metal2 s 289726 163200 289782 164400 6 la_iena[86]
port 180 nsew signal tristate
rlabel metal2 s 293038 163200 293094 164400 6 la_iena[87]
port 181 nsew signal tristate
rlabel metal2 s 296442 163200 296498 164400 6 la_iena[88]
port 182 nsew signal tristate
rlabel metal2 s 299754 163200 299810 164400 6 la_iena[89]
port 183 nsew signal tristate
rlabel metal2 s 27250 163200 27306 164400 6 la_iena[8]
port 184 nsew signal tristate
rlabel metal2 s 303158 163200 303214 164400 6 la_iena[90]
port 185 nsew signal tristate
rlabel metal2 s 306562 163200 306618 164400 6 la_iena[91]
port 186 nsew signal tristate
rlabel metal2 s 309874 163200 309930 164400 6 la_iena[92]
port 187 nsew signal tristate
rlabel metal2 s 313278 163200 313334 164400 6 la_iena[93]
port 188 nsew signal tristate
rlabel metal2 s 316590 163200 316646 164400 6 la_iena[94]
port 189 nsew signal tristate
rlabel metal2 s 319994 163200 320050 164400 6 la_iena[95]
port 190 nsew signal tristate
rlabel metal2 s 323306 163200 323362 164400 6 la_iena[96]
port 191 nsew signal tristate
rlabel metal2 s 326710 163200 326766 164400 6 la_iena[97]
port 192 nsew signal tristate
rlabel metal2 s 330114 163200 330170 164400 6 la_iena[98]
port 193 nsew signal tristate
rlabel metal2 s 333426 163200 333482 164400 6 la_iena[99]
port 194 nsew signal tristate
rlabel metal2 s 30654 163200 30710 164400 6 la_iena[9]
port 195 nsew signal tristate
rlabel metal2 s 1214 163200 1270 164400 6 la_input[0]
port 196 nsew signal input
rlabel metal2 s 337658 163200 337714 164400 6 la_input[100]
port 197 nsew signal input
rlabel metal2 s 340970 163200 341026 164400 6 la_input[101]
port 198 nsew signal input
rlabel metal2 s 344374 163200 344430 164400 6 la_input[102]
port 199 nsew signal input
rlabel metal2 s 347778 163200 347834 164400 6 la_input[103]
port 200 nsew signal input
rlabel metal2 s 351090 163200 351146 164400 6 la_input[104]
port 201 nsew signal input
rlabel metal2 s 354494 163200 354550 164400 6 la_input[105]
port 202 nsew signal input
rlabel metal2 s 357806 163200 357862 164400 6 la_input[106]
port 203 nsew signal input
rlabel metal2 s 361210 163200 361266 164400 6 la_input[107]
port 204 nsew signal input
rlabel metal2 s 364522 163200 364578 164400 6 la_input[108]
port 205 nsew signal input
rlabel metal2 s 367926 163200 367982 164400 6 la_input[109]
port 206 nsew signal input
rlabel metal2 s 34794 163200 34850 164400 6 la_input[10]
port 207 nsew signal input
rlabel metal2 s 371330 163200 371386 164400 6 la_input[110]
port 208 nsew signal input
rlabel metal2 s 374642 163200 374698 164400 6 la_input[111]
port 209 nsew signal input
rlabel metal2 s 378046 163200 378102 164400 6 la_input[112]
port 210 nsew signal input
rlabel metal2 s 381358 163200 381414 164400 6 la_input[113]
port 211 nsew signal input
rlabel metal2 s 384762 163200 384818 164400 6 la_input[114]
port 212 nsew signal input
rlabel metal2 s 388074 163200 388130 164400 6 la_input[115]
port 213 nsew signal input
rlabel metal2 s 391478 163200 391534 164400 6 la_input[116]
port 214 nsew signal input
rlabel metal2 s 394882 163200 394938 164400 6 la_input[117]
port 215 nsew signal input
rlabel metal2 s 398194 163200 398250 164400 6 la_input[118]
port 216 nsew signal input
rlabel metal2 s 401598 163200 401654 164400 6 la_input[119]
port 217 nsew signal input
rlabel metal2 s 38198 163200 38254 164400 6 la_input[11]
port 218 nsew signal input
rlabel metal2 s 404910 163200 404966 164400 6 la_input[120]
port 219 nsew signal input
rlabel metal2 s 408314 163200 408370 164400 6 la_input[121]
port 220 nsew signal input
rlabel metal2 s 411626 163200 411682 164400 6 la_input[122]
port 221 nsew signal input
rlabel metal2 s 415030 163200 415086 164400 6 la_input[123]
port 222 nsew signal input
rlabel metal2 s 418434 163200 418490 164400 6 la_input[124]
port 223 nsew signal input
rlabel metal2 s 421746 163200 421802 164400 6 la_input[125]
port 224 nsew signal input
rlabel metal2 s 425150 163200 425206 164400 6 la_input[126]
port 225 nsew signal input
rlabel metal2 s 428462 163200 428518 164400 6 la_input[127]
port 226 nsew signal input
rlabel metal2 s 41602 163200 41658 164400 6 la_input[12]
port 227 nsew signal input
rlabel metal2 s 44914 163200 44970 164400 6 la_input[13]
port 228 nsew signal input
rlabel metal2 s 48318 163200 48374 164400 6 la_input[14]
port 229 nsew signal input
rlabel metal2 s 51630 163200 51686 164400 6 la_input[15]
port 230 nsew signal input
rlabel metal2 s 55034 163200 55090 164400 6 la_input[16]
port 231 nsew signal input
rlabel metal2 s 58346 163200 58402 164400 6 la_input[17]
port 232 nsew signal input
rlabel metal2 s 61750 163200 61806 164400 6 la_input[18]
port 233 nsew signal input
rlabel metal2 s 65154 163200 65210 164400 6 la_input[19]
port 234 nsew signal input
rlabel metal2 s 4526 163200 4582 164400 6 la_input[1]
port 235 nsew signal input
rlabel metal2 s 68466 163200 68522 164400 6 la_input[20]
port 236 nsew signal input
rlabel metal2 s 71870 163200 71926 164400 6 la_input[21]
port 237 nsew signal input
rlabel metal2 s 75182 163200 75238 164400 6 la_input[22]
port 238 nsew signal input
rlabel metal2 s 78586 163200 78642 164400 6 la_input[23]
port 239 nsew signal input
rlabel metal2 s 81898 163200 81954 164400 6 la_input[24]
port 240 nsew signal input
rlabel metal2 s 85302 163200 85358 164400 6 la_input[25]
port 241 nsew signal input
rlabel metal2 s 88706 163200 88762 164400 6 la_input[26]
port 242 nsew signal input
rlabel metal2 s 92018 163200 92074 164400 6 la_input[27]
port 243 nsew signal input
rlabel metal2 s 95422 163200 95478 164400 6 la_input[28]
port 244 nsew signal input
rlabel metal2 s 98734 163200 98790 164400 6 la_input[29]
port 245 nsew signal input
rlabel metal2 s 7930 163200 7986 164400 6 la_input[2]
port 246 nsew signal input
rlabel metal2 s 102138 163200 102194 164400 6 la_input[30]
port 247 nsew signal input
rlabel metal2 s 105450 163200 105506 164400 6 la_input[31]
port 248 nsew signal input
rlabel metal2 s 108854 163200 108910 164400 6 la_input[32]
port 249 nsew signal input
rlabel metal2 s 112258 163200 112314 164400 6 la_input[33]
port 250 nsew signal input
rlabel metal2 s 115570 163200 115626 164400 6 la_input[34]
port 251 nsew signal input
rlabel metal2 s 118974 163200 119030 164400 6 la_input[35]
port 252 nsew signal input
rlabel metal2 s 122286 163200 122342 164400 6 la_input[36]
port 253 nsew signal input
rlabel metal2 s 125690 163200 125746 164400 6 la_input[37]
port 254 nsew signal input
rlabel metal2 s 129002 163200 129058 164400 6 la_input[38]
port 255 nsew signal input
rlabel metal2 s 132406 163200 132462 164400 6 la_input[39]
port 256 nsew signal input
rlabel metal2 s 11242 163200 11298 164400 6 la_input[3]
port 257 nsew signal input
rlabel metal2 s 135810 163200 135866 164400 6 la_input[40]
port 258 nsew signal input
rlabel metal2 s 139122 163200 139178 164400 6 la_input[41]
port 259 nsew signal input
rlabel metal2 s 142526 163200 142582 164400 6 la_input[42]
port 260 nsew signal input
rlabel metal2 s 145838 163200 145894 164400 6 la_input[43]
port 261 nsew signal input
rlabel metal2 s 149242 163200 149298 164400 6 la_input[44]
port 262 nsew signal input
rlabel metal2 s 152554 163200 152610 164400 6 la_input[45]
port 263 nsew signal input
rlabel metal2 s 155958 163200 156014 164400 6 la_input[46]
port 264 nsew signal input
rlabel metal2 s 159362 163200 159418 164400 6 la_input[47]
port 265 nsew signal input
rlabel metal2 s 162674 163200 162730 164400 6 la_input[48]
port 266 nsew signal input
rlabel metal2 s 166078 163200 166134 164400 6 la_input[49]
port 267 nsew signal input
rlabel metal2 s 14646 163200 14702 164400 6 la_input[4]
port 268 nsew signal input
rlabel metal2 s 169390 163200 169446 164400 6 la_input[50]
port 269 nsew signal input
rlabel metal2 s 172794 163200 172850 164400 6 la_input[51]
port 270 nsew signal input
rlabel metal2 s 176106 163200 176162 164400 6 la_input[52]
port 271 nsew signal input
rlabel metal2 s 179510 163200 179566 164400 6 la_input[53]
port 272 nsew signal input
rlabel metal2 s 182914 163200 182970 164400 6 la_input[54]
port 273 nsew signal input
rlabel metal2 s 186226 163200 186282 164400 6 la_input[55]
port 274 nsew signal input
rlabel metal2 s 189630 163200 189686 164400 6 la_input[56]
port 275 nsew signal input
rlabel metal2 s 192942 163200 192998 164400 6 la_input[57]
port 276 nsew signal input
rlabel metal2 s 196346 163200 196402 164400 6 la_input[58]
port 277 nsew signal input
rlabel metal2 s 199658 163200 199714 164400 6 la_input[59]
port 278 nsew signal input
rlabel metal2 s 18050 163200 18106 164400 6 la_input[5]
port 279 nsew signal input
rlabel metal2 s 203062 163200 203118 164400 6 la_input[60]
port 280 nsew signal input
rlabel metal2 s 206466 163200 206522 164400 6 la_input[61]
port 281 nsew signal input
rlabel metal2 s 209778 163200 209834 164400 6 la_input[62]
port 282 nsew signal input
rlabel metal2 s 213182 163200 213238 164400 6 la_input[63]
port 283 nsew signal input
rlabel metal2 s 216494 163200 216550 164400 6 la_input[64]
port 284 nsew signal input
rlabel metal2 s 219898 163200 219954 164400 6 la_input[65]
port 285 nsew signal input
rlabel metal2 s 223210 163200 223266 164400 6 la_input[66]
port 286 nsew signal input
rlabel metal2 s 226614 163200 226670 164400 6 la_input[67]
port 287 nsew signal input
rlabel metal2 s 230018 163200 230074 164400 6 la_input[68]
port 288 nsew signal input
rlabel metal2 s 233330 163200 233386 164400 6 la_input[69]
port 289 nsew signal input
rlabel metal2 s 21362 163200 21418 164400 6 la_input[6]
port 290 nsew signal input
rlabel metal2 s 236734 163200 236790 164400 6 la_input[70]
port 291 nsew signal input
rlabel metal2 s 240046 163200 240102 164400 6 la_input[71]
port 292 nsew signal input
rlabel metal2 s 243450 163200 243506 164400 6 la_input[72]
port 293 nsew signal input
rlabel metal2 s 246762 163200 246818 164400 6 la_input[73]
port 294 nsew signal input
rlabel metal2 s 250166 163200 250222 164400 6 la_input[74]
port 295 nsew signal input
rlabel metal2 s 253570 163200 253626 164400 6 la_input[75]
port 296 nsew signal input
rlabel metal2 s 256882 163200 256938 164400 6 la_input[76]
port 297 nsew signal input
rlabel metal2 s 260286 163200 260342 164400 6 la_input[77]
port 298 nsew signal input
rlabel metal2 s 263598 163200 263654 164400 6 la_input[78]
port 299 nsew signal input
rlabel metal2 s 267002 163200 267058 164400 6 la_input[79]
port 300 nsew signal input
rlabel metal2 s 24766 163200 24822 164400 6 la_input[7]
port 301 nsew signal input
rlabel metal2 s 270314 163200 270370 164400 6 la_input[80]
port 302 nsew signal input
rlabel metal2 s 273718 163200 273774 164400 6 la_input[81]
port 303 nsew signal input
rlabel metal2 s 277122 163200 277178 164400 6 la_input[82]
port 304 nsew signal input
rlabel metal2 s 280434 163200 280490 164400 6 la_input[83]
port 305 nsew signal input
rlabel metal2 s 283838 163200 283894 164400 6 la_input[84]
port 306 nsew signal input
rlabel metal2 s 287150 163200 287206 164400 6 la_input[85]
port 307 nsew signal input
rlabel metal2 s 290554 163200 290610 164400 6 la_input[86]
port 308 nsew signal input
rlabel metal2 s 293866 163200 293922 164400 6 la_input[87]
port 309 nsew signal input
rlabel metal2 s 297270 163200 297326 164400 6 la_input[88]
port 310 nsew signal input
rlabel metal2 s 300674 163200 300730 164400 6 la_input[89]
port 311 nsew signal input
rlabel metal2 s 28078 163200 28134 164400 6 la_input[8]
port 312 nsew signal input
rlabel metal2 s 303986 163200 304042 164400 6 la_input[90]
port 313 nsew signal input
rlabel metal2 s 307390 163200 307446 164400 6 la_input[91]
port 314 nsew signal input
rlabel metal2 s 310702 163200 310758 164400 6 la_input[92]
port 315 nsew signal input
rlabel metal2 s 314106 163200 314162 164400 6 la_input[93]
port 316 nsew signal input
rlabel metal2 s 317418 163200 317474 164400 6 la_input[94]
port 317 nsew signal input
rlabel metal2 s 320822 163200 320878 164400 6 la_input[95]
port 318 nsew signal input
rlabel metal2 s 324226 163200 324282 164400 6 la_input[96]
port 319 nsew signal input
rlabel metal2 s 327538 163200 327594 164400 6 la_input[97]
port 320 nsew signal input
rlabel metal2 s 330942 163200 330998 164400 6 la_input[98]
port 321 nsew signal input
rlabel metal2 s 334254 163200 334310 164400 6 la_input[99]
port 322 nsew signal input
rlabel metal2 s 31482 163200 31538 164400 6 la_input[9]
port 323 nsew signal input
rlabel metal2 s 2042 163200 2098 164400 6 la_oenb[0]
port 324 nsew signal tristate
rlabel metal2 s 338486 163200 338542 164400 6 la_oenb[100]
port 325 nsew signal tristate
rlabel metal2 s 341890 163200 341946 164400 6 la_oenb[101]
port 326 nsew signal tristate
rlabel metal2 s 345202 163200 345258 164400 6 la_oenb[102]
port 327 nsew signal tristate
rlabel metal2 s 348606 163200 348662 164400 6 la_oenb[103]
port 328 nsew signal tristate
rlabel metal2 s 351918 163200 351974 164400 6 la_oenb[104]
port 329 nsew signal tristate
rlabel metal2 s 355322 163200 355378 164400 6 la_oenb[105]
port 330 nsew signal tristate
rlabel metal2 s 358634 163200 358690 164400 6 la_oenb[106]
port 331 nsew signal tristate
rlabel metal2 s 362038 163200 362094 164400 6 la_oenb[107]
port 332 nsew signal tristate
rlabel metal2 s 365442 163200 365498 164400 6 la_oenb[108]
port 333 nsew signal tristate
rlabel metal2 s 368754 163200 368810 164400 6 la_oenb[109]
port 334 nsew signal tristate
rlabel metal2 s 35714 163200 35770 164400 6 la_oenb[10]
port 335 nsew signal tristate
rlabel metal2 s 372158 163200 372214 164400 6 la_oenb[110]
port 336 nsew signal tristate
rlabel metal2 s 375470 163200 375526 164400 6 la_oenb[111]
port 337 nsew signal tristate
rlabel metal2 s 378874 163200 378930 164400 6 la_oenb[112]
port 338 nsew signal tristate
rlabel metal2 s 382186 163200 382242 164400 6 la_oenb[113]
port 339 nsew signal tristate
rlabel metal2 s 385590 163200 385646 164400 6 la_oenb[114]
port 340 nsew signal tristate
rlabel metal2 s 388994 163200 389050 164400 6 la_oenb[115]
port 341 nsew signal tristate
rlabel metal2 s 392306 163200 392362 164400 6 la_oenb[116]
port 342 nsew signal tristate
rlabel metal2 s 395710 163200 395766 164400 6 la_oenb[117]
port 343 nsew signal tristate
rlabel metal2 s 399022 163200 399078 164400 6 la_oenb[118]
port 344 nsew signal tristate
rlabel metal2 s 402426 163200 402482 164400 6 la_oenb[119]
port 345 nsew signal tristate
rlabel metal2 s 39026 163200 39082 164400 6 la_oenb[11]
port 346 nsew signal tristate
rlabel metal2 s 405738 163200 405794 164400 6 la_oenb[120]
port 347 nsew signal tristate
rlabel metal2 s 409142 163200 409198 164400 6 la_oenb[121]
port 348 nsew signal tristate
rlabel metal2 s 412546 163200 412602 164400 6 la_oenb[122]
port 349 nsew signal tristate
rlabel metal2 s 415858 163200 415914 164400 6 la_oenb[123]
port 350 nsew signal tristate
rlabel metal2 s 419262 163200 419318 164400 6 la_oenb[124]
port 351 nsew signal tristate
rlabel metal2 s 422574 163200 422630 164400 6 la_oenb[125]
port 352 nsew signal tristate
rlabel metal2 s 425978 163200 426034 164400 6 la_oenb[126]
port 353 nsew signal tristate
rlabel metal2 s 429290 163200 429346 164400 6 la_oenb[127]
port 354 nsew signal tristate
rlabel metal2 s 42430 163200 42486 164400 6 la_oenb[12]
port 355 nsew signal tristate
rlabel metal2 s 45742 163200 45798 164400 6 la_oenb[13]
port 356 nsew signal tristate
rlabel metal2 s 49146 163200 49202 164400 6 la_oenb[14]
port 357 nsew signal tristate
rlabel metal2 s 52458 163200 52514 164400 6 la_oenb[15]
port 358 nsew signal tristate
rlabel metal2 s 55862 163200 55918 164400 6 la_oenb[16]
port 359 nsew signal tristate
rlabel metal2 s 59266 163200 59322 164400 6 la_oenb[17]
port 360 nsew signal tristate
rlabel metal2 s 62578 163200 62634 164400 6 la_oenb[18]
port 361 nsew signal tristate
rlabel metal2 s 65982 163200 66038 164400 6 la_oenb[19]
port 362 nsew signal tristate
rlabel metal2 s 5354 163200 5410 164400 6 la_oenb[1]
port 363 nsew signal tristate
rlabel metal2 s 69294 163200 69350 164400 6 la_oenb[20]
port 364 nsew signal tristate
rlabel metal2 s 72698 163200 72754 164400 6 la_oenb[21]
port 365 nsew signal tristate
rlabel metal2 s 76010 163200 76066 164400 6 la_oenb[22]
port 366 nsew signal tristate
rlabel metal2 s 79414 163200 79470 164400 6 la_oenb[23]
port 367 nsew signal tristate
rlabel metal2 s 82818 163200 82874 164400 6 la_oenb[24]
port 368 nsew signal tristate
rlabel metal2 s 86130 163200 86186 164400 6 la_oenb[25]
port 369 nsew signal tristate
rlabel metal2 s 89534 163200 89590 164400 6 la_oenb[26]
port 370 nsew signal tristate
rlabel metal2 s 92846 163200 92902 164400 6 la_oenb[27]
port 371 nsew signal tristate
rlabel metal2 s 96250 163200 96306 164400 6 la_oenb[28]
port 372 nsew signal tristate
rlabel metal2 s 99562 163200 99618 164400 6 la_oenb[29]
port 373 nsew signal tristate
rlabel metal2 s 8758 163200 8814 164400 6 la_oenb[2]
port 374 nsew signal tristate
rlabel metal2 s 102966 163200 103022 164400 6 la_oenb[30]
port 375 nsew signal tristate
rlabel metal2 s 106370 163200 106426 164400 6 la_oenb[31]
port 376 nsew signal tristate
rlabel metal2 s 109682 163200 109738 164400 6 la_oenb[32]
port 377 nsew signal tristate
rlabel metal2 s 113086 163200 113142 164400 6 la_oenb[33]
port 378 nsew signal tristate
rlabel metal2 s 116398 163200 116454 164400 6 la_oenb[34]
port 379 nsew signal tristate
rlabel metal2 s 119802 163200 119858 164400 6 la_oenb[35]
port 380 nsew signal tristate
rlabel metal2 s 123114 163200 123170 164400 6 la_oenb[36]
port 381 nsew signal tristate
rlabel metal2 s 126518 163200 126574 164400 6 la_oenb[37]
port 382 nsew signal tristate
rlabel metal2 s 129922 163200 129978 164400 6 la_oenb[38]
port 383 nsew signal tristate
rlabel metal2 s 133234 163200 133290 164400 6 la_oenb[39]
port 384 nsew signal tristate
rlabel metal2 s 12162 163200 12218 164400 6 la_oenb[3]
port 385 nsew signal tristate
rlabel metal2 s 136638 163200 136694 164400 6 la_oenb[40]
port 386 nsew signal tristate
rlabel metal2 s 139950 163200 140006 164400 6 la_oenb[41]
port 387 nsew signal tristate
rlabel metal2 s 143354 163200 143410 164400 6 la_oenb[42]
port 388 nsew signal tristate
rlabel metal2 s 146666 163200 146722 164400 6 la_oenb[43]
port 389 nsew signal tristate
rlabel metal2 s 150070 163200 150126 164400 6 la_oenb[44]
port 390 nsew signal tristate
rlabel metal2 s 153474 163200 153530 164400 6 la_oenb[45]
port 391 nsew signal tristate
rlabel metal2 s 156786 163200 156842 164400 6 la_oenb[46]
port 392 nsew signal tristate
rlabel metal2 s 160190 163200 160246 164400 6 la_oenb[47]
port 393 nsew signal tristate
rlabel metal2 s 163502 163200 163558 164400 6 la_oenb[48]
port 394 nsew signal tristate
rlabel metal2 s 166906 163200 166962 164400 6 la_oenb[49]
port 395 nsew signal tristate
rlabel metal2 s 15474 163200 15530 164400 6 la_oenb[4]
port 396 nsew signal tristate
rlabel metal2 s 170218 163200 170274 164400 6 la_oenb[50]
port 397 nsew signal tristate
rlabel metal2 s 173622 163200 173678 164400 6 la_oenb[51]
port 398 nsew signal tristate
rlabel metal2 s 177026 163200 177082 164400 6 la_oenb[52]
port 399 nsew signal tristate
rlabel metal2 s 180338 163200 180394 164400 6 la_oenb[53]
port 400 nsew signal tristate
rlabel metal2 s 183742 163200 183798 164400 6 la_oenb[54]
port 401 nsew signal tristate
rlabel metal2 s 187054 163200 187110 164400 6 la_oenb[55]
port 402 nsew signal tristate
rlabel metal2 s 190458 163200 190514 164400 6 la_oenb[56]
port 403 nsew signal tristate
rlabel metal2 s 193770 163200 193826 164400 6 la_oenb[57]
port 404 nsew signal tristate
rlabel metal2 s 197174 163200 197230 164400 6 la_oenb[58]
port 405 nsew signal tristate
rlabel metal2 s 200578 163200 200634 164400 6 la_oenb[59]
port 406 nsew signal tristate
rlabel metal2 s 18878 163200 18934 164400 6 la_oenb[5]
port 407 nsew signal tristate
rlabel metal2 s 203890 163200 203946 164400 6 la_oenb[60]
port 408 nsew signal tristate
rlabel metal2 s 207294 163200 207350 164400 6 la_oenb[61]
port 409 nsew signal tristate
rlabel metal2 s 210606 163200 210662 164400 6 la_oenb[62]
port 410 nsew signal tristate
rlabel metal2 s 214010 163200 214066 164400 6 la_oenb[63]
port 411 nsew signal tristate
rlabel metal2 s 217322 163200 217378 164400 6 la_oenb[64]
port 412 nsew signal tristate
rlabel metal2 s 220726 163200 220782 164400 6 la_oenb[65]
port 413 nsew signal tristate
rlabel metal2 s 224130 163200 224186 164400 6 la_oenb[66]
port 414 nsew signal tristate
rlabel metal2 s 227442 163200 227498 164400 6 la_oenb[67]
port 415 nsew signal tristate
rlabel metal2 s 230846 163200 230902 164400 6 la_oenb[68]
port 416 nsew signal tristate
rlabel metal2 s 234158 163200 234214 164400 6 la_oenb[69]
port 417 nsew signal tristate
rlabel metal2 s 22190 163200 22246 164400 6 la_oenb[6]
port 418 nsew signal tristate
rlabel metal2 s 237562 163200 237618 164400 6 la_oenb[70]
port 419 nsew signal tristate
rlabel metal2 s 240874 163200 240930 164400 6 la_oenb[71]
port 420 nsew signal tristate
rlabel metal2 s 244278 163200 244334 164400 6 la_oenb[72]
port 421 nsew signal tristate
rlabel metal2 s 247682 163200 247738 164400 6 la_oenb[73]
port 422 nsew signal tristate
rlabel metal2 s 250994 163200 251050 164400 6 la_oenb[74]
port 423 nsew signal tristate
rlabel metal2 s 254398 163200 254454 164400 6 la_oenb[75]
port 424 nsew signal tristate
rlabel metal2 s 257710 163200 257766 164400 6 la_oenb[76]
port 425 nsew signal tristate
rlabel metal2 s 261114 163200 261170 164400 6 la_oenb[77]
port 426 nsew signal tristate
rlabel metal2 s 264426 163200 264482 164400 6 la_oenb[78]
port 427 nsew signal tristate
rlabel metal2 s 267830 163200 267886 164400 6 la_oenb[79]
port 428 nsew signal tristate
rlabel metal2 s 25594 163200 25650 164400 6 la_oenb[7]
port 429 nsew signal tristate
rlabel metal2 s 271234 163200 271290 164400 6 la_oenb[80]
port 430 nsew signal tristate
rlabel metal2 s 274546 163200 274602 164400 6 la_oenb[81]
port 431 nsew signal tristate
rlabel metal2 s 277950 163200 278006 164400 6 la_oenb[82]
port 432 nsew signal tristate
rlabel metal2 s 281262 163200 281318 164400 6 la_oenb[83]
port 433 nsew signal tristate
rlabel metal2 s 284666 163200 284722 164400 6 la_oenb[84]
port 434 nsew signal tristate
rlabel metal2 s 287978 163200 288034 164400 6 la_oenb[85]
port 435 nsew signal tristate
rlabel metal2 s 291382 163200 291438 164400 6 la_oenb[86]
port 436 nsew signal tristate
rlabel metal2 s 294786 163200 294842 164400 6 la_oenb[87]
port 437 nsew signal tristate
rlabel metal2 s 298098 163200 298154 164400 6 la_oenb[88]
port 438 nsew signal tristate
rlabel metal2 s 301502 163200 301558 164400 6 la_oenb[89]
port 439 nsew signal tristate
rlabel metal2 s 28906 163200 28962 164400 6 la_oenb[8]
port 440 nsew signal tristate
rlabel metal2 s 304814 163200 304870 164400 6 la_oenb[90]
port 441 nsew signal tristate
rlabel metal2 s 308218 163200 308274 164400 6 la_oenb[91]
port 442 nsew signal tristate
rlabel metal2 s 311530 163200 311586 164400 6 la_oenb[92]
port 443 nsew signal tristate
rlabel metal2 s 314934 163200 314990 164400 6 la_oenb[93]
port 444 nsew signal tristate
rlabel metal2 s 318338 163200 318394 164400 6 la_oenb[94]
port 445 nsew signal tristate
rlabel metal2 s 321650 163200 321706 164400 6 la_oenb[95]
port 446 nsew signal tristate
rlabel metal2 s 325054 163200 325110 164400 6 la_oenb[96]
port 447 nsew signal tristate
rlabel metal2 s 328366 163200 328422 164400 6 la_oenb[97]
port 448 nsew signal tristate
rlabel metal2 s 331770 163200 331826 164400 6 la_oenb[98]
port 449 nsew signal tristate
rlabel metal2 s 335082 163200 335138 164400 6 la_oenb[99]
port 450 nsew signal tristate
rlabel metal2 s 32310 163200 32366 164400 6 la_oenb[9]
port 451 nsew signal tristate
rlabel metal2 s 2870 163200 2926 164400 6 la_output[0]
port 452 nsew signal tristate
rlabel metal2 s 339314 163200 339370 164400 6 la_output[100]
port 453 nsew signal tristate
rlabel metal2 s 342718 163200 342774 164400 6 la_output[101]
port 454 nsew signal tristate
rlabel metal2 s 346030 163200 346086 164400 6 la_output[102]
port 455 nsew signal tristate
rlabel metal2 s 349434 163200 349490 164400 6 la_output[103]
port 456 nsew signal tristate
rlabel metal2 s 352746 163200 352802 164400 6 la_output[104]
port 457 nsew signal tristate
rlabel metal2 s 356150 163200 356206 164400 6 la_output[105]
port 458 nsew signal tristate
rlabel metal2 s 359554 163200 359610 164400 6 la_output[106]
port 459 nsew signal tristate
rlabel metal2 s 362866 163200 362922 164400 6 la_output[107]
port 460 nsew signal tristate
rlabel metal2 s 366270 163200 366326 164400 6 la_output[108]
port 461 nsew signal tristate
rlabel metal2 s 369582 163200 369638 164400 6 la_output[109]
port 462 nsew signal tristate
rlabel metal2 s 36542 163200 36598 164400 6 la_output[10]
port 463 nsew signal tristate
rlabel metal2 s 372986 163200 373042 164400 6 la_output[110]
port 464 nsew signal tristate
rlabel metal2 s 376298 163200 376354 164400 6 la_output[111]
port 465 nsew signal tristate
rlabel metal2 s 379702 163200 379758 164400 6 la_output[112]
port 466 nsew signal tristate
rlabel metal2 s 383106 163200 383162 164400 6 la_output[113]
port 467 nsew signal tristate
rlabel metal2 s 386418 163200 386474 164400 6 la_output[114]
port 468 nsew signal tristate
rlabel metal2 s 389822 163200 389878 164400 6 la_output[115]
port 469 nsew signal tristate
rlabel metal2 s 393134 163200 393190 164400 6 la_output[116]
port 470 nsew signal tristate
rlabel metal2 s 396538 163200 396594 164400 6 la_output[117]
port 471 nsew signal tristate
rlabel metal2 s 399850 163200 399906 164400 6 la_output[118]
port 472 nsew signal tristate
rlabel metal2 s 403254 163200 403310 164400 6 la_output[119]
port 473 nsew signal tristate
rlabel metal2 s 39854 163200 39910 164400 6 la_output[11]
port 474 nsew signal tristate
rlabel metal2 s 406658 163200 406714 164400 6 la_output[120]
port 475 nsew signal tristate
rlabel metal2 s 409970 163200 410026 164400 6 la_output[121]
port 476 nsew signal tristate
rlabel metal2 s 413374 163200 413430 164400 6 la_output[122]
port 477 nsew signal tristate
rlabel metal2 s 416686 163200 416742 164400 6 la_output[123]
port 478 nsew signal tristate
rlabel metal2 s 420090 163200 420146 164400 6 la_output[124]
port 479 nsew signal tristate
rlabel metal2 s 423402 163200 423458 164400 6 la_output[125]
port 480 nsew signal tristate
rlabel metal2 s 426806 163200 426862 164400 6 la_output[126]
port 481 nsew signal tristate
rlabel metal2 s 430210 163200 430266 164400 6 la_output[127]
port 482 nsew signal tristate
rlabel metal2 s 43258 163200 43314 164400 6 la_output[12]
port 483 nsew signal tristate
rlabel metal2 s 46570 163200 46626 164400 6 la_output[13]
port 484 nsew signal tristate
rlabel metal2 s 49974 163200 50030 164400 6 la_output[14]
port 485 nsew signal tristate
rlabel metal2 s 53378 163200 53434 164400 6 la_output[15]
port 486 nsew signal tristate
rlabel metal2 s 56690 163200 56746 164400 6 la_output[16]
port 487 nsew signal tristate
rlabel metal2 s 60094 163200 60150 164400 6 la_output[17]
port 488 nsew signal tristate
rlabel metal2 s 63406 163200 63462 164400 6 la_output[18]
port 489 nsew signal tristate
rlabel metal2 s 66810 163200 66866 164400 6 la_output[19]
port 490 nsew signal tristate
rlabel metal2 s 6274 163200 6330 164400 6 la_output[1]
port 491 nsew signal tristate
rlabel metal2 s 70122 163200 70178 164400 6 la_output[20]
port 492 nsew signal tristate
rlabel metal2 s 73526 163200 73582 164400 6 la_output[21]
port 493 nsew signal tristate
rlabel metal2 s 76930 163200 76986 164400 6 la_output[22]
port 494 nsew signal tristate
rlabel metal2 s 80242 163200 80298 164400 6 la_output[23]
port 495 nsew signal tristate
rlabel metal2 s 83646 163200 83702 164400 6 la_output[24]
port 496 nsew signal tristate
rlabel metal2 s 86958 163200 87014 164400 6 la_output[25]
port 497 nsew signal tristate
rlabel metal2 s 90362 163200 90418 164400 6 la_output[26]
port 498 nsew signal tristate
rlabel metal2 s 93674 163200 93730 164400 6 la_output[27]
port 499 nsew signal tristate
rlabel metal2 s 97078 163200 97134 164400 6 la_output[28]
port 500 nsew signal tristate
rlabel metal2 s 100482 163200 100538 164400 6 la_output[29]
port 501 nsew signal tristate
rlabel metal2 s 9586 163200 9642 164400 6 la_output[2]
port 502 nsew signal tristate
rlabel metal2 s 103794 163200 103850 164400 6 la_output[30]
port 503 nsew signal tristate
rlabel metal2 s 107198 163200 107254 164400 6 la_output[31]
port 504 nsew signal tristate
rlabel metal2 s 110510 163200 110566 164400 6 la_output[32]
port 505 nsew signal tristate
rlabel metal2 s 113914 163200 113970 164400 6 la_output[33]
port 506 nsew signal tristate
rlabel metal2 s 117226 163200 117282 164400 6 la_output[34]
port 507 nsew signal tristate
rlabel metal2 s 120630 163200 120686 164400 6 la_output[35]
port 508 nsew signal tristate
rlabel metal2 s 124034 163200 124090 164400 6 la_output[36]
port 509 nsew signal tristate
rlabel metal2 s 127346 163200 127402 164400 6 la_output[37]
port 510 nsew signal tristate
rlabel metal2 s 130750 163200 130806 164400 6 la_output[38]
port 511 nsew signal tristate
rlabel metal2 s 134062 163200 134118 164400 6 la_output[39]
port 512 nsew signal tristate
rlabel metal2 s 12990 163200 13046 164400 6 la_output[3]
port 513 nsew signal tristate
rlabel metal2 s 137466 163200 137522 164400 6 la_output[40]
port 514 nsew signal tristate
rlabel metal2 s 140778 163200 140834 164400 6 la_output[41]
port 515 nsew signal tristate
rlabel metal2 s 144182 163200 144238 164400 6 la_output[42]
port 516 nsew signal tristate
rlabel metal2 s 147586 163200 147642 164400 6 la_output[43]
port 517 nsew signal tristate
rlabel metal2 s 150898 163200 150954 164400 6 la_output[44]
port 518 nsew signal tristate
rlabel metal2 s 154302 163200 154358 164400 6 la_output[45]
port 519 nsew signal tristate
rlabel metal2 s 157614 163200 157670 164400 6 la_output[46]
port 520 nsew signal tristate
rlabel metal2 s 161018 163200 161074 164400 6 la_output[47]
port 521 nsew signal tristate
rlabel metal2 s 164330 163200 164386 164400 6 la_output[48]
port 522 nsew signal tristate
rlabel metal2 s 167734 163200 167790 164400 6 la_output[49]
port 523 nsew signal tristate
rlabel metal2 s 16302 163200 16358 164400 6 la_output[4]
port 524 nsew signal tristate
rlabel metal2 s 171138 163200 171194 164400 6 la_output[50]
port 525 nsew signal tristate
rlabel metal2 s 174450 163200 174506 164400 6 la_output[51]
port 526 nsew signal tristate
rlabel metal2 s 177854 163200 177910 164400 6 la_output[52]
port 527 nsew signal tristate
rlabel metal2 s 181166 163200 181222 164400 6 la_output[53]
port 528 nsew signal tristate
rlabel metal2 s 184570 163200 184626 164400 6 la_output[54]
port 529 nsew signal tristate
rlabel metal2 s 187882 163200 187938 164400 6 la_output[55]
port 530 nsew signal tristate
rlabel metal2 s 191286 163200 191342 164400 6 la_output[56]
port 531 nsew signal tristate
rlabel metal2 s 194690 163200 194746 164400 6 la_output[57]
port 532 nsew signal tristate
rlabel metal2 s 198002 163200 198058 164400 6 la_output[58]
port 533 nsew signal tristate
rlabel metal2 s 201406 163200 201462 164400 6 la_output[59]
port 534 nsew signal tristate
rlabel metal2 s 19706 163200 19762 164400 6 la_output[5]
port 535 nsew signal tristate
rlabel metal2 s 204718 163200 204774 164400 6 la_output[60]
port 536 nsew signal tristate
rlabel metal2 s 208122 163200 208178 164400 6 la_output[61]
port 537 nsew signal tristate
rlabel metal2 s 211434 163200 211490 164400 6 la_output[62]
port 538 nsew signal tristate
rlabel metal2 s 214838 163200 214894 164400 6 la_output[63]
port 539 nsew signal tristate
rlabel metal2 s 218242 163200 218298 164400 6 la_output[64]
port 540 nsew signal tristate
rlabel metal2 s 221554 163200 221610 164400 6 la_output[65]
port 541 nsew signal tristate
rlabel metal2 s 224958 163200 225014 164400 6 la_output[66]
port 542 nsew signal tristate
rlabel metal2 s 228270 163200 228326 164400 6 la_output[67]
port 543 nsew signal tristate
rlabel metal2 s 231674 163200 231730 164400 6 la_output[68]
port 544 nsew signal tristate
rlabel metal2 s 234986 163200 235042 164400 6 la_output[69]
port 545 nsew signal tristate
rlabel metal2 s 23018 163200 23074 164400 6 la_output[6]
port 546 nsew signal tristate
rlabel metal2 s 238390 163200 238446 164400 6 la_output[70]
port 547 nsew signal tristate
rlabel metal2 s 241794 163200 241850 164400 6 la_output[71]
port 548 nsew signal tristate
rlabel metal2 s 245106 163200 245162 164400 6 la_output[72]
port 549 nsew signal tristate
rlabel metal2 s 248510 163200 248566 164400 6 la_output[73]
port 550 nsew signal tristate
rlabel metal2 s 251822 163200 251878 164400 6 la_output[74]
port 551 nsew signal tristate
rlabel metal2 s 255226 163200 255282 164400 6 la_output[75]
port 552 nsew signal tristate
rlabel metal2 s 258538 163200 258594 164400 6 la_output[76]
port 553 nsew signal tristate
rlabel metal2 s 261942 163200 261998 164400 6 la_output[77]
port 554 nsew signal tristate
rlabel metal2 s 265346 163200 265402 164400 6 la_output[78]
port 555 nsew signal tristate
rlabel metal2 s 268658 163200 268714 164400 6 la_output[79]
port 556 nsew signal tristate
rlabel metal2 s 26422 163200 26478 164400 6 la_output[7]
port 557 nsew signal tristate
rlabel metal2 s 272062 163200 272118 164400 6 la_output[80]
port 558 nsew signal tristate
rlabel metal2 s 275374 163200 275430 164400 6 la_output[81]
port 559 nsew signal tristate
rlabel metal2 s 278778 163200 278834 164400 6 la_output[82]
port 560 nsew signal tristate
rlabel metal2 s 282090 163200 282146 164400 6 la_output[83]
port 561 nsew signal tristate
rlabel metal2 s 285494 163200 285550 164400 6 la_output[84]
port 562 nsew signal tristate
rlabel metal2 s 288898 163200 288954 164400 6 la_output[85]
port 563 nsew signal tristate
rlabel metal2 s 292210 163200 292266 164400 6 la_output[86]
port 564 nsew signal tristate
rlabel metal2 s 295614 163200 295670 164400 6 la_output[87]
port 565 nsew signal tristate
rlabel metal2 s 298926 163200 298982 164400 6 la_output[88]
port 566 nsew signal tristate
rlabel metal2 s 302330 163200 302386 164400 6 la_output[89]
port 567 nsew signal tristate
rlabel metal2 s 29826 163200 29882 164400 6 la_output[8]
port 568 nsew signal tristate
rlabel metal2 s 305642 163200 305698 164400 6 la_output[90]
port 569 nsew signal tristate
rlabel metal2 s 309046 163200 309102 164400 6 la_output[91]
port 570 nsew signal tristate
rlabel metal2 s 312450 163200 312506 164400 6 la_output[92]
port 571 nsew signal tristate
rlabel metal2 s 315762 163200 315818 164400 6 la_output[93]
port 572 nsew signal tristate
rlabel metal2 s 319166 163200 319222 164400 6 la_output[94]
port 573 nsew signal tristate
rlabel metal2 s 322478 163200 322534 164400 6 la_output[95]
port 574 nsew signal tristate
rlabel metal2 s 325882 163200 325938 164400 6 la_output[96]
port 575 nsew signal tristate
rlabel metal2 s 329194 163200 329250 164400 6 la_output[97]
port 576 nsew signal tristate
rlabel metal2 s 332598 163200 332654 164400 6 la_output[98]
port 577 nsew signal tristate
rlabel metal2 s 336002 163200 336058 164400 6 la_output[99]
port 578 nsew signal tristate
rlabel metal2 s 33138 163200 33194 164400 6 la_output[9]
port 579 nsew signal tristate
rlabel metal2 s 431038 163200 431094 164400 6 mprj_ack_i
port 580 nsew signal input
rlabel metal2 s 435178 163200 435234 164400 6 mprj_adr_o[0]
port 581 nsew signal tristate
rlabel metal2 s 463790 163200 463846 164400 6 mprj_adr_o[10]
port 582 nsew signal tristate
rlabel metal2 s 466366 163200 466422 164400 6 mprj_adr_o[11]
port 583 nsew signal tristate
rlabel metal2 s 468850 163200 468906 164400 6 mprj_adr_o[12]
port 584 nsew signal tristate
rlabel metal2 s 471426 163200 471482 164400 6 mprj_adr_o[13]
port 585 nsew signal tristate
rlabel metal2 s 473910 163200 473966 164400 6 mprj_adr_o[14]
port 586 nsew signal tristate
rlabel metal2 s 476394 163200 476450 164400 6 mprj_adr_o[15]
port 587 nsew signal tristate
rlabel metal2 s 478970 163200 479026 164400 6 mprj_adr_o[16]
port 588 nsew signal tristate
rlabel metal2 s 481454 163200 481510 164400 6 mprj_adr_o[17]
port 589 nsew signal tristate
rlabel metal2 s 484030 163200 484086 164400 6 mprj_adr_o[18]
port 590 nsew signal tristate
rlabel metal2 s 486514 163200 486570 164400 6 mprj_adr_o[19]
port 591 nsew signal tristate
rlabel metal2 s 438582 163200 438638 164400 6 mprj_adr_o[1]
port 592 nsew signal tristate
rlabel metal2 s 489090 163200 489146 164400 6 mprj_adr_o[20]
port 593 nsew signal tristate
rlabel metal2 s 491574 163200 491630 164400 6 mprj_adr_o[21]
port 594 nsew signal tristate
rlabel metal2 s 494058 163200 494114 164400 6 mprj_adr_o[22]
port 595 nsew signal tristate
rlabel metal2 s 496634 163200 496690 164400 6 mprj_adr_o[23]
port 596 nsew signal tristate
rlabel metal2 s 499118 163200 499174 164400 6 mprj_adr_o[24]
port 597 nsew signal tristate
rlabel metal2 s 501694 163200 501750 164400 6 mprj_adr_o[25]
port 598 nsew signal tristate
rlabel metal2 s 504178 163200 504234 164400 6 mprj_adr_o[26]
port 599 nsew signal tristate
rlabel metal2 s 506754 163200 506810 164400 6 mprj_adr_o[27]
port 600 nsew signal tristate
rlabel metal2 s 509238 163200 509294 164400 6 mprj_adr_o[28]
port 601 nsew signal tristate
rlabel metal2 s 511722 163200 511778 164400 6 mprj_adr_o[29]
port 602 nsew signal tristate
rlabel metal2 s 441986 163200 442042 164400 6 mprj_adr_o[2]
port 603 nsew signal tristate
rlabel metal2 s 514298 163200 514354 164400 6 mprj_adr_o[30]
port 604 nsew signal tristate
rlabel metal2 s 516782 163200 516838 164400 6 mprj_adr_o[31]
port 605 nsew signal tristate
rlabel metal2 s 445298 163200 445354 164400 6 mprj_adr_o[3]
port 606 nsew signal tristate
rlabel metal2 s 448702 163200 448758 164400 6 mprj_adr_o[4]
port 607 nsew signal tristate
rlabel metal2 s 451186 163200 451242 164400 6 mprj_adr_o[5]
port 608 nsew signal tristate
rlabel metal2 s 453762 163200 453818 164400 6 mprj_adr_o[6]
port 609 nsew signal tristate
rlabel metal2 s 456246 163200 456302 164400 6 mprj_adr_o[7]
port 610 nsew signal tristate
rlabel metal2 s 458730 163200 458786 164400 6 mprj_adr_o[8]
port 611 nsew signal tristate
rlabel metal2 s 461306 163200 461362 164400 6 mprj_adr_o[9]
port 612 nsew signal tristate
rlabel metal2 s 431866 163200 431922 164400 6 mprj_cyc_o
port 613 nsew signal tristate
rlabel metal2 s 436098 163200 436154 164400 6 mprj_dat_i[0]
port 614 nsew signal input
rlabel metal2 s 464618 163200 464674 164400 6 mprj_dat_i[10]
port 615 nsew signal input
rlabel metal2 s 467194 163200 467250 164400 6 mprj_dat_i[11]
port 616 nsew signal input
rlabel metal2 s 469678 163200 469734 164400 6 mprj_dat_i[12]
port 617 nsew signal input
rlabel metal2 s 472254 163200 472310 164400 6 mprj_dat_i[13]
port 618 nsew signal input
rlabel metal2 s 474738 163200 474794 164400 6 mprj_dat_i[14]
port 619 nsew signal input
rlabel metal2 s 477314 163200 477370 164400 6 mprj_dat_i[15]
port 620 nsew signal input
rlabel metal2 s 479798 163200 479854 164400 6 mprj_dat_i[16]
port 621 nsew signal input
rlabel metal2 s 482282 163200 482338 164400 6 mprj_dat_i[17]
port 622 nsew signal input
rlabel metal2 s 484858 163200 484914 164400 6 mprj_dat_i[18]
port 623 nsew signal input
rlabel metal2 s 487342 163200 487398 164400 6 mprj_dat_i[19]
port 624 nsew signal input
rlabel metal2 s 439410 163200 439466 164400 6 mprj_dat_i[1]
port 625 nsew signal input
rlabel metal2 s 489918 163200 489974 164400 6 mprj_dat_i[20]
port 626 nsew signal input
rlabel metal2 s 492402 163200 492458 164400 6 mprj_dat_i[21]
port 627 nsew signal input
rlabel metal2 s 494978 163200 495034 164400 6 mprj_dat_i[22]
port 628 nsew signal input
rlabel metal2 s 497462 163200 497518 164400 6 mprj_dat_i[23]
port 629 nsew signal input
rlabel metal2 s 499946 163200 500002 164400 6 mprj_dat_i[24]
port 630 nsew signal input
rlabel metal2 s 502522 163200 502578 164400 6 mprj_dat_i[25]
port 631 nsew signal input
rlabel metal2 s 505006 163200 505062 164400 6 mprj_dat_i[26]
port 632 nsew signal input
rlabel metal2 s 507582 163200 507638 164400 6 mprj_dat_i[27]
port 633 nsew signal input
rlabel metal2 s 510066 163200 510122 164400 6 mprj_dat_i[28]
port 634 nsew signal input
rlabel metal2 s 512642 163200 512698 164400 6 mprj_dat_i[29]
port 635 nsew signal input
rlabel metal2 s 442814 163200 442870 164400 6 mprj_dat_i[2]
port 636 nsew signal input
rlabel metal2 s 515126 163200 515182 164400 6 mprj_dat_i[30]
port 637 nsew signal input
rlabel metal2 s 517610 163200 517666 164400 6 mprj_dat_i[31]
port 638 nsew signal input
rlabel metal2 s 446126 163200 446182 164400 6 mprj_dat_i[3]
port 639 nsew signal input
rlabel metal2 s 449530 163200 449586 164400 6 mprj_dat_i[4]
port 640 nsew signal input
rlabel metal2 s 452014 163200 452070 164400 6 mprj_dat_i[5]
port 641 nsew signal input
rlabel metal2 s 454590 163200 454646 164400 6 mprj_dat_i[6]
port 642 nsew signal input
rlabel metal2 s 457074 163200 457130 164400 6 mprj_dat_i[7]
port 643 nsew signal input
rlabel metal2 s 459650 163200 459706 164400 6 mprj_dat_i[8]
port 644 nsew signal input
rlabel metal2 s 462134 163200 462190 164400 6 mprj_dat_i[9]
port 645 nsew signal input
rlabel metal2 s 436926 163200 436982 164400 6 mprj_dat_o[0]
port 646 nsew signal tristate
rlabel metal2 s 465538 163200 465594 164400 6 mprj_dat_o[10]
port 647 nsew signal tristate
rlabel metal2 s 468022 163200 468078 164400 6 mprj_dat_o[11]
port 648 nsew signal tristate
rlabel metal2 s 470506 163200 470562 164400 6 mprj_dat_o[12]
port 649 nsew signal tristate
rlabel metal2 s 473082 163200 473138 164400 6 mprj_dat_o[13]
port 650 nsew signal tristate
rlabel metal2 s 475566 163200 475622 164400 6 mprj_dat_o[14]
port 651 nsew signal tristate
rlabel metal2 s 478142 163200 478198 164400 6 mprj_dat_o[15]
port 652 nsew signal tristate
rlabel metal2 s 480626 163200 480682 164400 6 mprj_dat_o[16]
port 653 nsew signal tristate
rlabel metal2 s 483202 163200 483258 164400 6 mprj_dat_o[17]
port 654 nsew signal tristate
rlabel metal2 s 485686 163200 485742 164400 6 mprj_dat_o[18]
port 655 nsew signal tristate
rlabel metal2 s 488170 163200 488226 164400 6 mprj_dat_o[19]
port 656 nsew signal tristate
rlabel metal2 s 440238 163200 440294 164400 6 mprj_dat_o[1]
port 657 nsew signal tristate
rlabel metal2 s 490746 163200 490802 164400 6 mprj_dat_o[20]
port 658 nsew signal tristate
rlabel metal2 s 493230 163200 493286 164400 6 mprj_dat_o[21]
port 659 nsew signal tristate
rlabel metal2 s 495806 163200 495862 164400 6 mprj_dat_o[22]
port 660 nsew signal tristate
rlabel metal2 s 498290 163200 498346 164400 6 mprj_dat_o[23]
port 661 nsew signal tristate
rlabel metal2 s 500866 163200 500922 164400 6 mprj_dat_o[24]
port 662 nsew signal tristate
rlabel metal2 s 503350 163200 503406 164400 6 mprj_dat_o[25]
port 663 nsew signal tristate
rlabel metal2 s 505834 163200 505890 164400 6 mprj_dat_o[26]
port 664 nsew signal tristate
rlabel metal2 s 508410 163200 508466 164400 6 mprj_dat_o[27]
port 665 nsew signal tristate
rlabel metal2 s 510894 163200 510950 164400 6 mprj_dat_o[28]
port 666 nsew signal tristate
rlabel metal2 s 513470 163200 513526 164400 6 mprj_dat_o[29]
port 667 nsew signal tristate
rlabel metal2 s 443642 163200 443698 164400 6 mprj_dat_o[2]
port 668 nsew signal tristate
rlabel metal2 s 515954 163200 516010 164400 6 mprj_dat_o[30]
port 669 nsew signal tristate
rlabel metal2 s 518530 163200 518586 164400 6 mprj_dat_o[31]
port 670 nsew signal tristate
rlabel metal2 s 446954 163200 447010 164400 6 mprj_dat_o[3]
port 671 nsew signal tristate
rlabel metal2 s 450358 163200 450414 164400 6 mprj_dat_o[4]
port 672 nsew signal tristate
rlabel metal2 s 452842 163200 452898 164400 6 mprj_dat_o[5]
port 673 nsew signal tristate
rlabel metal2 s 455418 163200 455474 164400 6 mprj_dat_o[6]
port 674 nsew signal tristate
rlabel metal2 s 457902 163200 457958 164400 6 mprj_dat_o[7]
port 675 nsew signal tristate
rlabel metal2 s 460478 163200 460534 164400 6 mprj_dat_o[8]
port 676 nsew signal tristate
rlabel metal2 s 462962 163200 463018 164400 6 mprj_dat_o[9]
port 677 nsew signal tristate
rlabel metal2 s 437754 163200 437810 164400 6 mprj_sel_o[0]
port 678 nsew signal tristate
rlabel metal2 s 441066 163200 441122 164400 6 mprj_sel_o[1]
port 679 nsew signal tristate
rlabel metal2 s 444470 163200 444526 164400 6 mprj_sel_o[2]
port 680 nsew signal tristate
rlabel metal2 s 447874 163200 447930 164400 6 mprj_sel_o[3]
port 681 nsew signal tristate
rlabel metal2 s 432694 163200 432750 164400 6 mprj_stb_o
port 682 nsew signal tristate
rlabel metal2 s 433522 163200 433578 164400 6 mprj_wb_iena
port 683 nsew signal tristate
rlabel metal2 s 434350 163200 434406 164400 6 mprj_we_o
port 684 nsew signal tristate
rlabel metal3 s 523200 90176 524400 90296 6 qspi_enabled
port 685 nsew signal tristate
rlabel metal3 s 523200 84192 524400 84312 6 ser_rx
port 686 nsew signal input
rlabel metal3 s 523200 85688 524400 85808 6 ser_tx
port 687 nsew signal tristate
rlabel metal3 s 523200 81064 524400 81184 6 spi_csb
port 688 nsew signal tristate
rlabel metal3 s 523200 87184 524400 87304 6 spi_enabled
port 689 nsew signal tristate
rlabel metal3 s 523200 79568 524400 79688 6 spi_sck
port 690 nsew signal tristate
rlabel metal3 s 523200 82696 524400 82816 6 spi_sdi
port 691 nsew signal input
rlabel metal3 s 523200 78072 524400 78192 6 spi_sdo
port 692 nsew signal tristate
rlabel metal3 s 523200 76576 524400 76696 6 spi_sdoenb
port 693 nsew signal tristate
rlabel metal3 s 523200 2184 524400 2304 6 sram_ro_addr[0]
port 694 nsew signal input
rlabel metal3 s 523200 3680 524400 3800 6 sram_ro_addr[1]
port 695 nsew signal input
rlabel metal3 s 523200 5176 524400 5296 6 sram_ro_addr[2]
port 696 nsew signal input
rlabel metal3 s 523200 6672 524400 6792 6 sram_ro_addr[3]
port 697 nsew signal input
rlabel metal3 s 523200 8168 524400 8288 6 sram_ro_addr[4]
port 698 nsew signal input
rlabel metal3 s 523200 9800 524400 9920 6 sram_ro_addr[5]
port 699 nsew signal input
rlabel metal3 s 523200 11296 524400 11416 6 sram_ro_addr[6]
port 700 nsew signal input
rlabel metal3 s 523200 12792 524400 12912 6 sram_ro_addr[7]
port 701 nsew signal input
rlabel metal3 s 523200 14288 524400 14408 6 sram_ro_clk
port 702 nsew signal input
rlabel metal3 s 523200 688 524400 808 6 sram_ro_csb
port 703 nsew signal input
rlabel metal3 s 523200 15784 524400 15904 6 sram_ro_data[0]
port 704 nsew signal tristate
rlabel metal3 s 523200 31016 524400 31136 6 sram_ro_data[10]
port 705 nsew signal tristate
rlabel metal3 s 523200 32512 524400 32632 6 sram_ro_data[11]
port 706 nsew signal tristate
rlabel metal3 s 523200 34008 524400 34128 6 sram_ro_data[12]
port 707 nsew signal tristate
rlabel metal3 s 523200 35504 524400 35624 6 sram_ro_data[13]
port 708 nsew signal tristate
rlabel metal3 s 523200 37136 524400 37256 6 sram_ro_data[14]
port 709 nsew signal tristate
rlabel metal3 s 523200 38632 524400 38752 6 sram_ro_data[15]
port 710 nsew signal tristate
rlabel metal3 s 523200 40128 524400 40248 6 sram_ro_data[16]
port 711 nsew signal tristate
rlabel metal3 s 523200 41624 524400 41744 6 sram_ro_data[17]
port 712 nsew signal tristate
rlabel metal3 s 523200 43120 524400 43240 6 sram_ro_data[18]
port 713 nsew signal tristate
rlabel metal3 s 523200 44616 524400 44736 6 sram_ro_data[19]
port 714 nsew signal tristate
rlabel metal3 s 523200 17280 524400 17400 6 sram_ro_data[1]
port 715 nsew signal tristate
rlabel metal3 s 523200 46248 524400 46368 6 sram_ro_data[20]
port 716 nsew signal tristate
rlabel metal3 s 523200 47744 524400 47864 6 sram_ro_data[21]
port 717 nsew signal tristate
rlabel metal3 s 523200 49240 524400 49360 6 sram_ro_data[22]
port 718 nsew signal tristate
rlabel metal3 s 523200 50736 524400 50856 6 sram_ro_data[23]
port 719 nsew signal tristate
rlabel metal3 s 523200 52232 524400 52352 6 sram_ro_data[24]
port 720 nsew signal tristate
rlabel metal3 s 523200 53728 524400 53848 6 sram_ro_data[25]
port 721 nsew signal tristate
rlabel metal3 s 523200 55360 524400 55480 6 sram_ro_data[26]
port 722 nsew signal tristate
rlabel metal3 s 523200 56856 524400 56976 6 sram_ro_data[27]
port 723 nsew signal tristate
rlabel metal3 s 523200 58352 524400 58472 6 sram_ro_data[28]
port 724 nsew signal tristate
rlabel metal3 s 523200 59848 524400 59968 6 sram_ro_data[29]
port 725 nsew signal tristate
rlabel metal3 s 523200 18912 524400 19032 6 sram_ro_data[2]
port 726 nsew signal tristate
rlabel metal3 s 523200 61344 524400 61464 6 sram_ro_data[30]
port 727 nsew signal tristate
rlabel metal3 s 523200 62840 524400 62960 6 sram_ro_data[31]
port 728 nsew signal tristate
rlabel metal3 s 523200 20408 524400 20528 6 sram_ro_data[3]
port 729 nsew signal tristate
rlabel metal3 s 523200 21904 524400 22024 6 sram_ro_data[4]
port 730 nsew signal tristate
rlabel metal3 s 523200 23400 524400 23520 6 sram_ro_data[5]
port 731 nsew signal tristate
rlabel metal3 s 523200 24896 524400 25016 6 sram_ro_data[6]
port 732 nsew signal tristate
rlabel metal3 s 523200 26392 524400 26512 6 sram_ro_data[7]
port 733 nsew signal tristate
rlabel metal3 s 523200 28024 524400 28144 6 sram_ro_data[8]
port 734 nsew signal tristate
rlabel metal3 s 523200 29520 524400 29640 6 sram_ro_data[9]
port 735 nsew signal tristate
rlabel metal3 s 523200 70456 524400 70576 6 trap
port 736 nsew signal tristate
rlabel metal3 s 523200 88680 524400 88800 6 uart_enabled
port 737 nsew signal tristate
rlabel metal2 s 519358 163200 519414 164400 6 user_irq_ena[0]
port 738 nsew signal tristate
rlabel metal2 s 520186 163200 520242 164400 6 user_irq_ena[1]
port 739 nsew signal tristate
rlabel metal2 s 521014 163200 521070 164400 6 user_irq_ena[2]
port 740 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 524000 164000
<< end >>
