VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DFFRAM
  CLASS BLOCK ;
  FOREIGN DFFRAM ;
  ORIGIN 0.000 0.000 ;
  SIZE 850.000 BY 550.000 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 546.000 33.030 550.000 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 546.000 98.350 550.000 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 546.000 163.670 550.000 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 546.000 228.990 550.000 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 546.000 294.310 550.000 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.350 546.000 359.630 550.000 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.670 546.000 424.950 550.000 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.450 546.000 490.730 550.000 ;
    END
  END A[7]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 0.000 425.410 4.000 ;
    END
  END CLK
  PIN Di[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 846.000 8.200 850.000 8.800 ;
    END
  END Di[0]
  PIN Di[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 846.000 179.560 850.000 180.160 ;
    END
  END Di[10]
  PIN Di[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 846.000 197.240 850.000 197.840 ;
    END
  END Di[11]
  PIN Di[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 846.000 214.240 850.000 214.840 ;
    END
  END Di[12]
  PIN Di[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 846.000 231.240 850.000 231.840 ;
    END
  END Di[13]
  PIN Di[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 846.000 248.240 850.000 248.840 ;
    END
  END Di[14]
  PIN Di[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 846.000 265.920 850.000 266.520 ;
    END
  END Di[15]
  PIN Di[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 846.000 282.920 850.000 283.520 ;
    END
  END Di[16]
  PIN Di[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 846.000 299.920 850.000 300.520 ;
    END
  END Di[17]
  PIN Di[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 846.000 317.600 850.000 318.200 ;
    END
  END Di[18]
  PIN Di[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 846.000 334.600 850.000 335.200 ;
    END
  END Di[19]
  PIN Di[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 846.000 25.200 850.000 25.800 ;
    END
  END Di[1]
  PIN Di[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 846.000 351.600 850.000 352.200 ;
    END
  END Di[20]
  PIN Di[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 846.000 368.600 850.000 369.200 ;
    END
  END Di[21]
  PIN Di[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 846.000 386.280 850.000 386.880 ;
    END
  END Di[22]
  PIN Di[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 846.000 403.280 850.000 403.880 ;
    END
  END Di[23]
  PIN Di[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 846.000 420.280 850.000 420.880 ;
    END
  END Di[24]
  PIN Di[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 846.000 437.960 850.000 438.560 ;
    END
  END Di[25]
  PIN Di[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 846.000 454.960 850.000 455.560 ;
    END
  END Di[26]
  PIN Di[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 846.000 471.960 850.000 472.560 ;
    END
  END Di[27]
  PIN Di[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 846.000 488.960 850.000 489.560 ;
    END
  END Di[28]
  PIN Di[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 846.000 506.640 850.000 507.240 ;
    END
  END Di[29]
  PIN Di[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 846.000 42.200 850.000 42.800 ;
    END
  END Di[2]
  PIN Di[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 846.000 523.640 850.000 524.240 ;
    END
  END Di[30]
  PIN Di[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 846.000 540.640 850.000 541.240 ;
    END
  END Di[31]
  PIN Di[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 846.000 59.200 850.000 59.800 ;
    END
  END Di[3]
  PIN Di[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 846.000 76.880 850.000 77.480 ;
    END
  END Di[4]
  PIN Di[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 846.000 93.880 850.000 94.480 ;
    END
  END Di[5]
  PIN Di[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 846.000 110.880 850.000 111.480 ;
    END
  END Di[6]
  PIN Di[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 846.000 127.880 850.000 128.480 ;
    END
  END Di[7]
  PIN Di[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 846.000 145.560 850.000 146.160 ;
    END
  END Di[8]
  PIN Di[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 846.000 162.560 850.000 163.160 ;
    END
  END Di[9]
  PIN Do[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END Do[0]
  PIN Do[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END Do[10]
  PIN Do[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END Do[11]
  PIN Do[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END Do[12]
  PIN Do[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END Do[13]
  PIN Do[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END Do[14]
  PIN Do[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.920 4.000 266.520 ;
    END
  END Do[15]
  PIN Do[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END Do[16]
  PIN Do[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.920 4.000 300.520 ;
    END
  END Do[17]
  PIN Do[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 317.600 4.000 318.200 ;
    END
  END Do[18]
  PIN Do[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.600 4.000 335.200 ;
    END
  END Do[19]
  PIN Do[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END Do[1]
  PIN Do[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 351.600 4.000 352.200 ;
    END
  END Do[20]
  PIN Do[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.600 4.000 369.200 ;
    END
  END Do[21]
  PIN Do[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.280 4.000 386.880 ;
    END
  END Do[22]
  PIN Do[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.280 4.000 403.880 ;
    END
  END Do[23]
  PIN Do[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.280 4.000 420.880 ;
    END
  END Do[24]
  PIN Do[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.960 4.000 438.560 ;
    END
  END Do[25]
  PIN Do[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 454.960 4.000 455.560 ;
    END
  END Do[26]
  PIN Do[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.960 4.000 472.560 ;
    END
  END Do[27]
  PIN Do[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.960 4.000 489.560 ;
    END
  END Do[28]
  PIN Do[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 506.640 4.000 507.240 ;
    END
  END Do[29]
  PIN Do[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END Do[2]
  PIN Do[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END Do[30]
  PIN Do[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 540.640 4.000 541.240 ;
    END
  END Do[31]
  PIN Do[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 4.000 59.800 ;
    END
  END Do[3]
  PIN Do[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 4.000 77.480 ;
    END
  END Do[4]
  PIN Do[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END Do[5]
  PIN Do[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.880 4.000 111.480 ;
    END
  END Do[6]
  PIN Do[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END Do[7]
  PIN Do[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END Do[8]
  PIN Do[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.560 4.000 163.160 ;
    END
  END Do[9]
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.050 546.000 817.330 550.000 ;
    END
  END EN
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 844.100 104.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 256.260 844.100 257.860 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 409.440 844.100 411.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 538.800 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 844.100 28.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 179.670 844.100 181.270 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 332.850 844.100 334.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 486.030 844.100 487.630 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 538.800 ;
    END
  END VPWR
  PIN WE[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.770 546.000 556.050 550.000 ;
    END
  END WE[0]
  PIN WE[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.090 546.000 621.370 550.000 ;
    END
  END WE[1]
  PIN WE[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.410 546.000 686.690 550.000 ;
    END
  END WE[2]
  PIN WE[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 751.730 546.000 752.010 550.000 ;
    END
  END WE[3]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 845.335 538.645 ;
      LAYER met1 ;
        RECT 5.520 10.240 845.395 538.800 ;
      LAYER met2 ;
        RECT 7.000 545.720 32.470 546.450 ;
        RECT 33.310 545.720 97.790 546.450 ;
        RECT 98.630 545.720 163.110 546.450 ;
        RECT 163.950 545.720 228.430 546.450 ;
        RECT 229.270 545.720 293.750 546.450 ;
        RECT 294.590 545.720 359.070 546.450 ;
        RECT 359.910 545.720 424.390 546.450 ;
        RECT 425.230 545.720 490.170 546.450 ;
        RECT 491.010 545.720 555.490 546.450 ;
        RECT 556.330 545.720 620.810 546.450 ;
        RECT 621.650 545.720 686.130 546.450 ;
        RECT 686.970 545.720 751.450 546.450 ;
        RECT 752.290 545.720 816.770 546.450 ;
        RECT 817.610 545.720 844.930 546.450 ;
        RECT 7.000 4.280 844.930 545.720 ;
        RECT 7.000 3.670 424.850 4.280 ;
        RECT 425.690 3.670 844.930 4.280 ;
      LAYER met3 ;
        RECT 4.400 540.240 845.600 541.105 ;
        RECT 4.000 524.640 846.000 540.240 ;
        RECT 4.400 523.240 845.600 524.640 ;
        RECT 4.000 507.640 846.000 523.240 ;
        RECT 4.400 506.240 845.600 507.640 ;
        RECT 4.000 489.960 846.000 506.240 ;
        RECT 4.400 488.560 845.600 489.960 ;
        RECT 4.000 472.960 846.000 488.560 ;
        RECT 4.400 471.560 845.600 472.960 ;
        RECT 4.000 455.960 846.000 471.560 ;
        RECT 4.400 454.560 845.600 455.960 ;
        RECT 4.000 438.960 846.000 454.560 ;
        RECT 4.400 437.560 845.600 438.960 ;
        RECT 4.000 421.280 846.000 437.560 ;
        RECT 4.400 419.880 845.600 421.280 ;
        RECT 4.000 404.280 846.000 419.880 ;
        RECT 4.400 402.880 845.600 404.280 ;
        RECT 4.000 387.280 846.000 402.880 ;
        RECT 4.400 385.880 845.600 387.280 ;
        RECT 4.000 369.600 846.000 385.880 ;
        RECT 4.400 368.200 845.600 369.600 ;
        RECT 4.000 352.600 846.000 368.200 ;
        RECT 4.400 351.200 845.600 352.600 ;
        RECT 4.000 335.600 846.000 351.200 ;
        RECT 4.400 334.200 845.600 335.600 ;
        RECT 4.000 318.600 846.000 334.200 ;
        RECT 4.400 317.200 845.600 318.600 ;
        RECT 4.000 300.920 846.000 317.200 ;
        RECT 4.400 299.520 845.600 300.920 ;
        RECT 4.000 283.920 846.000 299.520 ;
        RECT 4.400 282.520 845.600 283.920 ;
        RECT 4.000 266.920 846.000 282.520 ;
        RECT 4.400 265.520 845.600 266.920 ;
        RECT 4.000 249.240 846.000 265.520 ;
        RECT 4.400 247.840 845.600 249.240 ;
        RECT 4.000 232.240 846.000 247.840 ;
        RECT 4.400 230.840 845.600 232.240 ;
        RECT 4.000 215.240 846.000 230.840 ;
        RECT 4.400 213.840 845.600 215.240 ;
        RECT 4.000 198.240 846.000 213.840 ;
        RECT 4.400 196.840 845.600 198.240 ;
        RECT 4.000 180.560 846.000 196.840 ;
        RECT 4.400 179.160 845.600 180.560 ;
        RECT 4.000 163.560 846.000 179.160 ;
        RECT 4.400 162.160 845.600 163.560 ;
        RECT 4.000 146.560 846.000 162.160 ;
        RECT 4.400 145.160 845.600 146.560 ;
        RECT 4.000 128.880 846.000 145.160 ;
        RECT 4.400 127.480 845.600 128.880 ;
        RECT 4.000 111.880 846.000 127.480 ;
        RECT 4.400 110.480 845.600 111.880 ;
        RECT 4.000 94.880 846.000 110.480 ;
        RECT 4.400 93.480 845.600 94.880 ;
        RECT 4.000 77.880 846.000 93.480 ;
        RECT 4.400 76.480 845.600 77.880 ;
        RECT 4.000 60.200 846.000 76.480 ;
        RECT 4.400 58.800 845.600 60.200 ;
        RECT 4.000 43.200 846.000 58.800 ;
        RECT 4.400 41.800 845.600 43.200 ;
        RECT 4.000 26.200 846.000 41.800 ;
        RECT 4.400 24.800 845.600 26.200 ;
        RECT 4.000 9.200 846.000 24.800 ;
        RECT 4.400 8.335 845.600 9.200 ;
      LAYER met4 ;
        RECT 25.135 26.015 97.440 528.185 ;
        RECT 99.840 26.015 174.240 528.185 ;
        RECT 176.640 26.015 251.040 528.185 ;
        RECT 253.440 26.015 327.840 528.185 ;
        RECT 330.240 26.015 404.640 528.185 ;
        RECT 407.040 26.015 481.440 528.185 ;
        RECT 483.840 26.015 558.240 528.185 ;
        RECT 560.640 26.015 635.040 528.185 ;
        RECT 637.440 26.015 711.840 528.185 ;
        RECT 714.240 26.015 769.745 528.185 ;
  END
END DFFRAM
END LIBRARY

