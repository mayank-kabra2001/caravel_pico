magic
tech sky130A
magscale 1 2
timestamp 1637942417
<< obsli1 >>
rect 2024 2159 397900 145809
<< obsm1 >>
rect 290 1980 399726 147960
<< metal2 >>
rect 294 147200 350 148000
rect 846 147200 902 148000
rect 1490 147200 1546 148000
rect 2134 147200 2190 148000
rect 2778 147200 2834 148000
rect 3422 147200 3478 148000
rect 4066 147200 4122 148000
rect 4710 147200 4766 148000
rect 5354 147200 5410 148000
rect 5998 147200 6054 148000
rect 6642 147200 6698 148000
rect 7286 147200 7342 148000
rect 7930 147200 7986 148000
rect 8574 147200 8630 148000
rect 9218 147200 9274 148000
rect 9862 147200 9918 148000
rect 10506 147200 10562 148000
rect 11150 147200 11206 148000
rect 11794 147200 11850 148000
rect 12438 147200 12494 148000
rect 13082 147200 13138 148000
rect 13726 147200 13782 148000
rect 14370 147200 14426 148000
rect 15014 147200 15070 148000
rect 15658 147200 15714 148000
rect 16302 147200 16358 148000
rect 16946 147200 17002 148000
rect 17590 147200 17646 148000
rect 18234 147200 18290 148000
rect 18878 147200 18934 148000
rect 19522 147200 19578 148000
rect 20166 147200 20222 148000
rect 20810 147200 20866 148000
rect 21454 147200 21510 148000
rect 22098 147200 22154 148000
rect 22742 147200 22798 148000
rect 23386 147200 23442 148000
rect 24030 147200 24086 148000
rect 24674 147200 24730 148000
rect 25318 147200 25374 148000
rect 25962 147200 26018 148000
rect 26606 147200 26662 148000
rect 27250 147200 27306 148000
rect 27894 147200 27950 148000
rect 28538 147200 28594 148000
rect 29182 147200 29238 148000
rect 29826 147200 29882 148000
rect 30470 147200 30526 148000
rect 31022 147200 31078 148000
rect 31666 147200 31722 148000
rect 32310 147200 32366 148000
rect 32954 147200 33010 148000
rect 33598 147200 33654 148000
rect 34242 147200 34298 148000
rect 34886 147200 34942 148000
rect 35530 147200 35586 148000
rect 36174 147200 36230 148000
rect 36818 147200 36874 148000
rect 37462 147200 37518 148000
rect 38106 147200 38162 148000
rect 38750 147200 38806 148000
rect 39394 147200 39450 148000
rect 40038 147200 40094 148000
rect 40682 147200 40738 148000
rect 41326 147200 41382 148000
rect 41970 147200 42026 148000
rect 42614 147200 42670 148000
rect 43258 147200 43314 148000
rect 43902 147200 43958 148000
rect 44546 147200 44602 148000
rect 45190 147200 45246 148000
rect 45834 147200 45890 148000
rect 46478 147200 46534 148000
rect 47122 147200 47178 148000
rect 47766 147200 47822 148000
rect 48410 147200 48466 148000
rect 49054 147200 49110 148000
rect 49698 147200 49754 148000
rect 50342 147200 50398 148000
rect 50986 147200 51042 148000
rect 51630 147200 51686 148000
rect 52274 147200 52330 148000
rect 52918 147200 52974 148000
rect 53562 147200 53618 148000
rect 54206 147200 54262 148000
rect 54850 147200 54906 148000
rect 55494 147200 55550 148000
rect 56138 147200 56194 148000
rect 56782 147200 56838 148000
rect 57426 147200 57482 148000
rect 58070 147200 58126 148000
rect 58714 147200 58770 148000
rect 59358 147200 59414 148000
rect 60002 147200 60058 148000
rect 60646 147200 60702 148000
rect 61290 147200 61346 148000
rect 61842 147200 61898 148000
rect 62486 147200 62542 148000
rect 63130 147200 63186 148000
rect 63774 147200 63830 148000
rect 64418 147200 64474 148000
rect 65062 147200 65118 148000
rect 65706 147200 65762 148000
rect 66350 147200 66406 148000
rect 66994 147200 67050 148000
rect 67638 147200 67694 148000
rect 68282 147200 68338 148000
rect 68926 147200 68982 148000
rect 69570 147200 69626 148000
rect 70214 147200 70270 148000
rect 70858 147200 70914 148000
rect 71502 147200 71558 148000
rect 72146 147200 72202 148000
rect 72790 147200 72846 148000
rect 73434 147200 73490 148000
rect 74078 147200 74134 148000
rect 74722 147200 74778 148000
rect 75366 147200 75422 148000
rect 76010 147200 76066 148000
rect 76654 147200 76710 148000
rect 77298 147200 77354 148000
rect 77942 147200 77998 148000
rect 78586 147200 78642 148000
rect 79230 147200 79286 148000
rect 79874 147200 79930 148000
rect 80518 147200 80574 148000
rect 81162 147200 81218 148000
rect 81806 147200 81862 148000
rect 82450 147200 82506 148000
rect 83094 147200 83150 148000
rect 83738 147200 83794 148000
rect 84382 147200 84438 148000
rect 85026 147200 85082 148000
rect 85670 147200 85726 148000
rect 86314 147200 86370 148000
rect 86958 147200 87014 148000
rect 87602 147200 87658 148000
rect 88246 147200 88302 148000
rect 88890 147200 88946 148000
rect 89534 147200 89590 148000
rect 90178 147200 90234 148000
rect 90822 147200 90878 148000
rect 91466 147200 91522 148000
rect 92110 147200 92166 148000
rect 92662 147200 92718 148000
rect 93306 147200 93362 148000
rect 93950 147200 94006 148000
rect 94594 147200 94650 148000
rect 95238 147200 95294 148000
rect 95882 147200 95938 148000
rect 96526 147200 96582 148000
rect 97170 147200 97226 148000
rect 97814 147200 97870 148000
rect 98458 147200 98514 148000
rect 99102 147200 99158 148000
rect 99746 147200 99802 148000
rect 100390 147200 100446 148000
rect 101034 147200 101090 148000
rect 101678 147200 101734 148000
rect 102322 147200 102378 148000
rect 102966 147200 103022 148000
rect 103610 147200 103666 148000
rect 104254 147200 104310 148000
rect 104898 147200 104954 148000
rect 105542 147200 105598 148000
rect 106186 147200 106242 148000
rect 106830 147200 106886 148000
rect 107474 147200 107530 148000
rect 108118 147200 108174 148000
rect 108762 147200 108818 148000
rect 109406 147200 109462 148000
rect 110050 147200 110106 148000
rect 110694 147200 110750 148000
rect 111338 147200 111394 148000
rect 111982 147200 112038 148000
rect 112626 147200 112682 148000
rect 113270 147200 113326 148000
rect 113914 147200 113970 148000
rect 114558 147200 114614 148000
rect 115202 147200 115258 148000
rect 115846 147200 115902 148000
rect 116490 147200 116546 148000
rect 117134 147200 117190 148000
rect 117778 147200 117834 148000
rect 118422 147200 118478 148000
rect 119066 147200 119122 148000
rect 119710 147200 119766 148000
rect 120354 147200 120410 148000
rect 120998 147200 121054 148000
rect 121642 147200 121698 148000
rect 122286 147200 122342 148000
rect 122930 147200 122986 148000
rect 123482 147200 123538 148000
rect 124126 147200 124182 148000
rect 124770 147200 124826 148000
rect 125414 147200 125470 148000
rect 126058 147200 126114 148000
rect 126702 147200 126758 148000
rect 127346 147200 127402 148000
rect 127990 147200 128046 148000
rect 128634 147200 128690 148000
rect 129278 147200 129334 148000
rect 129922 147200 129978 148000
rect 130566 147200 130622 148000
rect 131210 147200 131266 148000
rect 131854 147200 131910 148000
rect 132498 147200 132554 148000
rect 133142 147200 133198 148000
rect 133786 147200 133842 148000
rect 134430 147200 134486 148000
rect 135074 147200 135130 148000
rect 135718 147200 135774 148000
rect 136362 147200 136418 148000
rect 137006 147200 137062 148000
rect 137650 147200 137706 148000
rect 138294 147200 138350 148000
rect 138938 147200 138994 148000
rect 139582 147200 139638 148000
rect 140226 147200 140282 148000
rect 140870 147200 140926 148000
rect 141514 147200 141570 148000
rect 142158 147200 142214 148000
rect 142802 147200 142858 148000
rect 143446 147200 143502 148000
rect 144090 147200 144146 148000
rect 144734 147200 144790 148000
rect 145378 147200 145434 148000
rect 146022 147200 146078 148000
rect 146666 147200 146722 148000
rect 147310 147200 147366 148000
rect 147954 147200 148010 148000
rect 148598 147200 148654 148000
rect 149242 147200 149298 148000
rect 149886 147200 149942 148000
rect 150530 147200 150586 148000
rect 151174 147200 151230 148000
rect 151818 147200 151874 148000
rect 152462 147200 152518 148000
rect 153106 147200 153162 148000
rect 153750 147200 153806 148000
rect 154302 147200 154358 148000
rect 154946 147200 155002 148000
rect 155590 147200 155646 148000
rect 156234 147200 156290 148000
rect 156878 147200 156934 148000
rect 157522 147200 157578 148000
rect 158166 147200 158222 148000
rect 158810 147200 158866 148000
rect 159454 147200 159510 148000
rect 160098 147200 160154 148000
rect 160742 147200 160798 148000
rect 161386 147200 161442 148000
rect 162030 147200 162086 148000
rect 162674 147200 162730 148000
rect 163318 147200 163374 148000
rect 163962 147200 164018 148000
rect 164606 147200 164662 148000
rect 165250 147200 165306 148000
rect 165894 147200 165950 148000
rect 166538 147200 166594 148000
rect 167182 147200 167238 148000
rect 167826 147200 167882 148000
rect 168470 147200 168526 148000
rect 169114 147200 169170 148000
rect 169758 147200 169814 148000
rect 170402 147200 170458 148000
rect 171046 147200 171102 148000
rect 171690 147200 171746 148000
rect 172334 147200 172390 148000
rect 172978 147200 173034 148000
rect 173622 147200 173678 148000
rect 174266 147200 174322 148000
rect 174910 147200 174966 148000
rect 175554 147200 175610 148000
rect 176198 147200 176254 148000
rect 176842 147200 176898 148000
rect 177486 147200 177542 148000
rect 178130 147200 178186 148000
rect 178774 147200 178830 148000
rect 179418 147200 179474 148000
rect 180062 147200 180118 148000
rect 180706 147200 180762 148000
rect 181350 147200 181406 148000
rect 181994 147200 182050 148000
rect 182638 147200 182694 148000
rect 183282 147200 183338 148000
rect 183926 147200 183982 148000
rect 184570 147200 184626 148000
rect 185122 147200 185178 148000
rect 185766 147200 185822 148000
rect 186410 147200 186466 148000
rect 187054 147200 187110 148000
rect 187698 147200 187754 148000
rect 188342 147200 188398 148000
rect 188986 147200 189042 148000
rect 189630 147200 189686 148000
rect 190274 147200 190330 148000
rect 190918 147200 190974 148000
rect 191562 147200 191618 148000
rect 192206 147200 192262 148000
rect 192850 147200 192906 148000
rect 193494 147200 193550 148000
rect 194138 147200 194194 148000
rect 194782 147200 194838 148000
rect 195426 147200 195482 148000
rect 196070 147200 196126 148000
rect 196714 147200 196770 148000
rect 197358 147200 197414 148000
rect 198002 147200 198058 148000
rect 198646 147200 198702 148000
rect 199290 147200 199346 148000
rect 199934 147200 199990 148000
rect 200578 147200 200634 148000
rect 201222 147200 201278 148000
rect 201866 147200 201922 148000
rect 202510 147200 202566 148000
rect 203154 147200 203210 148000
rect 203798 147200 203854 148000
rect 204442 147200 204498 148000
rect 205086 147200 205142 148000
rect 205730 147200 205786 148000
rect 206374 147200 206430 148000
rect 207018 147200 207074 148000
rect 207662 147200 207718 148000
rect 208306 147200 208362 148000
rect 208950 147200 209006 148000
rect 209594 147200 209650 148000
rect 210238 147200 210294 148000
rect 210882 147200 210938 148000
rect 211526 147200 211582 148000
rect 212170 147200 212226 148000
rect 212814 147200 212870 148000
rect 213458 147200 213514 148000
rect 214102 147200 214158 148000
rect 214746 147200 214802 148000
rect 215390 147200 215446 148000
rect 215942 147200 215998 148000
rect 216586 147200 216642 148000
rect 217230 147200 217286 148000
rect 217874 147200 217930 148000
rect 218518 147200 218574 148000
rect 219162 147200 219218 148000
rect 219806 147200 219862 148000
rect 220450 147200 220506 148000
rect 221094 147200 221150 148000
rect 221738 147200 221794 148000
rect 222382 147200 222438 148000
rect 223026 147200 223082 148000
rect 223670 147200 223726 148000
rect 224314 147200 224370 148000
rect 224958 147200 225014 148000
rect 225602 147200 225658 148000
rect 226246 147200 226302 148000
rect 226890 147200 226946 148000
rect 227534 147200 227590 148000
rect 228178 147200 228234 148000
rect 228822 147200 228878 148000
rect 229466 147200 229522 148000
rect 230110 147200 230166 148000
rect 230754 147200 230810 148000
rect 231398 147200 231454 148000
rect 232042 147200 232098 148000
rect 232686 147200 232742 148000
rect 233330 147200 233386 148000
rect 233974 147200 234030 148000
rect 234618 147200 234674 148000
rect 235262 147200 235318 148000
rect 235906 147200 235962 148000
rect 236550 147200 236606 148000
rect 237194 147200 237250 148000
rect 237838 147200 237894 148000
rect 238482 147200 238538 148000
rect 239126 147200 239182 148000
rect 239770 147200 239826 148000
rect 240414 147200 240470 148000
rect 241058 147200 241114 148000
rect 241702 147200 241758 148000
rect 242346 147200 242402 148000
rect 242990 147200 243046 148000
rect 243634 147200 243690 148000
rect 244278 147200 244334 148000
rect 244922 147200 244978 148000
rect 245566 147200 245622 148000
rect 246210 147200 246266 148000
rect 246762 147200 246818 148000
rect 247406 147200 247462 148000
rect 248050 147200 248106 148000
rect 248694 147200 248750 148000
rect 249338 147200 249394 148000
rect 249982 147200 250038 148000
rect 250626 147200 250682 148000
rect 251270 147200 251326 148000
rect 251914 147200 251970 148000
rect 252558 147200 252614 148000
rect 253202 147200 253258 148000
rect 253846 147200 253902 148000
rect 254490 147200 254546 148000
rect 255134 147200 255190 148000
rect 255778 147200 255834 148000
rect 256422 147200 256478 148000
rect 257066 147200 257122 148000
rect 257710 147200 257766 148000
rect 258354 147200 258410 148000
rect 258998 147200 259054 148000
rect 259642 147200 259698 148000
rect 260286 147200 260342 148000
rect 260930 147200 260986 148000
rect 261574 147200 261630 148000
rect 262218 147200 262274 148000
rect 262862 147200 262918 148000
rect 263506 147200 263562 148000
rect 264150 147200 264206 148000
rect 264794 147200 264850 148000
rect 265438 147200 265494 148000
rect 266082 147200 266138 148000
rect 266726 147200 266782 148000
rect 267370 147200 267426 148000
rect 268014 147200 268070 148000
rect 268658 147200 268714 148000
rect 269302 147200 269358 148000
rect 269946 147200 270002 148000
rect 270590 147200 270646 148000
rect 271234 147200 271290 148000
rect 271878 147200 271934 148000
rect 272522 147200 272578 148000
rect 273166 147200 273222 148000
rect 273810 147200 273866 148000
rect 274454 147200 274510 148000
rect 275098 147200 275154 148000
rect 275742 147200 275798 148000
rect 276386 147200 276442 148000
rect 277030 147200 277086 148000
rect 277582 147200 277638 148000
rect 278226 147200 278282 148000
rect 278870 147200 278926 148000
rect 279514 147200 279570 148000
rect 280158 147200 280214 148000
rect 280802 147200 280858 148000
rect 281446 147200 281502 148000
rect 282090 147200 282146 148000
rect 282734 147200 282790 148000
rect 283378 147200 283434 148000
rect 284022 147200 284078 148000
rect 284666 147200 284722 148000
rect 285310 147200 285366 148000
rect 285954 147200 286010 148000
rect 286598 147200 286654 148000
rect 287242 147200 287298 148000
rect 287886 147200 287942 148000
rect 288530 147200 288586 148000
rect 289174 147200 289230 148000
rect 289818 147200 289874 148000
rect 290462 147200 290518 148000
rect 291106 147200 291162 148000
rect 291750 147200 291806 148000
rect 292394 147200 292450 148000
rect 293038 147200 293094 148000
rect 293682 147200 293738 148000
rect 294326 147200 294382 148000
rect 294970 147200 295026 148000
rect 295614 147200 295670 148000
rect 296258 147200 296314 148000
rect 296902 147200 296958 148000
rect 297546 147200 297602 148000
rect 298190 147200 298246 148000
rect 298834 147200 298890 148000
rect 299478 147200 299534 148000
rect 300122 147200 300178 148000
rect 300766 147200 300822 148000
rect 301410 147200 301466 148000
rect 302054 147200 302110 148000
rect 302698 147200 302754 148000
rect 303342 147200 303398 148000
rect 303986 147200 304042 148000
rect 304630 147200 304686 148000
rect 305274 147200 305330 148000
rect 305918 147200 305974 148000
rect 306562 147200 306618 148000
rect 307206 147200 307262 148000
rect 307850 147200 307906 148000
rect 308402 147200 308458 148000
rect 309046 147200 309102 148000
rect 309690 147200 309746 148000
rect 310334 147200 310390 148000
rect 310978 147200 311034 148000
rect 311622 147200 311678 148000
rect 312266 147200 312322 148000
rect 312910 147200 312966 148000
rect 313554 147200 313610 148000
rect 314198 147200 314254 148000
rect 314842 147200 314898 148000
rect 315486 147200 315542 148000
rect 316130 147200 316186 148000
rect 316774 147200 316830 148000
rect 317418 147200 317474 148000
rect 318062 147200 318118 148000
rect 318706 147200 318762 148000
rect 319350 147200 319406 148000
rect 319994 147200 320050 148000
rect 320638 147200 320694 148000
rect 321282 147200 321338 148000
rect 321926 147200 321982 148000
rect 322570 147200 322626 148000
rect 323214 147200 323270 148000
rect 323858 147200 323914 148000
rect 324502 147200 324558 148000
rect 325146 147200 325202 148000
rect 325790 147200 325846 148000
rect 326434 147200 326490 148000
rect 327078 147200 327134 148000
rect 327722 147200 327778 148000
rect 328366 147200 328422 148000
rect 329010 147200 329066 148000
rect 329654 147200 329710 148000
rect 330298 147200 330354 148000
rect 330942 147200 330998 148000
rect 331586 147200 331642 148000
rect 332230 147200 332286 148000
rect 332874 147200 332930 148000
rect 333518 147200 333574 148000
rect 334162 147200 334218 148000
rect 334806 147200 334862 148000
rect 335450 147200 335506 148000
rect 336094 147200 336150 148000
rect 336738 147200 336794 148000
rect 337382 147200 337438 148000
rect 338026 147200 338082 148000
rect 338670 147200 338726 148000
rect 339222 147200 339278 148000
rect 339866 147200 339922 148000
rect 340510 147200 340566 148000
rect 341154 147200 341210 148000
rect 341798 147200 341854 148000
rect 342442 147200 342498 148000
rect 343086 147200 343142 148000
rect 343730 147200 343786 148000
rect 344374 147200 344430 148000
rect 345018 147200 345074 148000
rect 345662 147200 345718 148000
rect 346306 147200 346362 148000
rect 346950 147200 347006 148000
rect 347594 147200 347650 148000
rect 348238 147200 348294 148000
rect 348882 147200 348938 148000
rect 349526 147200 349582 148000
rect 350170 147200 350226 148000
rect 350814 147200 350870 148000
rect 351458 147200 351514 148000
rect 352102 147200 352158 148000
rect 352746 147200 352802 148000
rect 353390 147200 353446 148000
rect 354034 147200 354090 148000
rect 354678 147200 354734 148000
rect 355322 147200 355378 148000
rect 355966 147200 356022 148000
rect 356610 147200 356666 148000
rect 357254 147200 357310 148000
rect 357898 147200 357954 148000
rect 358542 147200 358598 148000
rect 359186 147200 359242 148000
rect 359830 147200 359886 148000
rect 360474 147200 360530 148000
rect 361118 147200 361174 148000
rect 361762 147200 361818 148000
rect 362406 147200 362462 148000
rect 363050 147200 363106 148000
rect 363694 147200 363750 148000
rect 364338 147200 364394 148000
rect 364982 147200 365038 148000
rect 365626 147200 365682 148000
rect 366270 147200 366326 148000
rect 366914 147200 366970 148000
rect 367558 147200 367614 148000
rect 368202 147200 368258 148000
rect 368846 147200 368902 148000
rect 369490 147200 369546 148000
rect 370042 147200 370098 148000
rect 370686 147200 370742 148000
rect 371330 147200 371386 148000
rect 371974 147200 372030 148000
rect 372618 147200 372674 148000
rect 373262 147200 373318 148000
rect 373906 147200 373962 148000
rect 374550 147200 374606 148000
rect 375194 147200 375250 148000
rect 375838 147200 375894 148000
rect 376482 147200 376538 148000
rect 377126 147200 377182 148000
rect 377770 147200 377826 148000
rect 378414 147200 378470 148000
rect 379058 147200 379114 148000
rect 379702 147200 379758 148000
rect 380346 147200 380402 148000
rect 380990 147200 381046 148000
rect 381634 147200 381690 148000
rect 382278 147200 382334 148000
rect 382922 147200 382978 148000
rect 383566 147200 383622 148000
rect 384210 147200 384266 148000
rect 384854 147200 384910 148000
rect 385498 147200 385554 148000
rect 386142 147200 386198 148000
rect 386786 147200 386842 148000
rect 387430 147200 387486 148000
rect 388074 147200 388130 148000
rect 388718 147200 388774 148000
rect 389362 147200 389418 148000
rect 390006 147200 390062 148000
rect 390650 147200 390706 148000
rect 391294 147200 391350 148000
rect 391938 147200 391994 148000
rect 392582 147200 392638 148000
rect 393226 147200 393282 148000
rect 393870 147200 393926 148000
rect 394514 147200 394570 148000
rect 395158 147200 395214 148000
rect 395802 147200 395858 148000
rect 396446 147200 396502 148000
rect 397090 147200 397146 148000
rect 397734 147200 397790 148000
rect 398378 147200 398434 148000
rect 399022 147200 399078 148000
rect 399666 147200 399722 148000
rect 24950 0 25006 800
rect 74906 0 74962 800
rect 124954 0 125010 800
rect 174910 0 174966 800
rect 224958 0 225014 800
rect 274914 0 274970 800
rect 324962 0 325018 800
rect 374918 0 374974 800
<< obsm2 >>
rect 406 147144 790 147966
rect 958 147144 1434 147966
rect 1602 147144 2078 147966
rect 2246 147144 2722 147966
rect 2890 147144 3366 147966
rect 3534 147144 4010 147966
rect 4178 147144 4654 147966
rect 4822 147144 5298 147966
rect 5466 147144 5942 147966
rect 6110 147144 6586 147966
rect 6754 147144 7230 147966
rect 7398 147144 7874 147966
rect 8042 147144 8518 147966
rect 8686 147144 9162 147966
rect 9330 147144 9806 147966
rect 9974 147144 10450 147966
rect 10618 147144 11094 147966
rect 11262 147144 11738 147966
rect 11906 147144 12382 147966
rect 12550 147144 13026 147966
rect 13194 147144 13670 147966
rect 13838 147144 14314 147966
rect 14482 147144 14958 147966
rect 15126 147144 15602 147966
rect 15770 147144 16246 147966
rect 16414 147144 16890 147966
rect 17058 147144 17534 147966
rect 17702 147144 18178 147966
rect 18346 147144 18822 147966
rect 18990 147144 19466 147966
rect 19634 147144 20110 147966
rect 20278 147144 20754 147966
rect 20922 147144 21398 147966
rect 21566 147144 22042 147966
rect 22210 147144 22686 147966
rect 22854 147144 23330 147966
rect 23498 147144 23974 147966
rect 24142 147144 24618 147966
rect 24786 147144 25262 147966
rect 25430 147144 25906 147966
rect 26074 147144 26550 147966
rect 26718 147144 27194 147966
rect 27362 147144 27838 147966
rect 28006 147144 28482 147966
rect 28650 147144 29126 147966
rect 29294 147144 29770 147966
rect 29938 147144 30414 147966
rect 30582 147144 30966 147966
rect 31134 147144 31610 147966
rect 31778 147144 32254 147966
rect 32422 147144 32898 147966
rect 33066 147144 33542 147966
rect 33710 147144 34186 147966
rect 34354 147144 34830 147966
rect 34998 147144 35474 147966
rect 35642 147144 36118 147966
rect 36286 147144 36762 147966
rect 36930 147144 37406 147966
rect 37574 147144 38050 147966
rect 38218 147144 38694 147966
rect 38862 147144 39338 147966
rect 39506 147144 39982 147966
rect 40150 147144 40626 147966
rect 40794 147144 41270 147966
rect 41438 147144 41914 147966
rect 42082 147144 42558 147966
rect 42726 147144 43202 147966
rect 43370 147144 43846 147966
rect 44014 147144 44490 147966
rect 44658 147144 45134 147966
rect 45302 147144 45778 147966
rect 45946 147144 46422 147966
rect 46590 147144 47066 147966
rect 47234 147144 47710 147966
rect 47878 147144 48354 147966
rect 48522 147144 48998 147966
rect 49166 147144 49642 147966
rect 49810 147144 50286 147966
rect 50454 147144 50930 147966
rect 51098 147144 51574 147966
rect 51742 147144 52218 147966
rect 52386 147144 52862 147966
rect 53030 147144 53506 147966
rect 53674 147144 54150 147966
rect 54318 147144 54794 147966
rect 54962 147144 55438 147966
rect 55606 147144 56082 147966
rect 56250 147144 56726 147966
rect 56894 147144 57370 147966
rect 57538 147144 58014 147966
rect 58182 147144 58658 147966
rect 58826 147144 59302 147966
rect 59470 147144 59946 147966
rect 60114 147144 60590 147966
rect 60758 147144 61234 147966
rect 61402 147144 61786 147966
rect 61954 147144 62430 147966
rect 62598 147144 63074 147966
rect 63242 147144 63718 147966
rect 63886 147144 64362 147966
rect 64530 147144 65006 147966
rect 65174 147144 65650 147966
rect 65818 147144 66294 147966
rect 66462 147144 66938 147966
rect 67106 147144 67582 147966
rect 67750 147144 68226 147966
rect 68394 147144 68870 147966
rect 69038 147144 69514 147966
rect 69682 147144 70158 147966
rect 70326 147144 70802 147966
rect 70970 147144 71446 147966
rect 71614 147144 72090 147966
rect 72258 147144 72734 147966
rect 72902 147144 73378 147966
rect 73546 147144 74022 147966
rect 74190 147144 74666 147966
rect 74834 147144 75310 147966
rect 75478 147144 75954 147966
rect 76122 147144 76598 147966
rect 76766 147144 77242 147966
rect 77410 147144 77886 147966
rect 78054 147144 78530 147966
rect 78698 147144 79174 147966
rect 79342 147144 79818 147966
rect 79986 147144 80462 147966
rect 80630 147144 81106 147966
rect 81274 147144 81750 147966
rect 81918 147144 82394 147966
rect 82562 147144 83038 147966
rect 83206 147144 83682 147966
rect 83850 147144 84326 147966
rect 84494 147144 84970 147966
rect 85138 147144 85614 147966
rect 85782 147144 86258 147966
rect 86426 147144 86902 147966
rect 87070 147144 87546 147966
rect 87714 147144 88190 147966
rect 88358 147144 88834 147966
rect 89002 147144 89478 147966
rect 89646 147144 90122 147966
rect 90290 147144 90766 147966
rect 90934 147144 91410 147966
rect 91578 147144 92054 147966
rect 92222 147144 92606 147966
rect 92774 147144 93250 147966
rect 93418 147144 93894 147966
rect 94062 147144 94538 147966
rect 94706 147144 95182 147966
rect 95350 147144 95826 147966
rect 95994 147144 96470 147966
rect 96638 147144 97114 147966
rect 97282 147144 97758 147966
rect 97926 147144 98402 147966
rect 98570 147144 99046 147966
rect 99214 147144 99690 147966
rect 99858 147144 100334 147966
rect 100502 147144 100978 147966
rect 101146 147144 101622 147966
rect 101790 147144 102266 147966
rect 102434 147144 102910 147966
rect 103078 147144 103554 147966
rect 103722 147144 104198 147966
rect 104366 147144 104842 147966
rect 105010 147144 105486 147966
rect 105654 147144 106130 147966
rect 106298 147144 106774 147966
rect 106942 147144 107418 147966
rect 107586 147144 108062 147966
rect 108230 147144 108706 147966
rect 108874 147144 109350 147966
rect 109518 147144 109994 147966
rect 110162 147144 110638 147966
rect 110806 147144 111282 147966
rect 111450 147144 111926 147966
rect 112094 147144 112570 147966
rect 112738 147144 113214 147966
rect 113382 147144 113858 147966
rect 114026 147144 114502 147966
rect 114670 147144 115146 147966
rect 115314 147144 115790 147966
rect 115958 147144 116434 147966
rect 116602 147144 117078 147966
rect 117246 147144 117722 147966
rect 117890 147144 118366 147966
rect 118534 147144 119010 147966
rect 119178 147144 119654 147966
rect 119822 147144 120298 147966
rect 120466 147144 120942 147966
rect 121110 147144 121586 147966
rect 121754 147144 122230 147966
rect 122398 147144 122874 147966
rect 123042 147144 123426 147966
rect 123594 147144 124070 147966
rect 124238 147144 124714 147966
rect 124882 147144 125358 147966
rect 125526 147144 126002 147966
rect 126170 147144 126646 147966
rect 126814 147144 127290 147966
rect 127458 147144 127934 147966
rect 128102 147144 128578 147966
rect 128746 147144 129222 147966
rect 129390 147144 129866 147966
rect 130034 147144 130510 147966
rect 130678 147144 131154 147966
rect 131322 147144 131798 147966
rect 131966 147144 132442 147966
rect 132610 147144 133086 147966
rect 133254 147144 133730 147966
rect 133898 147144 134374 147966
rect 134542 147144 135018 147966
rect 135186 147144 135662 147966
rect 135830 147144 136306 147966
rect 136474 147144 136950 147966
rect 137118 147144 137594 147966
rect 137762 147144 138238 147966
rect 138406 147144 138882 147966
rect 139050 147144 139526 147966
rect 139694 147144 140170 147966
rect 140338 147144 140814 147966
rect 140982 147144 141458 147966
rect 141626 147144 142102 147966
rect 142270 147144 142746 147966
rect 142914 147144 143390 147966
rect 143558 147144 144034 147966
rect 144202 147144 144678 147966
rect 144846 147144 145322 147966
rect 145490 147144 145966 147966
rect 146134 147144 146610 147966
rect 146778 147144 147254 147966
rect 147422 147144 147898 147966
rect 148066 147144 148542 147966
rect 148710 147144 149186 147966
rect 149354 147144 149830 147966
rect 149998 147144 150474 147966
rect 150642 147144 151118 147966
rect 151286 147144 151762 147966
rect 151930 147144 152406 147966
rect 152574 147144 153050 147966
rect 153218 147144 153694 147966
rect 153862 147144 154246 147966
rect 154414 147144 154890 147966
rect 155058 147144 155534 147966
rect 155702 147144 156178 147966
rect 156346 147144 156822 147966
rect 156990 147144 157466 147966
rect 157634 147144 158110 147966
rect 158278 147144 158754 147966
rect 158922 147144 159398 147966
rect 159566 147144 160042 147966
rect 160210 147144 160686 147966
rect 160854 147144 161330 147966
rect 161498 147144 161974 147966
rect 162142 147144 162618 147966
rect 162786 147144 163262 147966
rect 163430 147144 163906 147966
rect 164074 147144 164550 147966
rect 164718 147144 165194 147966
rect 165362 147144 165838 147966
rect 166006 147144 166482 147966
rect 166650 147144 167126 147966
rect 167294 147144 167770 147966
rect 167938 147144 168414 147966
rect 168582 147144 169058 147966
rect 169226 147144 169702 147966
rect 169870 147144 170346 147966
rect 170514 147144 170990 147966
rect 171158 147144 171634 147966
rect 171802 147144 172278 147966
rect 172446 147144 172922 147966
rect 173090 147144 173566 147966
rect 173734 147144 174210 147966
rect 174378 147144 174854 147966
rect 175022 147144 175498 147966
rect 175666 147144 176142 147966
rect 176310 147144 176786 147966
rect 176954 147144 177430 147966
rect 177598 147144 178074 147966
rect 178242 147144 178718 147966
rect 178886 147144 179362 147966
rect 179530 147144 180006 147966
rect 180174 147144 180650 147966
rect 180818 147144 181294 147966
rect 181462 147144 181938 147966
rect 182106 147144 182582 147966
rect 182750 147144 183226 147966
rect 183394 147144 183870 147966
rect 184038 147144 184514 147966
rect 184682 147144 185066 147966
rect 185234 147144 185710 147966
rect 185878 147144 186354 147966
rect 186522 147144 186998 147966
rect 187166 147144 187642 147966
rect 187810 147144 188286 147966
rect 188454 147144 188930 147966
rect 189098 147144 189574 147966
rect 189742 147144 190218 147966
rect 190386 147144 190862 147966
rect 191030 147144 191506 147966
rect 191674 147144 192150 147966
rect 192318 147144 192794 147966
rect 192962 147144 193438 147966
rect 193606 147144 194082 147966
rect 194250 147144 194726 147966
rect 194894 147144 195370 147966
rect 195538 147144 196014 147966
rect 196182 147144 196658 147966
rect 196826 147144 197302 147966
rect 197470 147144 197946 147966
rect 198114 147144 198590 147966
rect 198758 147144 199234 147966
rect 199402 147144 199878 147966
rect 200046 147144 200522 147966
rect 200690 147144 201166 147966
rect 201334 147144 201810 147966
rect 201978 147144 202454 147966
rect 202622 147144 203098 147966
rect 203266 147144 203742 147966
rect 203910 147144 204386 147966
rect 204554 147144 205030 147966
rect 205198 147144 205674 147966
rect 205842 147144 206318 147966
rect 206486 147144 206962 147966
rect 207130 147144 207606 147966
rect 207774 147144 208250 147966
rect 208418 147144 208894 147966
rect 209062 147144 209538 147966
rect 209706 147144 210182 147966
rect 210350 147144 210826 147966
rect 210994 147144 211470 147966
rect 211638 147144 212114 147966
rect 212282 147144 212758 147966
rect 212926 147144 213402 147966
rect 213570 147144 214046 147966
rect 214214 147144 214690 147966
rect 214858 147144 215334 147966
rect 215502 147144 215886 147966
rect 216054 147144 216530 147966
rect 216698 147144 217174 147966
rect 217342 147144 217818 147966
rect 217986 147144 218462 147966
rect 218630 147144 219106 147966
rect 219274 147144 219750 147966
rect 219918 147144 220394 147966
rect 220562 147144 221038 147966
rect 221206 147144 221682 147966
rect 221850 147144 222326 147966
rect 222494 147144 222970 147966
rect 223138 147144 223614 147966
rect 223782 147144 224258 147966
rect 224426 147144 224902 147966
rect 225070 147144 225546 147966
rect 225714 147144 226190 147966
rect 226358 147144 226834 147966
rect 227002 147144 227478 147966
rect 227646 147144 228122 147966
rect 228290 147144 228766 147966
rect 228934 147144 229410 147966
rect 229578 147144 230054 147966
rect 230222 147144 230698 147966
rect 230866 147144 231342 147966
rect 231510 147144 231986 147966
rect 232154 147144 232630 147966
rect 232798 147144 233274 147966
rect 233442 147144 233918 147966
rect 234086 147144 234562 147966
rect 234730 147144 235206 147966
rect 235374 147144 235850 147966
rect 236018 147144 236494 147966
rect 236662 147144 237138 147966
rect 237306 147144 237782 147966
rect 237950 147144 238426 147966
rect 238594 147144 239070 147966
rect 239238 147144 239714 147966
rect 239882 147144 240358 147966
rect 240526 147144 241002 147966
rect 241170 147144 241646 147966
rect 241814 147144 242290 147966
rect 242458 147144 242934 147966
rect 243102 147144 243578 147966
rect 243746 147144 244222 147966
rect 244390 147144 244866 147966
rect 245034 147144 245510 147966
rect 245678 147144 246154 147966
rect 246322 147144 246706 147966
rect 246874 147144 247350 147966
rect 247518 147144 247994 147966
rect 248162 147144 248638 147966
rect 248806 147144 249282 147966
rect 249450 147144 249926 147966
rect 250094 147144 250570 147966
rect 250738 147144 251214 147966
rect 251382 147144 251858 147966
rect 252026 147144 252502 147966
rect 252670 147144 253146 147966
rect 253314 147144 253790 147966
rect 253958 147144 254434 147966
rect 254602 147144 255078 147966
rect 255246 147144 255722 147966
rect 255890 147144 256366 147966
rect 256534 147144 257010 147966
rect 257178 147144 257654 147966
rect 257822 147144 258298 147966
rect 258466 147144 258942 147966
rect 259110 147144 259586 147966
rect 259754 147144 260230 147966
rect 260398 147144 260874 147966
rect 261042 147144 261518 147966
rect 261686 147144 262162 147966
rect 262330 147144 262806 147966
rect 262974 147144 263450 147966
rect 263618 147144 264094 147966
rect 264262 147144 264738 147966
rect 264906 147144 265382 147966
rect 265550 147144 266026 147966
rect 266194 147144 266670 147966
rect 266838 147144 267314 147966
rect 267482 147144 267958 147966
rect 268126 147144 268602 147966
rect 268770 147144 269246 147966
rect 269414 147144 269890 147966
rect 270058 147144 270534 147966
rect 270702 147144 271178 147966
rect 271346 147144 271822 147966
rect 271990 147144 272466 147966
rect 272634 147144 273110 147966
rect 273278 147144 273754 147966
rect 273922 147144 274398 147966
rect 274566 147144 275042 147966
rect 275210 147144 275686 147966
rect 275854 147144 276330 147966
rect 276498 147144 276974 147966
rect 277142 147144 277526 147966
rect 277694 147144 278170 147966
rect 278338 147144 278814 147966
rect 278982 147144 279458 147966
rect 279626 147144 280102 147966
rect 280270 147144 280746 147966
rect 280914 147144 281390 147966
rect 281558 147144 282034 147966
rect 282202 147144 282678 147966
rect 282846 147144 283322 147966
rect 283490 147144 283966 147966
rect 284134 147144 284610 147966
rect 284778 147144 285254 147966
rect 285422 147144 285898 147966
rect 286066 147144 286542 147966
rect 286710 147144 287186 147966
rect 287354 147144 287830 147966
rect 287998 147144 288474 147966
rect 288642 147144 289118 147966
rect 289286 147144 289762 147966
rect 289930 147144 290406 147966
rect 290574 147144 291050 147966
rect 291218 147144 291694 147966
rect 291862 147144 292338 147966
rect 292506 147144 292982 147966
rect 293150 147144 293626 147966
rect 293794 147144 294270 147966
rect 294438 147144 294914 147966
rect 295082 147144 295558 147966
rect 295726 147144 296202 147966
rect 296370 147144 296846 147966
rect 297014 147144 297490 147966
rect 297658 147144 298134 147966
rect 298302 147144 298778 147966
rect 298946 147144 299422 147966
rect 299590 147144 300066 147966
rect 300234 147144 300710 147966
rect 300878 147144 301354 147966
rect 301522 147144 301998 147966
rect 302166 147144 302642 147966
rect 302810 147144 303286 147966
rect 303454 147144 303930 147966
rect 304098 147144 304574 147966
rect 304742 147144 305218 147966
rect 305386 147144 305862 147966
rect 306030 147144 306506 147966
rect 306674 147144 307150 147966
rect 307318 147144 307794 147966
rect 307962 147144 308346 147966
rect 308514 147144 308990 147966
rect 309158 147144 309634 147966
rect 309802 147144 310278 147966
rect 310446 147144 310922 147966
rect 311090 147144 311566 147966
rect 311734 147144 312210 147966
rect 312378 147144 312854 147966
rect 313022 147144 313498 147966
rect 313666 147144 314142 147966
rect 314310 147144 314786 147966
rect 314954 147144 315430 147966
rect 315598 147144 316074 147966
rect 316242 147144 316718 147966
rect 316886 147144 317362 147966
rect 317530 147144 318006 147966
rect 318174 147144 318650 147966
rect 318818 147144 319294 147966
rect 319462 147144 319938 147966
rect 320106 147144 320582 147966
rect 320750 147144 321226 147966
rect 321394 147144 321870 147966
rect 322038 147144 322514 147966
rect 322682 147144 323158 147966
rect 323326 147144 323802 147966
rect 323970 147144 324446 147966
rect 324614 147144 325090 147966
rect 325258 147144 325734 147966
rect 325902 147144 326378 147966
rect 326546 147144 327022 147966
rect 327190 147144 327666 147966
rect 327834 147144 328310 147966
rect 328478 147144 328954 147966
rect 329122 147144 329598 147966
rect 329766 147144 330242 147966
rect 330410 147144 330886 147966
rect 331054 147144 331530 147966
rect 331698 147144 332174 147966
rect 332342 147144 332818 147966
rect 332986 147144 333462 147966
rect 333630 147144 334106 147966
rect 334274 147144 334750 147966
rect 334918 147144 335394 147966
rect 335562 147144 336038 147966
rect 336206 147144 336682 147966
rect 336850 147144 337326 147966
rect 337494 147144 337970 147966
rect 338138 147144 338614 147966
rect 338782 147144 339166 147966
rect 339334 147144 339810 147966
rect 339978 147144 340454 147966
rect 340622 147144 341098 147966
rect 341266 147144 341742 147966
rect 341910 147144 342386 147966
rect 342554 147144 343030 147966
rect 343198 147144 343674 147966
rect 343842 147144 344318 147966
rect 344486 147144 344962 147966
rect 345130 147144 345606 147966
rect 345774 147144 346250 147966
rect 346418 147144 346894 147966
rect 347062 147144 347538 147966
rect 347706 147144 348182 147966
rect 348350 147144 348826 147966
rect 348994 147144 349470 147966
rect 349638 147144 350114 147966
rect 350282 147144 350758 147966
rect 350926 147144 351402 147966
rect 351570 147144 352046 147966
rect 352214 147144 352690 147966
rect 352858 147144 353334 147966
rect 353502 147144 353978 147966
rect 354146 147144 354622 147966
rect 354790 147144 355266 147966
rect 355434 147144 355910 147966
rect 356078 147144 356554 147966
rect 356722 147144 357198 147966
rect 357366 147144 357842 147966
rect 358010 147144 358486 147966
rect 358654 147144 359130 147966
rect 359298 147144 359774 147966
rect 359942 147144 360418 147966
rect 360586 147144 361062 147966
rect 361230 147144 361706 147966
rect 361874 147144 362350 147966
rect 362518 147144 362994 147966
rect 363162 147144 363638 147966
rect 363806 147144 364282 147966
rect 364450 147144 364926 147966
rect 365094 147144 365570 147966
rect 365738 147144 366214 147966
rect 366382 147144 366858 147966
rect 367026 147144 367502 147966
rect 367670 147144 368146 147966
rect 368314 147144 368790 147966
rect 368958 147144 369434 147966
rect 369602 147144 369986 147966
rect 370154 147144 370630 147966
rect 370798 147144 371274 147966
rect 371442 147144 371918 147966
rect 372086 147144 372562 147966
rect 372730 147144 373206 147966
rect 373374 147144 373850 147966
rect 374018 147144 374494 147966
rect 374662 147144 375138 147966
rect 375306 147144 375782 147966
rect 375950 147144 376426 147966
rect 376594 147144 377070 147966
rect 377238 147144 377714 147966
rect 377882 147144 378358 147966
rect 378526 147144 379002 147966
rect 379170 147144 379646 147966
rect 379814 147144 380290 147966
rect 380458 147144 380934 147966
rect 381102 147144 381578 147966
rect 381746 147144 382222 147966
rect 382390 147144 382866 147966
rect 383034 147144 383510 147966
rect 383678 147144 384154 147966
rect 384322 147144 384798 147966
rect 384966 147144 385442 147966
rect 385610 147144 386086 147966
rect 386254 147144 386730 147966
rect 386898 147144 387374 147966
rect 387542 147144 388018 147966
rect 388186 147144 388662 147966
rect 388830 147144 389306 147966
rect 389474 147144 389950 147966
rect 390118 147144 390594 147966
rect 390762 147144 391238 147966
rect 391406 147144 391882 147966
rect 392050 147144 392526 147966
rect 392694 147144 393170 147966
rect 393338 147144 393814 147966
rect 393982 147144 394458 147966
rect 394626 147144 395102 147966
rect 395270 147144 395746 147966
rect 395914 147144 396390 147966
rect 396558 147144 397034 147966
rect 397202 147144 397678 147966
rect 397846 147144 398322 147966
rect 398490 147144 398966 147966
rect 399134 147144 399610 147966
rect 296 856 399720 147144
rect 296 711 24894 856
rect 25062 711 74850 856
rect 75018 711 124898 856
rect 125066 711 174854 856
rect 175022 711 224902 856
rect 225070 711 274858 856
rect 275026 711 324906 856
rect 325074 711 374862 856
rect 375030 711 399720 856
<< metal3 >>
rect 399200 147160 400000 147280
rect 0 146888 800 147008
rect 399200 145800 400000 145920
rect 0 144984 800 145104
rect 399200 144440 400000 144560
rect 0 143080 800 143200
rect 399200 143080 400000 143200
rect 399200 141720 400000 141840
rect 0 141176 800 141296
rect 399200 140360 400000 140480
rect 0 139272 800 139392
rect 399200 139000 400000 139120
rect 399200 137640 400000 137760
rect 0 137368 800 137488
rect 399200 136280 400000 136400
rect 0 135464 800 135584
rect 399200 134920 400000 135040
rect 0 133424 800 133544
rect 399200 133560 400000 133680
rect 399200 132200 400000 132320
rect 0 131520 800 131640
rect 399200 130840 400000 130960
rect 0 129616 800 129736
rect 399200 129344 400000 129464
rect 399200 127984 400000 128104
rect 0 127712 800 127832
rect 399200 126624 400000 126744
rect 0 125808 800 125928
rect 399200 125264 400000 125384
rect 0 123904 800 124024
rect 399200 123904 400000 124024
rect 399200 122544 400000 122664
rect 0 122000 800 122120
rect 399200 121184 400000 121304
rect 0 120096 800 120216
rect 399200 119824 400000 119944
rect 399200 118464 400000 118584
rect 0 118056 800 118176
rect 399200 117104 400000 117224
rect 0 116152 800 116272
rect 399200 115744 400000 115864
rect 0 114248 800 114368
rect 399200 114384 400000 114504
rect 399200 113024 400000 113144
rect 0 112344 800 112464
rect 399200 111664 400000 111784
rect 0 110440 800 110560
rect 399200 110168 400000 110288
rect 399200 108808 400000 108928
rect 0 108536 800 108656
rect 399200 107448 400000 107568
rect 0 106632 800 106752
rect 399200 106088 400000 106208
rect 0 104728 800 104848
rect 399200 104728 400000 104848
rect 399200 103368 400000 103488
rect 0 102688 800 102808
rect 399200 102008 400000 102128
rect 0 100784 800 100904
rect 399200 100648 400000 100768
rect 399200 99288 400000 99408
rect 0 98880 800 99000
rect 399200 97928 400000 98048
rect 0 96976 800 97096
rect 399200 96568 400000 96688
rect 0 95072 800 95192
rect 399200 95208 400000 95328
rect 399200 93848 400000 93968
rect 0 93168 800 93288
rect 399200 92352 400000 92472
rect 0 91264 800 91384
rect 399200 90992 400000 91112
rect 399200 89632 400000 89752
rect 0 89224 800 89344
rect 399200 88272 400000 88392
rect 0 87320 800 87440
rect 399200 86912 400000 87032
rect 0 85416 800 85536
rect 399200 85552 400000 85672
rect 399200 84192 400000 84312
rect 0 83512 800 83632
rect 399200 82832 400000 82952
rect 0 81608 800 81728
rect 399200 81472 400000 81592
rect 399200 80112 400000 80232
rect 0 79704 800 79824
rect 399200 78752 400000 78872
rect 0 77800 800 77920
rect 399200 77392 400000 77512
rect 0 75896 800 76016
rect 399200 76032 400000 76152
rect 399200 74672 400000 74792
rect 0 73856 800 73976
rect 399200 73176 400000 73296
rect 0 71952 800 72072
rect 399200 71816 400000 71936
rect 399200 70456 400000 70576
rect 0 70048 800 70168
rect 399200 69096 400000 69216
rect 0 68144 800 68264
rect 399200 67736 400000 67856
rect 0 66240 800 66360
rect 399200 66376 400000 66496
rect 399200 65016 400000 65136
rect 0 64336 800 64456
rect 399200 63656 400000 63776
rect 0 62432 800 62552
rect 399200 62296 400000 62416
rect 399200 60936 400000 61056
rect 0 60528 800 60648
rect 399200 59576 400000 59696
rect 0 58488 800 58608
rect 399200 58216 400000 58336
rect 399200 56856 400000 56976
rect 0 56584 800 56704
rect 399200 55360 400000 55480
rect 0 54680 800 54800
rect 399200 54000 400000 54120
rect 0 52776 800 52896
rect 399200 52640 400000 52760
rect 399200 51280 400000 51400
rect 0 50872 800 50992
rect 399200 49920 400000 50040
rect 0 48968 800 49088
rect 399200 48560 400000 48680
rect 0 47064 800 47184
rect 399200 47200 400000 47320
rect 399200 45840 400000 45960
rect 0 45024 800 45144
rect 399200 44480 400000 44600
rect 0 43120 800 43240
rect 399200 43120 400000 43240
rect 399200 41760 400000 41880
rect 0 41216 800 41336
rect 399200 40400 400000 40520
rect 0 39312 800 39432
rect 399200 39040 400000 39160
rect 399200 37680 400000 37800
rect 0 37408 800 37528
rect 399200 36184 400000 36304
rect 0 35504 800 35624
rect 399200 34824 400000 34944
rect 0 33600 800 33720
rect 399200 33464 400000 33584
rect 399200 32104 400000 32224
rect 0 31696 800 31816
rect 399200 30744 400000 30864
rect 0 29656 800 29776
rect 399200 29384 400000 29504
rect 399200 28024 400000 28144
rect 0 27752 800 27872
rect 399200 26664 400000 26784
rect 0 25848 800 25968
rect 399200 25304 400000 25424
rect 0 23944 800 24064
rect 399200 23944 400000 24064
rect 399200 22584 400000 22704
rect 0 22040 800 22160
rect 399200 21224 400000 21344
rect 0 20136 800 20256
rect 399200 19864 400000 19984
rect 0 18232 800 18352
rect 399200 18368 400000 18488
rect 399200 17008 400000 17128
rect 0 16328 800 16448
rect 399200 15648 400000 15768
rect 0 14288 800 14408
rect 399200 14288 400000 14408
rect 399200 12928 400000 13048
rect 0 12384 800 12504
rect 399200 11568 400000 11688
rect 0 10480 800 10600
rect 399200 10208 400000 10328
rect 399200 8848 400000 8968
rect 0 8576 800 8696
rect 399200 7488 400000 7608
rect 0 6672 800 6792
rect 399200 6128 400000 6248
rect 0 4768 800 4888
rect 399200 4768 400000 4888
rect 399200 3408 400000 3528
rect 0 2864 800 2984
rect 399200 2048 400000 2168
rect 0 960 800 1080
rect 399200 688 400000 808
<< obsm3 >>
rect 800 147360 399200 147389
rect 800 147088 399120 147360
rect 880 147080 399120 147088
rect 880 146808 399200 147080
rect 800 146000 399200 146808
rect 800 145720 399120 146000
rect 800 145184 399200 145720
rect 880 144904 399200 145184
rect 800 144640 399200 144904
rect 800 144360 399120 144640
rect 800 143280 399200 144360
rect 880 143000 399120 143280
rect 800 141920 399200 143000
rect 800 141640 399120 141920
rect 800 141376 399200 141640
rect 880 141096 399200 141376
rect 800 140560 399200 141096
rect 800 140280 399120 140560
rect 800 139472 399200 140280
rect 880 139200 399200 139472
rect 880 139192 399120 139200
rect 800 138920 399120 139192
rect 800 137840 399200 138920
rect 800 137568 399120 137840
rect 880 137560 399120 137568
rect 880 137288 399200 137560
rect 800 136480 399200 137288
rect 800 136200 399120 136480
rect 800 135664 399200 136200
rect 880 135384 399200 135664
rect 800 135120 399200 135384
rect 800 134840 399120 135120
rect 800 133760 399200 134840
rect 800 133624 399120 133760
rect 880 133480 399120 133624
rect 880 133344 399200 133480
rect 800 132400 399200 133344
rect 800 132120 399120 132400
rect 800 131720 399200 132120
rect 880 131440 399200 131720
rect 800 131040 399200 131440
rect 800 130760 399120 131040
rect 800 129816 399200 130760
rect 880 129544 399200 129816
rect 880 129536 399120 129544
rect 800 129264 399120 129536
rect 800 128184 399200 129264
rect 800 127912 399120 128184
rect 880 127904 399120 127912
rect 880 127632 399200 127904
rect 800 126824 399200 127632
rect 800 126544 399120 126824
rect 800 126008 399200 126544
rect 880 125728 399200 126008
rect 800 125464 399200 125728
rect 800 125184 399120 125464
rect 800 124104 399200 125184
rect 880 123824 399120 124104
rect 800 122744 399200 123824
rect 800 122464 399120 122744
rect 800 122200 399200 122464
rect 880 121920 399200 122200
rect 800 121384 399200 121920
rect 800 121104 399120 121384
rect 800 120296 399200 121104
rect 880 120024 399200 120296
rect 880 120016 399120 120024
rect 800 119744 399120 120016
rect 800 118664 399200 119744
rect 800 118384 399120 118664
rect 800 118256 399200 118384
rect 880 117976 399200 118256
rect 800 117304 399200 117976
rect 800 117024 399120 117304
rect 800 116352 399200 117024
rect 880 116072 399200 116352
rect 800 115944 399200 116072
rect 800 115664 399120 115944
rect 800 114584 399200 115664
rect 800 114448 399120 114584
rect 880 114304 399120 114448
rect 880 114168 399200 114304
rect 800 113224 399200 114168
rect 800 112944 399120 113224
rect 800 112544 399200 112944
rect 880 112264 399200 112544
rect 800 111864 399200 112264
rect 800 111584 399120 111864
rect 800 110640 399200 111584
rect 880 110368 399200 110640
rect 880 110360 399120 110368
rect 800 110088 399120 110360
rect 800 109008 399200 110088
rect 800 108736 399120 109008
rect 880 108728 399120 108736
rect 880 108456 399200 108728
rect 800 107648 399200 108456
rect 800 107368 399120 107648
rect 800 106832 399200 107368
rect 880 106552 399200 106832
rect 800 106288 399200 106552
rect 800 106008 399120 106288
rect 800 104928 399200 106008
rect 880 104648 399120 104928
rect 800 103568 399200 104648
rect 800 103288 399120 103568
rect 800 102888 399200 103288
rect 880 102608 399200 102888
rect 800 102208 399200 102608
rect 800 101928 399120 102208
rect 800 100984 399200 101928
rect 880 100848 399200 100984
rect 880 100704 399120 100848
rect 800 100568 399120 100704
rect 800 99488 399200 100568
rect 800 99208 399120 99488
rect 800 99080 399200 99208
rect 880 98800 399200 99080
rect 800 98128 399200 98800
rect 800 97848 399120 98128
rect 800 97176 399200 97848
rect 880 96896 399200 97176
rect 800 96768 399200 96896
rect 800 96488 399120 96768
rect 800 95408 399200 96488
rect 800 95272 399120 95408
rect 880 95128 399120 95272
rect 880 94992 399200 95128
rect 800 94048 399200 94992
rect 800 93768 399120 94048
rect 800 93368 399200 93768
rect 880 93088 399200 93368
rect 800 92552 399200 93088
rect 800 92272 399120 92552
rect 800 91464 399200 92272
rect 880 91192 399200 91464
rect 880 91184 399120 91192
rect 800 90912 399120 91184
rect 800 89832 399200 90912
rect 800 89552 399120 89832
rect 800 89424 399200 89552
rect 880 89144 399200 89424
rect 800 88472 399200 89144
rect 800 88192 399120 88472
rect 800 87520 399200 88192
rect 880 87240 399200 87520
rect 800 87112 399200 87240
rect 800 86832 399120 87112
rect 800 85752 399200 86832
rect 800 85616 399120 85752
rect 880 85472 399120 85616
rect 880 85336 399200 85472
rect 800 84392 399200 85336
rect 800 84112 399120 84392
rect 800 83712 399200 84112
rect 880 83432 399200 83712
rect 800 83032 399200 83432
rect 800 82752 399120 83032
rect 800 81808 399200 82752
rect 880 81672 399200 81808
rect 880 81528 399120 81672
rect 800 81392 399120 81528
rect 800 80312 399200 81392
rect 800 80032 399120 80312
rect 800 79904 399200 80032
rect 880 79624 399200 79904
rect 800 78952 399200 79624
rect 800 78672 399120 78952
rect 800 78000 399200 78672
rect 880 77720 399200 78000
rect 800 77592 399200 77720
rect 800 77312 399120 77592
rect 800 76232 399200 77312
rect 800 76096 399120 76232
rect 880 75952 399120 76096
rect 880 75816 399200 75952
rect 800 74872 399200 75816
rect 800 74592 399120 74872
rect 800 74056 399200 74592
rect 880 73776 399200 74056
rect 800 73376 399200 73776
rect 800 73096 399120 73376
rect 800 72152 399200 73096
rect 880 72016 399200 72152
rect 880 71872 399120 72016
rect 800 71736 399120 71872
rect 800 70656 399200 71736
rect 800 70376 399120 70656
rect 800 70248 399200 70376
rect 880 69968 399200 70248
rect 800 69296 399200 69968
rect 800 69016 399120 69296
rect 800 68344 399200 69016
rect 880 68064 399200 68344
rect 800 67936 399200 68064
rect 800 67656 399120 67936
rect 800 66576 399200 67656
rect 800 66440 399120 66576
rect 880 66296 399120 66440
rect 880 66160 399200 66296
rect 800 65216 399200 66160
rect 800 64936 399120 65216
rect 800 64536 399200 64936
rect 880 64256 399200 64536
rect 800 63856 399200 64256
rect 800 63576 399120 63856
rect 800 62632 399200 63576
rect 880 62496 399200 62632
rect 880 62352 399120 62496
rect 800 62216 399120 62352
rect 800 61136 399200 62216
rect 800 60856 399120 61136
rect 800 60728 399200 60856
rect 880 60448 399200 60728
rect 800 59776 399200 60448
rect 800 59496 399120 59776
rect 800 58688 399200 59496
rect 880 58416 399200 58688
rect 880 58408 399120 58416
rect 800 58136 399120 58408
rect 800 57056 399200 58136
rect 800 56784 399120 57056
rect 880 56776 399120 56784
rect 880 56504 399200 56776
rect 800 55560 399200 56504
rect 800 55280 399120 55560
rect 800 54880 399200 55280
rect 880 54600 399200 54880
rect 800 54200 399200 54600
rect 800 53920 399120 54200
rect 800 52976 399200 53920
rect 880 52840 399200 52976
rect 880 52696 399120 52840
rect 800 52560 399120 52696
rect 800 51480 399200 52560
rect 800 51200 399120 51480
rect 800 51072 399200 51200
rect 880 50792 399200 51072
rect 800 50120 399200 50792
rect 800 49840 399120 50120
rect 800 49168 399200 49840
rect 880 48888 399200 49168
rect 800 48760 399200 48888
rect 800 48480 399120 48760
rect 800 47400 399200 48480
rect 800 47264 399120 47400
rect 880 47120 399120 47264
rect 880 46984 399200 47120
rect 800 46040 399200 46984
rect 800 45760 399120 46040
rect 800 45224 399200 45760
rect 880 44944 399200 45224
rect 800 44680 399200 44944
rect 800 44400 399120 44680
rect 800 43320 399200 44400
rect 880 43040 399120 43320
rect 800 41960 399200 43040
rect 800 41680 399120 41960
rect 800 41416 399200 41680
rect 880 41136 399200 41416
rect 800 40600 399200 41136
rect 800 40320 399120 40600
rect 800 39512 399200 40320
rect 880 39240 399200 39512
rect 880 39232 399120 39240
rect 800 38960 399120 39232
rect 800 37880 399200 38960
rect 800 37608 399120 37880
rect 880 37600 399120 37608
rect 880 37328 399200 37600
rect 800 36384 399200 37328
rect 800 36104 399120 36384
rect 800 35704 399200 36104
rect 880 35424 399200 35704
rect 800 35024 399200 35424
rect 800 34744 399120 35024
rect 800 33800 399200 34744
rect 880 33664 399200 33800
rect 880 33520 399120 33664
rect 800 33384 399120 33520
rect 800 32304 399200 33384
rect 800 32024 399120 32304
rect 800 31896 399200 32024
rect 880 31616 399200 31896
rect 800 30944 399200 31616
rect 800 30664 399120 30944
rect 800 29856 399200 30664
rect 880 29584 399200 29856
rect 880 29576 399120 29584
rect 800 29304 399120 29576
rect 800 28224 399200 29304
rect 800 27952 399120 28224
rect 880 27944 399120 27952
rect 880 27672 399200 27944
rect 800 26864 399200 27672
rect 800 26584 399120 26864
rect 800 26048 399200 26584
rect 880 25768 399200 26048
rect 800 25504 399200 25768
rect 800 25224 399120 25504
rect 800 24144 399200 25224
rect 880 23864 399120 24144
rect 800 22784 399200 23864
rect 800 22504 399120 22784
rect 800 22240 399200 22504
rect 880 21960 399200 22240
rect 800 21424 399200 21960
rect 800 21144 399120 21424
rect 800 20336 399200 21144
rect 880 20064 399200 20336
rect 880 20056 399120 20064
rect 800 19784 399120 20056
rect 800 18568 399200 19784
rect 800 18432 399120 18568
rect 880 18288 399120 18432
rect 880 18152 399200 18288
rect 800 17208 399200 18152
rect 800 16928 399120 17208
rect 800 16528 399200 16928
rect 880 16248 399200 16528
rect 800 15848 399200 16248
rect 800 15568 399120 15848
rect 800 14488 399200 15568
rect 880 14208 399120 14488
rect 800 13128 399200 14208
rect 800 12848 399120 13128
rect 800 12584 399200 12848
rect 880 12304 399200 12584
rect 800 11768 399200 12304
rect 800 11488 399120 11768
rect 800 10680 399200 11488
rect 880 10408 399200 10680
rect 880 10400 399120 10408
rect 800 10128 399120 10400
rect 800 9048 399200 10128
rect 800 8776 399120 9048
rect 880 8768 399120 8776
rect 880 8496 399200 8768
rect 800 7688 399200 8496
rect 800 7408 399120 7688
rect 800 6872 399200 7408
rect 880 6592 399200 6872
rect 800 6328 399200 6592
rect 800 6048 399120 6328
rect 800 4968 399200 6048
rect 880 4688 399120 4968
rect 800 3608 399200 4688
rect 800 3328 399120 3608
rect 800 3064 399200 3328
rect 880 2784 399200 3064
rect 800 2248 399200 2784
rect 800 1968 399120 2248
rect 800 1160 399200 1968
rect 880 888 399200 1160
rect 880 880 399120 888
rect 800 715 399120 880
<< metal4 >>
rect 4 156 324 147812
rect 664 816 984 147152
rect 5128 156 5448 147812
rect 10128 156 10448 147812
rect 15128 156 15448 147812
rect 20128 107460 20448 147812
rect 25128 107460 25448 147812
rect 30128 107460 30448 147812
rect 35128 107460 35448 147812
rect 40128 107460 40448 147812
rect 45128 107460 45448 147812
rect 50128 107460 50448 147812
rect 55128 107460 55448 147812
rect 60128 107460 60448 147812
rect 65128 107460 65448 147812
rect 70128 107460 70448 147812
rect 75128 107460 75448 147812
rect 80128 107460 80448 147812
rect 85128 107460 85448 147812
rect 90128 107460 90448 147812
rect 95128 107460 95448 147812
rect 100128 107460 100448 147812
rect 105128 107460 105448 147812
rect 110128 107460 110448 147812
rect 115128 107460 115448 147812
rect 120128 107460 120448 147812
rect 125128 107460 125448 147812
rect 130128 107460 130448 147812
rect 135128 107460 135448 147812
rect 140128 107460 140448 147812
rect 145128 107460 145448 147812
rect 150128 107460 150448 147812
rect 155128 107460 155448 147812
rect 20128 156 20448 20248
rect 25128 156 25448 20248
rect 30128 156 30448 20248
rect 35128 156 35448 20248
rect 40128 156 40448 20248
rect 45128 156 45448 20248
rect 50128 156 50448 20248
rect 55128 156 55448 20248
rect 60128 156 60448 20248
rect 65128 156 65448 20248
rect 70128 156 70448 20248
rect 75128 156 75448 20248
rect 80128 156 80448 20248
rect 85128 156 85448 20248
rect 90128 156 90448 20248
rect 95128 156 95448 20248
rect 100128 156 100448 20248
rect 105128 156 105448 20248
rect 110128 156 110448 20248
rect 115128 156 115448 20248
rect 120128 156 120448 20248
rect 125128 156 125448 20248
rect 130128 156 130448 20248
rect 135128 156 135448 20248
rect 140128 156 140448 20248
rect 145128 156 145448 20248
rect 150128 156 150448 20248
rect 155128 156 155448 20248
rect 160128 156 160448 147812
rect 165128 156 165448 147812
rect 170128 156 170448 147812
rect 175128 156 175448 147812
rect 180128 156 180448 147812
rect 185128 156 185448 147812
rect 190128 156 190448 147812
rect 195128 156 195448 147812
rect 200128 156 200448 147812
rect 205128 156 205448 147812
rect 210128 156 210448 147812
rect 215128 156 215448 147812
rect 220128 156 220448 147812
rect 225128 156 225448 147812
rect 230128 156 230448 147812
rect 235128 156 235448 147812
rect 240128 156 240448 147812
rect 245128 156 245448 147812
rect 250128 156 250448 147812
rect 255128 156 255448 147812
rect 260128 156 260448 147812
rect 265128 156 265448 147812
rect 270128 156 270448 147812
rect 275128 156 275448 147812
rect 280128 156 280448 147812
rect 285128 156 285448 147812
rect 290128 156 290448 147812
rect 295128 156 295448 147812
rect 300128 156 300448 147812
rect 305128 156 305448 147812
rect 310128 156 310448 147812
rect 315128 156 315448 147812
rect 320128 156 320448 147812
rect 325128 156 325448 147812
rect 330128 156 330448 147812
rect 335128 156 335448 147812
rect 340128 156 340448 147812
rect 345128 156 345448 147812
rect 350128 156 350448 147812
rect 355128 156 355448 147812
rect 360128 156 360448 147812
rect 365128 156 365448 147812
rect 370128 156 370448 147812
rect 375128 156 375448 147812
rect 380128 156 380448 147812
rect 385128 156 385448 147812
rect 390128 156 390448 147812
rect 395128 156 395448 147812
rect 398940 816 399260 147152
rect 399600 156 399920 147812
<< obsm4 >>
rect 4291 9555 5048 147253
rect 5528 9555 10048 147253
rect 10528 9555 15048 147253
rect 15528 107380 20048 147253
rect 20528 107380 25048 147253
rect 25528 107380 30048 147253
rect 30528 107380 35048 147253
rect 35528 107380 40048 147253
rect 40528 107380 45048 147253
rect 45528 107380 50048 147253
rect 50528 107380 55048 147253
rect 55528 107380 60048 147253
rect 60528 107380 65048 147253
rect 65528 107380 70048 147253
rect 70528 107380 75048 147253
rect 75528 107380 80048 147253
rect 80528 107380 85048 147253
rect 85528 107380 90048 147253
rect 90528 107380 95048 147253
rect 95528 107380 100048 147253
rect 100528 107380 105048 147253
rect 105528 107380 110048 147253
rect 110528 107380 115048 147253
rect 115528 107380 120048 147253
rect 120528 107380 125048 147253
rect 125528 107380 130048 147253
rect 130528 107380 135048 147253
rect 135528 107380 140048 147253
rect 140528 107380 145048 147253
rect 145528 107380 150048 147253
rect 150528 107380 155048 147253
rect 155528 107380 160048 147253
rect 15528 20328 160048 107380
rect 15528 9555 20048 20328
rect 20528 9555 25048 20328
rect 25528 9555 30048 20328
rect 30528 9555 35048 20328
rect 35528 9555 40048 20328
rect 40528 9555 45048 20328
rect 45528 9555 50048 20328
rect 50528 9555 55048 20328
rect 55528 9555 60048 20328
rect 60528 9555 65048 20328
rect 65528 9555 70048 20328
rect 70528 9555 75048 20328
rect 75528 9555 80048 20328
rect 80528 9555 85048 20328
rect 85528 9555 90048 20328
rect 90528 9555 95048 20328
rect 95528 9555 100048 20328
rect 100528 9555 105048 20328
rect 105528 9555 110048 20328
rect 110528 9555 115048 20328
rect 115528 9555 120048 20328
rect 120528 9555 125048 20328
rect 125528 9555 130048 20328
rect 130528 9555 135048 20328
rect 135528 9555 140048 20328
rect 140528 9555 145048 20328
rect 145528 9555 150048 20328
rect 150528 9555 155048 20328
rect 155528 9555 160048 20328
rect 160528 9555 165048 147253
rect 165528 9555 170048 147253
rect 170528 9555 175048 147253
rect 175528 9555 180048 147253
rect 180528 9555 185048 147253
rect 185528 9555 190048 147253
rect 190528 9555 195048 147253
rect 195528 9555 200048 147253
rect 200528 9555 205048 147253
rect 205528 9555 210048 147253
rect 210528 9555 215048 147253
rect 215528 9555 220048 147253
rect 220528 9555 225048 147253
rect 225528 9555 230048 147253
rect 230528 9555 235048 147253
rect 235528 9555 240048 147253
rect 240528 9555 245048 147253
rect 245528 9555 250048 147253
rect 250528 9555 255048 147253
rect 255528 9555 260048 147253
rect 260528 9555 265048 147253
rect 265528 9555 270048 147253
rect 270528 9555 275048 147253
rect 275528 9555 280048 147253
rect 280528 9555 285048 147253
rect 285528 9555 290048 147253
rect 290528 9555 295048 147253
rect 295528 9555 300048 147253
rect 300528 9555 305048 147253
rect 305528 9555 310048 147253
rect 310528 9555 315048 147253
rect 315528 9555 320048 147253
rect 320528 9555 325048 147253
rect 325528 9555 330048 147253
rect 330528 9555 335048 147253
rect 335528 9555 340048 147253
rect 340528 9555 345048 147253
rect 345528 9555 350048 147253
rect 350528 9555 355048 147253
rect 355528 9555 360048 147253
rect 360528 9555 365048 147253
rect 365528 9555 370048 147253
rect 370528 9555 375048 147253
rect 375528 9555 376589 147253
<< metal5 >>
rect 4 147492 399920 147812
rect 664 146832 399260 147152
rect 4 135298 399920 135618
rect 4 122298 399920 122618
rect 4 109298 399920 109618
rect 4 96298 399920 96618
rect 4 83298 399920 83618
rect 4 70298 399920 70618
rect 4 57298 399920 57618
rect 4 44298 399920 44618
rect 4 31298 399920 31618
rect 4 18298 399920 18618
rect 4 5298 399920 5618
rect 664 816 399260 1136
rect 4 156 399920 476
<< obsm5 >>
rect 6188 135938 314892 146020
rect 6188 122938 314892 134978
rect 6188 109938 314892 121978
rect 6188 96938 314892 108978
rect 6188 83938 314892 95978
rect 6188 70938 314892 82978
rect 6188 57938 314892 69978
rect 6188 44938 314892 56978
rect 6188 31938 314892 43978
rect 6188 18938 314892 30978
rect 6188 17180 314892 17978
<< labels >>
rlabel metal5 s 4 156 399920 476 6 VGND
port 1 nsew ground input
rlabel metal5 s 4 18298 399920 18618 6 VGND
port 1 nsew ground input
rlabel metal5 s 4 44298 399920 44618 6 VGND
port 1 nsew ground input
rlabel metal5 s 4 70298 399920 70618 6 VGND
port 1 nsew ground input
rlabel metal5 s 4 96298 399920 96618 6 VGND
port 1 nsew ground input
rlabel metal5 s 4 122298 399920 122618 6 VGND
port 1 nsew ground input
rlabel metal5 s 4 147492 399920 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 20128 156 20448 20248 6 VGND
port 1 nsew ground input
rlabel metal4 s 30128 156 30448 20248 6 VGND
port 1 nsew ground input
rlabel metal4 s 40128 156 40448 20248 6 VGND
port 1 nsew ground input
rlabel metal4 s 50128 156 50448 20248 6 VGND
port 1 nsew ground input
rlabel metal4 s 60128 156 60448 20248 6 VGND
port 1 nsew ground input
rlabel metal4 s 70128 156 70448 20248 6 VGND
port 1 nsew ground input
rlabel metal4 s 80128 156 80448 20248 6 VGND
port 1 nsew ground input
rlabel metal4 s 90128 156 90448 20248 6 VGND
port 1 nsew ground input
rlabel metal4 s 100128 156 100448 20248 6 VGND
port 1 nsew ground input
rlabel metal4 s 110128 156 110448 20248 6 VGND
port 1 nsew ground input
rlabel metal4 s 120128 156 120448 20248 6 VGND
port 1 nsew ground input
rlabel metal4 s 130128 156 130448 20248 6 VGND
port 1 nsew ground input
rlabel metal4 s 140128 156 140448 20248 6 VGND
port 1 nsew ground input
rlabel metal4 s 150128 156 150448 20248 6 VGND
port 1 nsew ground input
rlabel metal4 s 4 156 324 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 10128 156 10448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 20128 107460 20448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 30128 107460 30448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 40128 107460 40448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 50128 107460 50448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 60128 107460 60448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 70128 107460 70448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 80128 107460 80448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 90128 107460 90448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 100128 107460 100448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 110128 107460 110448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 120128 107460 120448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 130128 107460 130448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 140128 107460 140448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 150128 107460 150448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 160128 156 160448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 170128 156 170448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 180128 156 180448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 190128 156 190448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 200128 156 200448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 210128 156 210448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 220128 156 220448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 230128 156 230448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 240128 156 240448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 250128 156 250448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 260128 156 260448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 270128 156 270448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 280128 156 280448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 290128 156 290448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 300128 156 300448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 310128 156 310448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 320128 156 320448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 330128 156 330448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 340128 156 340448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 350128 156 350448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 360128 156 360448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 370128 156 370448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 380128 156 380448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 390128 156 390448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 399600 156 399920 147812 6 VGND
port 1 nsew ground input
rlabel metal5 s 664 816 399260 1136 6 VPWR
port 2 nsew power input
rlabel metal5 s 4 5298 399920 5618 6 VPWR
port 2 nsew power input
rlabel metal5 s 4 31298 399920 31618 6 VPWR
port 2 nsew power input
rlabel metal5 s 4 57298 399920 57618 6 VPWR
port 2 nsew power input
rlabel metal5 s 4 83298 399920 83618 6 VPWR
port 2 nsew power input
rlabel metal5 s 4 109298 399920 109618 6 VPWR
port 2 nsew power input
rlabel metal5 s 4 135298 399920 135618 6 VPWR
port 2 nsew power input
rlabel metal5 s 664 146832 399260 147152 6 VPWR
port 2 nsew power input
rlabel metal4 s 25128 156 25448 20248 6 VPWR
port 2 nsew power input
rlabel metal4 s 35128 156 35448 20248 6 VPWR
port 2 nsew power input
rlabel metal4 s 45128 156 45448 20248 6 VPWR
port 2 nsew power input
rlabel metal4 s 55128 156 55448 20248 6 VPWR
port 2 nsew power input
rlabel metal4 s 65128 156 65448 20248 6 VPWR
port 2 nsew power input
rlabel metal4 s 75128 156 75448 20248 6 VPWR
port 2 nsew power input
rlabel metal4 s 85128 156 85448 20248 6 VPWR
port 2 nsew power input
rlabel metal4 s 95128 156 95448 20248 6 VPWR
port 2 nsew power input
rlabel metal4 s 105128 156 105448 20248 6 VPWR
port 2 nsew power input
rlabel metal4 s 115128 156 115448 20248 6 VPWR
port 2 nsew power input
rlabel metal4 s 125128 156 125448 20248 6 VPWR
port 2 nsew power input
rlabel metal4 s 135128 156 135448 20248 6 VPWR
port 2 nsew power input
rlabel metal4 s 145128 156 145448 20248 6 VPWR
port 2 nsew power input
rlabel metal4 s 155128 156 155448 20248 6 VPWR
port 2 nsew power input
rlabel metal4 s 664 816 984 147152 6 VPWR
port 2 nsew power input
rlabel metal4 s 398940 816 399260 147152 6 VPWR
port 2 nsew power input
rlabel metal4 s 5128 156 5448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 15128 156 15448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 25128 107460 25448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 35128 107460 35448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 45128 107460 45448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 55128 107460 55448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 65128 107460 65448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 75128 107460 75448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 85128 107460 85448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 95128 107460 95448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 105128 107460 105448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 115128 107460 115448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 125128 107460 125448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 135128 107460 135448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 145128 107460 145448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 155128 107460 155448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 165128 156 165448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 175128 156 175448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 185128 156 185448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 195128 156 195448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 205128 156 205448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 215128 156 215448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 225128 156 225448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 235128 156 235448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 245128 156 245448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 255128 156 255448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 265128 156 265448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 275128 156 275448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 285128 156 285448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 295128 156 295448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 305128 156 305448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 315128 156 315448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 325128 156 325448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 335128 156 335448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 345128 156 345448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 355128 156 355448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 365128 156 365448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 375128 156 375448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 385128 156 385448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 395128 156 395448 147812 6 VPWR
port 2 nsew power input
rlabel metal2 s 224958 0 225014 800 6 clk
port 3 nsew signal input
rlabel metal3 s 399200 58216 400000 58336 6 debug_in
port 4 nsew signal input
rlabel metal3 s 399200 59576 400000 59696 6 debug_mode
port 5 nsew signal output
rlabel metal3 s 399200 60936 400000 61056 6 debug_oeb
port 6 nsew signal output
rlabel metal3 s 399200 62296 400000 62416 6 debug_out
port 7 nsew signal output
rlabel metal3 s 399200 130840 400000 130960 6 flash_clk
port 8 nsew signal output
rlabel metal3 s 399200 129344 400000 129464 6 flash_csb
port 9 nsew signal output
rlabel metal3 s 399200 132200 400000 132320 6 flash_io0_di
port 10 nsew signal input
rlabel metal3 s 399200 133560 400000 133680 6 flash_io0_do
port 11 nsew signal output
rlabel metal3 s 399200 134920 400000 135040 6 flash_io0_oeb
port 12 nsew signal output
rlabel metal3 s 399200 136280 400000 136400 6 flash_io1_di
port 13 nsew signal input
rlabel metal3 s 399200 137640 400000 137760 6 flash_io1_do
port 14 nsew signal output
rlabel metal3 s 399200 139000 400000 139120 6 flash_io1_oeb
port 15 nsew signal output
rlabel metal3 s 399200 140360 400000 140480 6 flash_io2_di
port 16 nsew signal input
rlabel metal3 s 399200 141720 400000 141840 6 flash_io2_do
port 17 nsew signal output
rlabel metal3 s 399200 143080 400000 143200 6 flash_io2_oeb
port 18 nsew signal output
rlabel metal3 s 399200 144440 400000 144560 6 flash_io3_di
port 19 nsew signal input
rlabel metal3 s 399200 145800 400000 145920 6 flash_io3_do
port 20 nsew signal output
rlabel metal3 s 399200 147160 400000 147280 6 flash_io3_oeb
port 21 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 gpio_in_pad
port 22 nsew signal input
rlabel metal2 s 124954 0 125010 800 6 gpio_inenb_pad
port 23 nsew signal output
rlabel metal2 s 174910 0 174966 800 6 gpio_mode0_pad
port 24 nsew signal output
rlabel metal2 s 274914 0 274970 800 6 gpio_mode1_pad
port 25 nsew signal output
rlabel metal2 s 324962 0 325018 800 6 gpio_out_pad
port 26 nsew signal output
rlabel metal2 s 374918 0 374974 800 6 gpio_outenb_pad
port 27 nsew signal output
rlabel metal3 s 399200 82832 400000 82952 6 hk_ack_i
port 28 nsew signal input
rlabel metal3 s 399200 85552 400000 85672 6 hk_dat_i[0]
port 29 nsew signal input
rlabel metal3 s 399200 99288 400000 99408 6 hk_dat_i[10]
port 30 nsew signal input
rlabel metal3 s 399200 100648 400000 100768 6 hk_dat_i[11]
port 31 nsew signal input
rlabel metal3 s 399200 102008 400000 102128 6 hk_dat_i[12]
port 32 nsew signal input
rlabel metal3 s 399200 103368 400000 103488 6 hk_dat_i[13]
port 33 nsew signal input
rlabel metal3 s 399200 104728 400000 104848 6 hk_dat_i[14]
port 34 nsew signal input
rlabel metal3 s 399200 106088 400000 106208 6 hk_dat_i[15]
port 35 nsew signal input
rlabel metal3 s 399200 107448 400000 107568 6 hk_dat_i[16]
port 36 nsew signal input
rlabel metal3 s 399200 108808 400000 108928 6 hk_dat_i[17]
port 37 nsew signal input
rlabel metal3 s 399200 110168 400000 110288 6 hk_dat_i[18]
port 38 nsew signal input
rlabel metal3 s 399200 111664 400000 111784 6 hk_dat_i[19]
port 39 nsew signal input
rlabel metal3 s 399200 86912 400000 87032 6 hk_dat_i[1]
port 40 nsew signal input
rlabel metal3 s 399200 113024 400000 113144 6 hk_dat_i[20]
port 41 nsew signal input
rlabel metal3 s 399200 114384 400000 114504 6 hk_dat_i[21]
port 42 nsew signal input
rlabel metal3 s 399200 115744 400000 115864 6 hk_dat_i[22]
port 43 nsew signal input
rlabel metal3 s 399200 117104 400000 117224 6 hk_dat_i[23]
port 44 nsew signal input
rlabel metal3 s 399200 118464 400000 118584 6 hk_dat_i[24]
port 45 nsew signal input
rlabel metal3 s 399200 119824 400000 119944 6 hk_dat_i[25]
port 46 nsew signal input
rlabel metal3 s 399200 121184 400000 121304 6 hk_dat_i[26]
port 47 nsew signal input
rlabel metal3 s 399200 122544 400000 122664 6 hk_dat_i[27]
port 48 nsew signal input
rlabel metal3 s 399200 123904 400000 124024 6 hk_dat_i[28]
port 49 nsew signal input
rlabel metal3 s 399200 125264 400000 125384 6 hk_dat_i[29]
port 50 nsew signal input
rlabel metal3 s 399200 88272 400000 88392 6 hk_dat_i[2]
port 51 nsew signal input
rlabel metal3 s 399200 126624 400000 126744 6 hk_dat_i[30]
port 52 nsew signal input
rlabel metal3 s 399200 127984 400000 128104 6 hk_dat_i[31]
port 53 nsew signal input
rlabel metal3 s 399200 89632 400000 89752 6 hk_dat_i[3]
port 54 nsew signal input
rlabel metal3 s 399200 90992 400000 91112 6 hk_dat_i[4]
port 55 nsew signal input
rlabel metal3 s 399200 92352 400000 92472 6 hk_dat_i[5]
port 56 nsew signal input
rlabel metal3 s 399200 93848 400000 93968 6 hk_dat_i[6]
port 57 nsew signal input
rlabel metal3 s 399200 95208 400000 95328 6 hk_dat_i[7]
port 58 nsew signal input
rlabel metal3 s 399200 96568 400000 96688 6 hk_dat_i[8]
port 59 nsew signal input
rlabel metal3 s 399200 97928 400000 98048 6 hk_dat_i[9]
port 60 nsew signal input
rlabel metal3 s 399200 84192 400000 84312 6 hk_stb_o
port 61 nsew signal output
rlabel metal2 s 398378 147200 398434 148000 6 irq[0]
port 62 nsew signal input
rlabel metal2 s 399022 147200 399078 148000 6 irq[1]
port 63 nsew signal input
rlabel metal2 s 399666 147200 399722 148000 6 irq[2]
port 64 nsew signal input
rlabel metal3 s 399200 67736 400000 67856 6 irq[3]
port 65 nsew signal input
rlabel metal3 s 399200 66376 400000 66496 6 irq[4]
port 66 nsew signal input
rlabel metal3 s 399200 65016 400000 65136 6 irq[5]
port 67 nsew signal input
rlabel metal2 s 294 147200 350 148000 6 la_iena[0]
port 68 nsew signal output
rlabel metal2 s 257066 147200 257122 148000 6 la_iena[100]
port 69 nsew signal output
rlabel metal2 s 259642 147200 259698 148000 6 la_iena[101]
port 70 nsew signal output
rlabel metal2 s 262218 147200 262274 148000 6 la_iena[102]
port 71 nsew signal output
rlabel metal2 s 264794 147200 264850 148000 6 la_iena[103]
port 72 nsew signal output
rlabel metal2 s 267370 147200 267426 148000 6 la_iena[104]
port 73 nsew signal output
rlabel metal2 s 269946 147200 270002 148000 6 la_iena[105]
port 74 nsew signal output
rlabel metal2 s 272522 147200 272578 148000 6 la_iena[106]
port 75 nsew signal output
rlabel metal2 s 275098 147200 275154 148000 6 la_iena[107]
port 76 nsew signal output
rlabel metal2 s 277582 147200 277638 148000 6 la_iena[108]
port 77 nsew signal output
rlabel metal2 s 280158 147200 280214 148000 6 la_iena[109]
port 78 nsew signal output
rlabel metal2 s 25962 147200 26018 148000 6 la_iena[10]
port 79 nsew signal output
rlabel metal2 s 282734 147200 282790 148000 6 la_iena[110]
port 80 nsew signal output
rlabel metal2 s 285310 147200 285366 148000 6 la_iena[111]
port 81 nsew signal output
rlabel metal2 s 287886 147200 287942 148000 6 la_iena[112]
port 82 nsew signal output
rlabel metal2 s 290462 147200 290518 148000 6 la_iena[113]
port 83 nsew signal output
rlabel metal2 s 293038 147200 293094 148000 6 la_iena[114]
port 84 nsew signal output
rlabel metal2 s 295614 147200 295670 148000 6 la_iena[115]
port 85 nsew signal output
rlabel metal2 s 298190 147200 298246 148000 6 la_iena[116]
port 86 nsew signal output
rlabel metal2 s 300766 147200 300822 148000 6 la_iena[117]
port 87 nsew signal output
rlabel metal2 s 303342 147200 303398 148000 6 la_iena[118]
port 88 nsew signal output
rlabel metal2 s 305918 147200 305974 148000 6 la_iena[119]
port 89 nsew signal output
rlabel metal2 s 28538 147200 28594 148000 6 la_iena[11]
port 90 nsew signal output
rlabel metal2 s 308402 147200 308458 148000 6 la_iena[120]
port 91 nsew signal output
rlabel metal2 s 310978 147200 311034 148000 6 la_iena[121]
port 92 nsew signal output
rlabel metal2 s 313554 147200 313610 148000 6 la_iena[122]
port 93 nsew signal output
rlabel metal2 s 316130 147200 316186 148000 6 la_iena[123]
port 94 nsew signal output
rlabel metal2 s 318706 147200 318762 148000 6 la_iena[124]
port 95 nsew signal output
rlabel metal2 s 321282 147200 321338 148000 6 la_iena[125]
port 96 nsew signal output
rlabel metal2 s 323858 147200 323914 148000 6 la_iena[126]
port 97 nsew signal output
rlabel metal2 s 326434 147200 326490 148000 6 la_iena[127]
port 98 nsew signal output
rlabel metal2 s 31022 147200 31078 148000 6 la_iena[12]
port 99 nsew signal output
rlabel metal2 s 33598 147200 33654 148000 6 la_iena[13]
port 100 nsew signal output
rlabel metal2 s 36174 147200 36230 148000 6 la_iena[14]
port 101 nsew signal output
rlabel metal2 s 38750 147200 38806 148000 6 la_iena[15]
port 102 nsew signal output
rlabel metal2 s 41326 147200 41382 148000 6 la_iena[16]
port 103 nsew signal output
rlabel metal2 s 43902 147200 43958 148000 6 la_iena[17]
port 104 nsew signal output
rlabel metal2 s 46478 147200 46534 148000 6 la_iena[18]
port 105 nsew signal output
rlabel metal2 s 49054 147200 49110 148000 6 la_iena[19]
port 106 nsew signal output
rlabel metal2 s 2778 147200 2834 148000 6 la_iena[1]
port 107 nsew signal output
rlabel metal2 s 51630 147200 51686 148000 6 la_iena[20]
port 108 nsew signal output
rlabel metal2 s 54206 147200 54262 148000 6 la_iena[21]
port 109 nsew signal output
rlabel metal2 s 56782 147200 56838 148000 6 la_iena[22]
port 110 nsew signal output
rlabel metal2 s 59358 147200 59414 148000 6 la_iena[23]
port 111 nsew signal output
rlabel metal2 s 61842 147200 61898 148000 6 la_iena[24]
port 112 nsew signal output
rlabel metal2 s 64418 147200 64474 148000 6 la_iena[25]
port 113 nsew signal output
rlabel metal2 s 66994 147200 67050 148000 6 la_iena[26]
port 114 nsew signal output
rlabel metal2 s 69570 147200 69626 148000 6 la_iena[27]
port 115 nsew signal output
rlabel metal2 s 72146 147200 72202 148000 6 la_iena[28]
port 116 nsew signal output
rlabel metal2 s 74722 147200 74778 148000 6 la_iena[29]
port 117 nsew signal output
rlabel metal2 s 5354 147200 5410 148000 6 la_iena[2]
port 118 nsew signal output
rlabel metal2 s 77298 147200 77354 148000 6 la_iena[30]
port 119 nsew signal output
rlabel metal2 s 79874 147200 79930 148000 6 la_iena[31]
port 120 nsew signal output
rlabel metal2 s 82450 147200 82506 148000 6 la_iena[32]
port 121 nsew signal output
rlabel metal2 s 85026 147200 85082 148000 6 la_iena[33]
port 122 nsew signal output
rlabel metal2 s 87602 147200 87658 148000 6 la_iena[34]
port 123 nsew signal output
rlabel metal2 s 90178 147200 90234 148000 6 la_iena[35]
port 124 nsew signal output
rlabel metal2 s 92662 147200 92718 148000 6 la_iena[36]
port 125 nsew signal output
rlabel metal2 s 95238 147200 95294 148000 6 la_iena[37]
port 126 nsew signal output
rlabel metal2 s 97814 147200 97870 148000 6 la_iena[38]
port 127 nsew signal output
rlabel metal2 s 100390 147200 100446 148000 6 la_iena[39]
port 128 nsew signal output
rlabel metal2 s 7930 147200 7986 148000 6 la_iena[3]
port 129 nsew signal output
rlabel metal2 s 102966 147200 103022 148000 6 la_iena[40]
port 130 nsew signal output
rlabel metal2 s 105542 147200 105598 148000 6 la_iena[41]
port 131 nsew signal output
rlabel metal2 s 108118 147200 108174 148000 6 la_iena[42]
port 132 nsew signal output
rlabel metal2 s 110694 147200 110750 148000 6 la_iena[43]
port 133 nsew signal output
rlabel metal2 s 113270 147200 113326 148000 6 la_iena[44]
port 134 nsew signal output
rlabel metal2 s 115846 147200 115902 148000 6 la_iena[45]
port 135 nsew signal output
rlabel metal2 s 118422 147200 118478 148000 6 la_iena[46]
port 136 nsew signal output
rlabel metal2 s 120998 147200 121054 148000 6 la_iena[47]
port 137 nsew signal output
rlabel metal2 s 123482 147200 123538 148000 6 la_iena[48]
port 138 nsew signal output
rlabel metal2 s 126058 147200 126114 148000 6 la_iena[49]
port 139 nsew signal output
rlabel metal2 s 10506 147200 10562 148000 6 la_iena[4]
port 140 nsew signal output
rlabel metal2 s 128634 147200 128690 148000 6 la_iena[50]
port 141 nsew signal output
rlabel metal2 s 131210 147200 131266 148000 6 la_iena[51]
port 142 nsew signal output
rlabel metal2 s 133786 147200 133842 148000 6 la_iena[52]
port 143 nsew signal output
rlabel metal2 s 136362 147200 136418 148000 6 la_iena[53]
port 144 nsew signal output
rlabel metal2 s 138938 147200 138994 148000 6 la_iena[54]
port 145 nsew signal output
rlabel metal2 s 141514 147200 141570 148000 6 la_iena[55]
port 146 nsew signal output
rlabel metal2 s 144090 147200 144146 148000 6 la_iena[56]
port 147 nsew signal output
rlabel metal2 s 146666 147200 146722 148000 6 la_iena[57]
port 148 nsew signal output
rlabel metal2 s 149242 147200 149298 148000 6 la_iena[58]
port 149 nsew signal output
rlabel metal2 s 151818 147200 151874 148000 6 la_iena[59]
port 150 nsew signal output
rlabel metal2 s 13082 147200 13138 148000 6 la_iena[5]
port 151 nsew signal output
rlabel metal2 s 154302 147200 154358 148000 6 la_iena[60]
port 152 nsew signal output
rlabel metal2 s 156878 147200 156934 148000 6 la_iena[61]
port 153 nsew signal output
rlabel metal2 s 159454 147200 159510 148000 6 la_iena[62]
port 154 nsew signal output
rlabel metal2 s 162030 147200 162086 148000 6 la_iena[63]
port 155 nsew signal output
rlabel metal2 s 164606 147200 164662 148000 6 la_iena[64]
port 156 nsew signal output
rlabel metal2 s 167182 147200 167238 148000 6 la_iena[65]
port 157 nsew signal output
rlabel metal2 s 169758 147200 169814 148000 6 la_iena[66]
port 158 nsew signal output
rlabel metal2 s 172334 147200 172390 148000 6 la_iena[67]
port 159 nsew signal output
rlabel metal2 s 174910 147200 174966 148000 6 la_iena[68]
port 160 nsew signal output
rlabel metal2 s 177486 147200 177542 148000 6 la_iena[69]
port 161 nsew signal output
rlabel metal2 s 15658 147200 15714 148000 6 la_iena[6]
port 162 nsew signal output
rlabel metal2 s 180062 147200 180118 148000 6 la_iena[70]
port 163 nsew signal output
rlabel metal2 s 182638 147200 182694 148000 6 la_iena[71]
port 164 nsew signal output
rlabel metal2 s 185122 147200 185178 148000 6 la_iena[72]
port 165 nsew signal output
rlabel metal2 s 187698 147200 187754 148000 6 la_iena[73]
port 166 nsew signal output
rlabel metal2 s 190274 147200 190330 148000 6 la_iena[74]
port 167 nsew signal output
rlabel metal2 s 192850 147200 192906 148000 6 la_iena[75]
port 168 nsew signal output
rlabel metal2 s 195426 147200 195482 148000 6 la_iena[76]
port 169 nsew signal output
rlabel metal2 s 198002 147200 198058 148000 6 la_iena[77]
port 170 nsew signal output
rlabel metal2 s 200578 147200 200634 148000 6 la_iena[78]
port 171 nsew signal output
rlabel metal2 s 203154 147200 203210 148000 6 la_iena[79]
port 172 nsew signal output
rlabel metal2 s 18234 147200 18290 148000 6 la_iena[7]
port 173 nsew signal output
rlabel metal2 s 205730 147200 205786 148000 6 la_iena[80]
port 174 nsew signal output
rlabel metal2 s 208306 147200 208362 148000 6 la_iena[81]
port 175 nsew signal output
rlabel metal2 s 210882 147200 210938 148000 6 la_iena[82]
port 176 nsew signal output
rlabel metal2 s 213458 147200 213514 148000 6 la_iena[83]
port 177 nsew signal output
rlabel metal2 s 215942 147200 215998 148000 6 la_iena[84]
port 178 nsew signal output
rlabel metal2 s 218518 147200 218574 148000 6 la_iena[85]
port 179 nsew signal output
rlabel metal2 s 221094 147200 221150 148000 6 la_iena[86]
port 180 nsew signal output
rlabel metal2 s 223670 147200 223726 148000 6 la_iena[87]
port 181 nsew signal output
rlabel metal2 s 226246 147200 226302 148000 6 la_iena[88]
port 182 nsew signal output
rlabel metal2 s 228822 147200 228878 148000 6 la_iena[89]
port 183 nsew signal output
rlabel metal2 s 20810 147200 20866 148000 6 la_iena[8]
port 184 nsew signal output
rlabel metal2 s 231398 147200 231454 148000 6 la_iena[90]
port 185 nsew signal output
rlabel metal2 s 233974 147200 234030 148000 6 la_iena[91]
port 186 nsew signal output
rlabel metal2 s 236550 147200 236606 148000 6 la_iena[92]
port 187 nsew signal output
rlabel metal2 s 239126 147200 239182 148000 6 la_iena[93]
port 188 nsew signal output
rlabel metal2 s 241702 147200 241758 148000 6 la_iena[94]
port 189 nsew signal output
rlabel metal2 s 244278 147200 244334 148000 6 la_iena[95]
port 190 nsew signal output
rlabel metal2 s 246762 147200 246818 148000 6 la_iena[96]
port 191 nsew signal output
rlabel metal2 s 249338 147200 249394 148000 6 la_iena[97]
port 192 nsew signal output
rlabel metal2 s 251914 147200 251970 148000 6 la_iena[98]
port 193 nsew signal output
rlabel metal2 s 254490 147200 254546 148000 6 la_iena[99]
port 194 nsew signal output
rlabel metal2 s 23386 147200 23442 148000 6 la_iena[9]
port 195 nsew signal output
rlabel metal2 s 846 147200 902 148000 6 la_input[0]
port 196 nsew signal input
rlabel metal2 s 257710 147200 257766 148000 6 la_input[100]
port 197 nsew signal input
rlabel metal2 s 260286 147200 260342 148000 6 la_input[101]
port 198 nsew signal input
rlabel metal2 s 262862 147200 262918 148000 6 la_input[102]
port 199 nsew signal input
rlabel metal2 s 265438 147200 265494 148000 6 la_input[103]
port 200 nsew signal input
rlabel metal2 s 268014 147200 268070 148000 6 la_input[104]
port 201 nsew signal input
rlabel metal2 s 270590 147200 270646 148000 6 la_input[105]
port 202 nsew signal input
rlabel metal2 s 273166 147200 273222 148000 6 la_input[106]
port 203 nsew signal input
rlabel metal2 s 275742 147200 275798 148000 6 la_input[107]
port 204 nsew signal input
rlabel metal2 s 278226 147200 278282 148000 6 la_input[108]
port 205 nsew signal input
rlabel metal2 s 280802 147200 280858 148000 6 la_input[109]
port 206 nsew signal input
rlabel metal2 s 26606 147200 26662 148000 6 la_input[10]
port 207 nsew signal input
rlabel metal2 s 283378 147200 283434 148000 6 la_input[110]
port 208 nsew signal input
rlabel metal2 s 285954 147200 286010 148000 6 la_input[111]
port 209 nsew signal input
rlabel metal2 s 288530 147200 288586 148000 6 la_input[112]
port 210 nsew signal input
rlabel metal2 s 291106 147200 291162 148000 6 la_input[113]
port 211 nsew signal input
rlabel metal2 s 293682 147200 293738 148000 6 la_input[114]
port 212 nsew signal input
rlabel metal2 s 296258 147200 296314 148000 6 la_input[115]
port 213 nsew signal input
rlabel metal2 s 298834 147200 298890 148000 6 la_input[116]
port 214 nsew signal input
rlabel metal2 s 301410 147200 301466 148000 6 la_input[117]
port 215 nsew signal input
rlabel metal2 s 303986 147200 304042 148000 6 la_input[118]
port 216 nsew signal input
rlabel metal2 s 306562 147200 306618 148000 6 la_input[119]
port 217 nsew signal input
rlabel metal2 s 29182 147200 29238 148000 6 la_input[11]
port 218 nsew signal input
rlabel metal2 s 309046 147200 309102 148000 6 la_input[120]
port 219 nsew signal input
rlabel metal2 s 311622 147200 311678 148000 6 la_input[121]
port 220 nsew signal input
rlabel metal2 s 314198 147200 314254 148000 6 la_input[122]
port 221 nsew signal input
rlabel metal2 s 316774 147200 316830 148000 6 la_input[123]
port 222 nsew signal input
rlabel metal2 s 319350 147200 319406 148000 6 la_input[124]
port 223 nsew signal input
rlabel metal2 s 321926 147200 321982 148000 6 la_input[125]
port 224 nsew signal input
rlabel metal2 s 324502 147200 324558 148000 6 la_input[126]
port 225 nsew signal input
rlabel metal2 s 327078 147200 327134 148000 6 la_input[127]
port 226 nsew signal input
rlabel metal2 s 31666 147200 31722 148000 6 la_input[12]
port 227 nsew signal input
rlabel metal2 s 34242 147200 34298 148000 6 la_input[13]
port 228 nsew signal input
rlabel metal2 s 36818 147200 36874 148000 6 la_input[14]
port 229 nsew signal input
rlabel metal2 s 39394 147200 39450 148000 6 la_input[15]
port 230 nsew signal input
rlabel metal2 s 41970 147200 42026 148000 6 la_input[16]
port 231 nsew signal input
rlabel metal2 s 44546 147200 44602 148000 6 la_input[17]
port 232 nsew signal input
rlabel metal2 s 47122 147200 47178 148000 6 la_input[18]
port 233 nsew signal input
rlabel metal2 s 49698 147200 49754 148000 6 la_input[19]
port 234 nsew signal input
rlabel metal2 s 3422 147200 3478 148000 6 la_input[1]
port 235 nsew signal input
rlabel metal2 s 52274 147200 52330 148000 6 la_input[20]
port 236 nsew signal input
rlabel metal2 s 54850 147200 54906 148000 6 la_input[21]
port 237 nsew signal input
rlabel metal2 s 57426 147200 57482 148000 6 la_input[22]
port 238 nsew signal input
rlabel metal2 s 60002 147200 60058 148000 6 la_input[23]
port 239 nsew signal input
rlabel metal2 s 62486 147200 62542 148000 6 la_input[24]
port 240 nsew signal input
rlabel metal2 s 65062 147200 65118 148000 6 la_input[25]
port 241 nsew signal input
rlabel metal2 s 67638 147200 67694 148000 6 la_input[26]
port 242 nsew signal input
rlabel metal2 s 70214 147200 70270 148000 6 la_input[27]
port 243 nsew signal input
rlabel metal2 s 72790 147200 72846 148000 6 la_input[28]
port 244 nsew signal input
rlabel metal2 s 75366 147200 75422 148000 6 la_input[29]
port 245 nsew signal input
rlabel metal2 s 5998 147200 6054 148000 6 la_input[2]
port 246 nsew signal input
rlabel metal2 s 77942 147200 77998 148000 6 la_input[30]
port 247 nsew signal input
rlabel metal2 s 80518 147200 80574 148000 6 la_input[31]
port 248 nsew signal input
rlabel metal2 s 83094 147200 83150 148000 6 la_input[32]
port 249 nsew signal input
rlabel metal2 s 85670 147200 85726 148000 6 la_input[33]
port 250 nsew signal input
rlabel metal2 s 88246 147200 88302 148000 6 la_input[34]
port 251 nsew signal input
rlabel metal2 s 90822 147200 90878 148000 6 la_input[35]
port 252 nsew signal input
rlabel metal2 s 93306 147200 93362 148000 6 la_input[36]
port 253 nsew signal input
rlabel metal2 s 95882 147200 95938 148000 6 la_input[37]
port 254 nsew signal input
rlabel metal2 s 98458 147200 98514 148000 6 la_input[38]
port 255 nsew signal input
rlabel metal2 s 101034 147200 101090 148000 6 la_input[39]
port 256 nsew signal input
rlabel metal2 s 8574 147200 8630 148000 6 la_input[3]
port 257 nsew signal input
rlabel metal2 s 103610 147200 103666 148000 6 la_input[40]
port 258 nsew signal input
rlabel metal2 s 106186 147200 106242 148000 6 la_input[41]
port 259 nsew signal input
rlabel metal2 s 108762 147200 108818 148000 6 la_input[42]
port 260 nsew signal input
rlabel metal2 s 111338 147200 111394 148000 6 la_input[43]
port 261 nsew signal input
rlabel metal2 s 113914 147200 113970 148000 6 la_input[44]
port 262 nsew signal input
rlabel metal2 s 116490 147200 116546 148000 6 la_input[45]
port 263 nsew signal input
rlabel metal2 s 119066 147200 119122 148000 6 la_input[46]
port 264 nsew signal input
rlabel metal2 s 121642 147200 121698 148000 6 la_input[47]
port 265 nsew signal input
rlabel metal2 s 124126 147200 124182 148000 6 la_input[48]
port 266 nsew signal input
rlabel metal2 s 126702 147200 126758 148000 6 la_input[49]
port 267 nsew signal input
rlabel metal2 s 11150 147200 11206 148000 6 la_input[4]
port 268 nsew signal input
rlabel metal2 s 129278 147200 129334 148000 6 la_input[50]
port 269 nsew signal input
rlabel metal2 s 131854 147200 131910 148000 6 la_input[51]
port 270 nsew signal input
rlabel metal2 s 134430 147200 134486 148000 6 la_input[52]
port 271 nsew signal input
rlabel metal2 s 137006 147200 137062 148000 6 la_input[53]
port 272 nsew signal input
rlabel metal2 s 139582 147200 139638 148000 6 la_input[54]
port 273 nsew signal input
rlabel metal2 s 142158 147200 142214 148000 6 la_input[55]
port 274 nsew signal input
rlabel metal2 s 144734 147200 144790 148000 6 la_input[56]
port 275 nsew signal input
rlabel metal2 s 147310 147200 147366 148000 6 la_input[57]
port 276 nsew signal input
rlabel metal2 s 149886 147200 149942 148000 6 la_input[58]
port 277 nsew signal input
rlabel metal2 s 152462 147200 152518 148000 6 la_input[59]
port 278 nsew signal input
rlabel metal2 s 13726 147200 13782 148000 6 la_input[5]
port 279 nsew signal input
rlabel metal2 s 154946 147200 155002 148000 6 la_input[60]
port 280 nsew signal input
rlabel metal2 s 157522 147200 157578 148000 6 la_input[61]
port 281 nsew signal input
rlabel metal2 s 160098 147200 160154 148000 6 la_input[62]
port 282 nsew signal input
rlabel metal2 s 162674 147200 162730 148000 6 la_input[63]
port 283 nsew signal input
rlabel metal2 s 165250 147200 165306 148000 6 la_input[64]
port 284 nsew signal input
rlabel metal2 s 167826 147200 167882 148000 6 la_input[65]
port 285 nsew signal input
rlabel metal2 s 170402 147200 170458 148000 6 la_input[66]
port 286 nsew signal input
rlabel metal2 s 172978 147200 173034 148000 6 la_input[67]
port 287 nsew signal input
rlabel metal2 s 175554 147200 175610 148000 6 la_input[68]
port 288 nsew signal input
rlabel metal2 s 178130 147200 178186 148000 6 la_input[69]
port 289 nsew signal input
rlabel metal2 s 16302 147200 16358 148000 6 la_input[6]
port 290 nsew signal input
rlabel metal2 s 180706 147200 180762 148000 6 la_input[70]
port 291 nsew signal input
rlabel metal2 s 183282 147200 183338 148000 6 la_input[71]
port 292 nsew signal input
rlabel metal2 s 185766 147200 185822 148000 6 la_input[72]
port 293 nsew signal input
rlabel metal2 s 188342 147200 188398 148000 6 la_input[73]
port 294 nsew signal input
rlabel metal2 s 190918 147200 190974 148000 6 la_input[74]
port 295 nsew signal input
rlabel metal2 s 193494 147200 193550 148000 6 la_input[75]
port 296 nsew signal input
rlabel metal2 s 196070 147200 196126 148000 6 la_input[76]
port 297 nsew signal input
rlabel metal2 s 198646 147200 198702 148000 6 la_input[77]
port 298 nsew signal input
rlabel metal2 s 201222 147200 201278 148000 6 la_input[78]
port 299 nsew signal input
rlabel metal2 s 203798 147200 203854 148000 6 la_input[79]
port 300 nsew signal input
rlabel metal2 s 18878 147200 18934 148000 6 la_input[7]
port 301 nsew signal input
rlabel metal2 s 206374 147200 206430 148000 6 la_input[80]
port 302 nsew signal input
rlabel metal2 s 208950 147200 209006 148000 6 la_input[81]
port 303 nsew signal input
rlabel metal2 s 211526 147200 211582 148000 6 la_input[82]
port 304 nsew signal input
rlabel metal2 s 214102 147200 214158 148000 6 la_input[83]
port 305 nsew signal input
rlabel metal2 s 216586 147200 216642 148000 6 la_input[84]
port 306 nsew signal input
rlabel metal2 s 219162 147200 219218 148000 6 la_input[85]
port 307 nsew signal input
rlabel metal2 s 221738 147200 221794 148000 6 la_input[86]
port 308 nsew signal input
rlabel metal2 s 224314 147200 224370 148000 6 la_input[87]
port 309 nsew signal input
rlabel metal2 s 226890 147200 226946 148000 6 la_input[88]
port 310 nsew signal input
rlabel metal2 s 229466 147200 229522 148000 6 la_input[89]
port 311 nsew signal input
rlabel metal2 s 21454 147200 21510 148000 6 la_input[8]
port 312 nsew signal input
rlabel metal2 s 232042 147200 232098 148000 6 la_input[90]
port 313 nsew signal input
rlabel metal2 s 234618 147200 234674 148000 6 la_input[91]
port 314 nsew signal input
rlabel metal2 s 237194 147200 237250 148000 6 la_input[92]
port 315 nsew signal input
rlabel metal2 s 239770 147200 239826 148000 6 la_input[93]
port 316 nsew signal input
rlabel metal2 s 242346 147200 242402 148000 6 la_input[94]
port 317 nsew signal input
rlabel metal2 s 244922 147200 244978 148000 6 la_input[95]
port 318 nsew signal input
rlabel metal2 s 247406 147200 247462 148000 6 la_input[96]
port 319 nsew signal input
rlabel metal2 s 249982 147200 250038 148000 6 la_input[97]
port 320 nsew signal input
rlabel metal2 s 252558 147200 252614 148000 6 la_input[98]
port 321 nsew signal input
rlabel metal2 s 255134 147200 255190 148000 6 la_input[99]
port 322 nsew signal input
rlabel metal2 s 24030 147200 24086 148000 6 la_input[9]
port 323 nsew signal input
rlabel metal2 s 1490 147200 1546 148000 6 la_oenb[0]
port 324 nsew signal output
rlabel metal2 s 258354 147200 258410 148000 6 la_oenb[100]
port 325 nsew signal output
rlabel metal2 s 260930 147200 260986 148000 6 la_oenb[101]
port 326 nsew signal output
rlabel metal2 s 263506 147200 263562 148000 6 la_oenb[102]
port 327 nsew signal output
rlabel metal2 s 266082 147200 266138 148000 6 la_oenb[103]
port 328 nsew signal output
rlabel metal2 s 268658 147200 268714 148000 6 la_oenb[104]
port 329 nsew signal output
rlabel metal2 s 271234 147200 271290 148000 6 la_oenb[105]
port 330 nsew signal output
rlabel metal2 s 273810 147200 273866 148000 6 la_oenb[106]
port 331 nsew signal output
rlabel metal2 s 276386 147200 276442 148000 6 la_oenb[107]
port 332 nsew signal output
rlabel metal2 s 278870 147200 278926 148000 6 la_oenb[108]
port 333 nsew signal output
rlabel metal2 s 281446 147200 281502 148000 6 la_oenb[109]
port 334 nsew signal output
rlabel metal2 s 27250 147200 27306 148000 6 la_oenb[10]
port 335 nsew signal output
rlabel metal2 s 284022 147200 284078 148000 6 la_oenb[110]
port 336 nsew signal output
rlabel metal2 s 286598 147200 286654 148000 6 la_oenb[111]
port 337 nsew signal output
rlabel metal2 s 289174 147200 289230 148000 6 la_oenb[112]
port 338 nsew signal output
rlabel metal2 s 291750 147200 291806 148000 6 la_oenb[113]
port 339 nsew signal output
rlabel metal2 s 294326 147200 294382 148000 6 la_oenb[114]
port 340 nsew signal output
rlabel metal2 s 296902 147200 296958 148000 6 la_oenb[115]
port 341 nsew signal output
rlabel metal2 s 299478 147200 299534 148000 6 la_oenb[116]
port 342 nsew signal output
rlabel metal2 s 302054 147200 302110 148000 6 la_oenb[117]
port 343 nsew signal output
rlabel metal2 s 304630 147200 304686 148000 6 la_oenb[118]
port 344 nsew signal output
rlabel metal2 s 307206 147200 307262 148000 6 la_oenb[119]
port 345 nsew signal output
rlabel metal2 s 29826 147200 29882 148000 6 la_oenb[11]
port 346 nsew signal output
rlabel metal2 s 309690 147200 309746 148000 6 la_oenb[120]
port 347 nsew signal output
rlabel metal2 s 312266 147200 312322 148000 6 la_oenb[121]
port 348 nsew signal output
rlabel metal2 s 314842 147200 314898 148000 6 la_oenb[122]
port 349 nsew signal output
rlabel metal2 s 317418 147200 317474 148000 6 la_oenb[123]
port 350 nsew signal output
rlabel metal2 s 319994 147200 320050 148000 6 la_oenb[124]
port 351 nsew signal output
rlabel metal2 s 322570 147200 322626 148000 6 la_oenb[125]
port 352 nsew signal output
rlabel metal2 s 325146 147200 325202 148000 6 la_oenb[126]
port 353 nsew signal output
rlabel metal2 s 327722 147200 327778 148000 6 la_oenb[127]
port 354 nsew signal output
rlabel metal2 s 32310 147200 32366 148000 6 la_oenb[12]
port 355 nsew signal output
rlabel metal2 s 34886 147200 34942 148000 6 la_oenb[13]
port 356 nsew signal output
rlabel metal2 s 37462 147200 37518 148000 6 la_oenb[14]
port 357 nsew signal output
rlabel metal2 s 40038 147200 40094 148000 6 la_oenb[15]
port 358 nsew signal output
rlabel metal2 s 42614 147200 42670 148000 6 la_oenb[16]
port 359 nsew signal output
rlabel metal2 s 45190 147200 45246 148000 6 la_oenb[17]
port 360 nsew signal output
rlabel metal2 s 47766 147200 47822 148000 6 la_oenb[18]
port 361 nsew signal output
rlabel metal2 s 50342 147200 50398 148000 6 la_oenb[19]
port 362 nsew signal output
rlabel metal2 s 4066 147200 4122 148000 6 la_oenb[1]
port 363 nsew signal output
rlabel metal2 s 52918 147200 52974 148000 6 la_oenb[20]
port 364 nsew signal output
rlabel metal2 s 55494 147200 55550 148000 6 la_oenb[21]
port 365 nsew signal output
rlabel metal2 s 58070 147200 58126 148000 6 la_oenb[22]
port 366 nsew signal output
rlabel metal2 s 60646 147200 60702 148000 6 la_oenb[23]
port 367 nsew signal output
rlabel metal2 s 63130 147200 63186 148000 6 la_oenb[24]
port 368 nsew signal output
rlabel metal2 s 65706 147200 65762 148000 6 la_oenb[25]
port 369 nsew signal output
rlabel metal2 s 68282 147200 68338 148000 6 la_oenb[26]
port 370 nsew signal output
rlabel metal2 s 70858 147200 70914 148000 6 la_oenb[27]
port 371 nsew signal output
rlabel metal2 s 73434 147200 73490 148000 6 la_oenb[28]
port 372 nsew signal output
rlabel metal2 s 76010 147200 76066 148000 6 la_oenb[29]
port 373 nsew signal output
rlabel metal2 s 6642 147200 6698 148000 6 la_oenb[2]
port 374 nsew signal output
rlabel metal2 s 78586 147200 78642 148000 6 la_oenb[30]
port 375 nsew signal output
rlabel metal2 s 81162 147200 81218 148000 6 la_oenb[31]
port 376 nsew signal output
rlabel metal2 s 83738 147200 83794 148000 6 la_oenb[32]
port 377 nsew signal output
rlabel metal2 s 86314 147200 86370 148000 6 la_oenb[33]
port 378 nsew signal output
rlabel metal2 s 88890 147200 88946 148000 6 la_oenb[34]
port 379 nsew signal output
rlabel metal2 s 91466 147200 91522 148000 6 la_oenb[35]
port 380 nsew signal output
rlabel metal2 s 93950 147200 94006 148000 6 la_oenb[36]
port 381 nsew signal output
rlabel metal2 s 96526 147200 96582 148000 6 la_oenb[37]
port 382 nsew signal output
rlabel metal2 s 99102 147200 99158 148000 6 la_oenb[38]
port 383 nsew signal output
rlabel metal2 s 101678 147200 101734 148000 6 la_oenb[39]
port 384 nsew signal output
rlabel metal2 s 9218 147200 9274 148000 6 la_oenb[3]
port 385 nsew signal output
rlabel metal2 s 104254 147200 104310 148000 6 la_oenb[40]
port 386 nsew signal output
rlabel metal2 s 106830 147200 106886 148000 6 la_oenb[41]
port 387 nsew signal output
rlabel metal2 s 109406 147200 109462 148000 6 la_oenb[42]
port 388 nsew signal output
rlabel metal2 s 111982 147200 112038 148000 6 la_oenb[43]
port 389 nsew signal output
rlabel metal2 s 114558 147200 114614 148000 6 la_oenb[44]
port 390 nsew signal output
rlabel metal2 s 117134 147200 117190 148000 6 la_oenb[45]
port 391 nsew signal output
rlabel metal2 s 119710 147200 119766 148000 6 la_oenb[46]
port 392 nsew signal output
rlabel metal2 s 122286 147200 122342 148000 6 la_oenb[47]
port 393 nsew signal output
rlabel metal2 s 124770 147200 124826 148000 6 la_oenb[48]
port 394 nsew signal output
rlabel metal2 s 127346 147200 127402 148000 6 la_oenb[49]
port 395 nsew signal output
rlabel metal2 s 11794 147200 11850 148000 6 la_oenb[4]
port 396 nsew signal output
rlabel metal2 s 129922 147200 129978 148000 6 la_oenb[50]
port 397 nsew signal output
rlabel metal2 s 132498 147200 132554 148000 6 la_oenb[51]
port 398 nsew signal output
rlabel metal2 s 135074 147200 135130 148000 6 la_oenb[52]
port 399 nsew signal output
rlabel metal2 s 137650 147200 137706 148000 6 la_oenb[53]
port 400 nsew signal output
rlabel metal2 s 140226 147200 140282 148000 6 la_oenb[54]
port 401 nsew signal output
rlabel metal2 s 142802 147200 142858 148000 6 la_oenb[55]
port 402 nsew signal output
rlabel metal2 s 145378 147200 145434 148000 6 la_oenb[56]
port 403 nsew signal output
rlabel metal2 s 147954 147200 148010 148000 6 la_oenb[57]
port 404 nsew signal output
rlabel metal2 s 150530 147200 150586 148000 6 la_oenb[58]
port 405 nsew signal output
rlabel metal2 s 153106 147200 153162 148000 6 la_oenb[59]
port 406 nsew signal output
rlabel metal2 s 14370 147200 14426 148000 6 la_oenb[5]
port 407 nsew signal output
rlabel metal2 s 155590 147200 155646 148000 6 la_oenb[60]
port 408 nsew signal output
rlabel metal2 s 158166 147200 158222 148000 6 la_oenb[61]
port 409 nsew signal output
rlabel metal2 s 160742 147200 160798 148000 6 la_oenb[62]
port 410 nsew signal output
rlabel metal2 s 163318 147200 163374 148000 6 la_oenb[63]
port 411 nsew signal output
rlabel metal2 s 165894 147200 165950 148000 6 la_oenb[64]
port 412 nsew signal output
rlabel metal2 s 168470 147200 168526 148000 6 la_oenb[65]
port 413 nsew signal output
rlabel metal2 s 171046 147200 171102 148000 6 la_oenb[66]
port 414 nsew signal output
rlabel metal2 s 173622 147200 173678 148000 6 la_oenb[67]
port 415 nsew signal output
rlabel metal2 s 176198 147200 176254 148000 6 la_oenb[68]
port 416 nsew signal output
rlabel metal2 s 178774 147200 178830 148000 6 la_oenb[69]
port 417 nsew signal output
rlabel metal2 s 16946 147200 17002 148000 6 la_oenb[6]
port 418 nsew signal output
rlabel metal2 s 181350 147200 181406 148000 6 la_oenb[70]
port 419 nsew signal output
rlabel metal2 s 183926 147200 183982 148000 6 la_oenb[71]
port 420 nsew signal output
rlabel metal2 s 186410 147200 186466 148000 6 la_oenb[72]
port 421 nsew signal output
rlabel metal2 s 188986 147200 189042 148000 6 la_oenb[73]
port 422 nsew signal output
rlabel metal2 s 191562 147200 191618 148000 6 la_oenb[74]
port 423 nsew signal output
rlabel metal2 s 194138 147200 194194 148000 6 la_oenb[75]
port 424 nsew signal output
rlabel metal2 s 196714 147200 196770 148000 6 la_oenb[76]
port 425 nsew signal output
rlabel metal2 s 199290 147200 199346 148000 6 la_oenb[77]
port 426 nsew signal output
rlabel metal2 s 201866 147200 201922 148000 6 la_oenb[78]
port 427 nsew signal output
rlabel metal2 s 204442 147200 204498 148000 6 la_oenb[79]
port 428 nsew signal output
rlabel metal2 s 19522 147200 19578 148000 6 la_oenb[7]
port 429 nsew signal output
rlabel metal2 s 207018 147200 207074 148000 6 la_oenb[80]
port 430 nsew signal output
rlabel metal2 s 209594 147200 209650 148000 6 la_oenb[81]
port 431 nsew signal output
rlabel metal2 s 212170 147200 212226 148000 6 la_oenb[82]
port 432 nsew signal output
rlabel metal2 s 214746 147200 214802 148000 6 la_oenb[83]
port 433 nsew signal output
rlabel metal2 s 217230 147200 217286 148000 6 la_oenb[84]
port 434 nsew signal output
rlabel metal2 s 219806 147200 219862 148000 6 la_oenb[85]
port 435 nsew signal output
rlabel metal2 s 222382 147200 222438 148000 6 la_oenb[86]
port 436 nsew signal output
rlabel metal2 s 224958 147200 225014 148000 6 la_oenb[87]
port 437 nsew signal output
rlabel metal2 s 227534 147200 227590 148000 6 la_oenb[88]
port 438 nsew signal output
rlabel metal2 s 230110 147200 230166 148000 6 la_oenb[89]
port 439 nsew signal output
rlabel metal2 s 22098 147200 22154 148000 6 la_oenb[8]
port 440 nsew signal output
rlabel metal2 s 232686 147200 232742 148000 6 la_oenb[90]
port 441 nsew signal output
rlabel metal2 s 235262 147200 235318 148000 6 la_oenb[91]
port 442 nsew signal output
rlabel metal2 s 237838 147200 237894 148000 6 la_oenb[92]
port 443 nsew signal output
rlabel metal2 s 240414 147200 240470 148000 6 la_oenb[93]
port 444 nsew signal output
rlabel metal2 s 242990 147200 243046 148000 6 la_oenb[94]
port 445 nsew signal output
rlabel metal2 s 245566 147200 245622 148000 6 la_oenb[95]
port 446 nsew signal output
rlabel metal2 s 248050 147200 248106 148000 6 la_oenb[96]
port 447 nsew signal output
rlabel metal2 s 250626 147200 250682 148000 6 la_oenb[97]
port 448 nsew signal output
rlabel metal2 s 253202 147200 253258 148000 6 la_oenb[98]
port 449 nsew signal output
rlabel metal2 s 255778 147200 255834 148000 6 la_oenb[99]
port 450 nsew signal output
rlabel metal2 s 24674 147200 24730 148000 6 la_oenb[9]
port 451 nsew signal output
rlabel metal2 s 2134 147200 2190 148000 6 la_output[0]
port 452 nsew signal output
rlabel metal2 s 258998 147200 259054 148000 6 la_output[100]
port 453 nsew signal output
rlabel metal2 s 261574 147200 261630 148000 6 la_output[101]
port 454 nsew signal output
rlabel metal2 s 264150 147200 264206 148000 6 la_output[102]
port 455 nsew signal output
rlabel metal2 s 266726 147200 266782 148000 6 la_output[103]
port 456 nsew signal output
rlabel metal2 s 269302 147200 269358 148000 6 la_output[104]
port 457 nsew signal output
rlabel metal2 s 271878 147200 271934 148000 6 la_output[105]
port 458 nsew signal output
rlabel metal2 s 274454 147200 274510 148000 6 la_output[106]
port 459 nsew signal output
rlabel metal2 s 277030 147200 277086 148000 6 la_output[107]
port 460 nsew signal output
rlabel metal2 s 279514 147200 279570 148000 6 la_output[108]
port 461 nsew signal output
rlabel metal2 s 282090 147200 282146 148000 6 la_output[109]
port 462 nsew signal output
rlabel metal2 s 27894 147200 27950 148000 6 la_output[10]
port 463 nsew signal output
rlabel metal2 s 284666 147200 284722 148000 6 la_output[110]
port 464 nsew signal output
rlabel metal2 s 287242 147200 287298 148000 6 la_output[111]
port 465 nsew signal output
rlabel metal2 s 289818 147200 289874 148000 6 la_output[112]
port 466 nsew signal output
rlabel metal2 s 292394 147200 292450 148000 6 la_output[113]
port 467 nsew signal output
rlabel metal2 s 294970 147200 295026 148000 6 la_output[114]
port 468 nsew signal output
rlabel metal2 s 297546 147200 297602 148000 6 la_output[115]
port 469 nsew signal output
rlabel metal2 s 300122 147200 300178 148000 6 la_output[116]
port 470 nsew signal output
rlabel metal2 s 302698 147200 302754 148000 6 la_output[117]
port 471 nsew signal output
rlabel metal2 s 305274 147200 305330 148000 6 la_output[118]
port 472 nsew signal output
rlabel metal2 s 307850 147200 307906 148000 6 la_output[119]
port 473 nsew signal output
rlabel metal2 s 30470 147200 30526 148000 6 la_output[11]
port 474 nsew signal output
rlabel metal2 s 310334 147200 310390 148000 6 la_output[120]
port 475 nsew signal output
rlabel metal2 s 312910 147200 312966 148000 6 la_output[121]
port 476 nsew signal output
rlabel metal2 s 315486 147200 315542 148000 6 la_output[122]
port 477 nsew signal output
rlabel metal2 s 318062 147200 318118 148000 6 la_output[123]
port 478 nsew signal output
rlabel metal2 s 320638 147200 320694 148000 6 la_output[124]
port 479 nsew signal output
rlabel metal2 s 323214 147200 323270 148000 6 la_output[125]
port 480 nsew signal output
rlabel metal2 s 325790 147200 325846 148000 6 la_output[126]
port 481 nsew signal output
rlabel metal2 s 328366 147200 328422 148000 6 la_output[127]
port 482 nsew signal output
rlabel metal2 s 32954 147200 33010 148000 6 la_output[12]
port 483 nsew signal output
rlabel metal2 s 35530 147200 35586 148000 6 la_output[13]
port 484 nsew signal output
rlabel metal2 s 38106 147200 38162 148000 6 la_output[14]
port 485 nsew signal output
rlabel metal2 s 40682 147200 40738 148000 6 la_output[15]
port 486 nsew signal output
rlabel metal2 s 43258 147200 43314 148000 6 la_output[16]
port 487 nsew signal output
rlabel metal2 s 45834 147200 45890 148000 6 la_output[17]
port 488 nsew signal output
rlabel metal2 s 48410 147200 48466 148000 6 la_output[18]
port 489 nsew signal output
rlabel metal2 s 50986 147200 51042 148000 6 la_output[19]
port 490 nsew signal output
rlabel metal2 s 4710 147200 4766 148000 6 la_output[1]
port 491 nsew signal output
rlabel metal2 s 53562 147200 53618 148000 6 la_output[20]
port 492 nsew signal output
rlabel metal2 s 56138 147200 56194 148000 6 la_output[21]
port 493 nsew signal output
rlabel metal2 s 58714 147200 58770 148000 6 la_output[22]
port 494 nsew signal output
rlabel metal2 s 61290 147200 61346 148000 6 la_output[23]
port 495 nsew signal output
rlabel metal2 s 63774 147200 63830 148000 6 la_output[24]
port 496 nsew signal output
rlabel metal2 s 66350 147200 66406 148000 6 la_output[25]
port 497 nsew signal output
rlabel metal2 s 68926 147200 68982 148000 6 la_output[26]
port 498 nsew signal output
rlabel metal2 s 71502 147200 71558 148000 6 la_output[27]
port 499 nsew signal output
rlabel metal2 s 74078 147200 74134 148000 6 la_output[28]
port 500 nsew signal output
rlabel metal2 s 76654 147200 76710 148000 6 la_output[29]
port 501 nsew signal output
rlabel metal2 s 7286 147200 7342 148000 6 la_output[2]
port 502 nsew signal output
rlabel metal2 s 79230 147200 79286 148000 6 la_output[30]
port 503 nsew signal output
rlabel metal2 s 81806 147200 81862 148000 6 la_output[31]
port 504 nsew signal output
rlabel metal2 s 84382 147200 84438 148000 6 la_output[32]
port 505 nsew signal output
rlabel metal2 s 86958 147200 87014 148000 6 la_output[33]
port 506 nsew signal output
rlabel metal2 s 89534 147200 89590 148000 6 la_output[34]
port 507 nsew signal output
rlabel metal2 s 92110 147200 92166 148000 6 la_output[35]
port 508 nsew signal output
rlabel metal2 s 94594 147200 94650 148000 6 la_output[36]
port 509 nsew signal output
rlabel metal2 s 97170 147200 97226 148000 6 la_output[37]
port 510 nsew signal output
rlabel metal2 s 99746 147200 99802 148000 6 la_output[38]
port 511 nsew signal output
rlabel metal2 s 102322 147200 102378 148000 6 la_output[39]
port 512 nsew signal output
rlabel metal2 s 9862 147200 9918 148000 6 la_output[3]
port 513 nsew signal output
rlabel metal2 s 104898 147200 104954 148000 6 la_output[40]
port 514 nsew signal output
rlabel metal2 s 107474 147200 107530 148000 6 la_output[41]
port 515 nsew signal output
rlabel metal2 s 110050 147200 110106 148000 6 la_output[42]
port 516 nsew signal output
rlabel metal2 s 112626 147200 112682 148000 6 la_output[43]
port 517 nsew signal output
rlabel metal2 s 115202 147200 115258 148000 6 la_output[44]
port 518 nsew signal output
rlabel metal2 s 117778 147200 117834 148000 6 la_output[45]
port 519 nsew signal output
rlabel metal2 s 120354 147200 120410 148000 6 la_output[46]
port 520 nsew signal output
rlabel metal2 s 122930 147200 122986 148000 6 la_output[47]
port 521 nsew signal output
rlabel metal2 s 125414 147200 125470 148000 6 la_output[48]
port 522 nsew signal output
rlabel metal2 s 127990 147200 128046 148000 6 la_output[49]
port 523 nsew signal output
rlabel metal2 s 12438 147200 12494 148000 6 la_output[4]
port 524 nsew signal output
rlabel metal2 s 130566 147200 130622 148000 6 la_output[50]
port 525 nsew signal output
rlabel metal2 s 133142 147200 133198 148000 6 la_output[51]
port 526 nsew signal output
rlabel metal2 s 135718 147200 135774 148000 6 la_output[52]
port 527 nsew signal output
rlabel metal2 s 138294 147200 138350 148000 6 la_output[53]
port 528 nsew signal output
rlabel metal2 s 140870 147200 140926 148000 6 la_output[54]
port 529 nsew signal output
rlabel metal2 s 143446 147200 143502 148000 6 la_output[55]
port 530 nsew signal output
rlabel metal2 s 146022 147200 146078 148000 6 la_output[56]
port 531 nsew signal output
rlabel metal2 s 148598 147200 148654 148000 6 la_output[57]
port 532 nsew signal output
rlabel metal2 s 151174 147200 151230 148000 6 la_output[58]
port 533 nsew signal output
rlabel metal2 s 153750 147200 153806 148000 6 la_output[59]
port 534 nsew signal output
rlabel metal2 s 15014 147200 15070 148000 6 la_output[5]
port 535 nsew signal output
rlabel metal2 s 156234 147200 156290 148000 6 la_output[60]
port 536 nsew signal output
rlabel metal2 s 158810 147200 158866 148000 6 la_output[61]
port 537 nsew signal output
rlabel metal2 s 161386 147200 161442 148000 6 la_output[62]
port 538 nsew signal output
rlabel metal2 s 163962 147200 164018 148000 6 la_output[63]
port 539 nsew signal output
rlabel metal2 s 166538 147200 166594 148000 6 la_output[64]
port 540 nsew signal output
rlabel metal2 s 169114 147200 169170 148000 6 la_output[65]
port 541 nsew signal output
rlabel metal2 s 171690 147200 171746 148000 6 la_output[66]
port 542 nsew signal output
rlabel metal2 s 174266 147200 174322 148000 6 la_output[67]
port 543 nsew signal output
rlabel metal2 s 176842 147200 176898 148000 6 la_output[68]
port 544 nsew signal output
rlabel metal2 s 179418 147200 179474 148000 6 la_output[69]
port 545 nsew signal output
rlabel metal2 s 17590 147200 17646 148000 6 la_output[6]
port 546 nsew signal output
rlabel metal2 s 181994 147200 182050 148000 6 la_output[70]
port 547 nsew signal output
rlabel metal2 s 184570 147200 184626 148000 6 la_output[71]
port 548 nsew signal output
rlabel metal2 s 187054 147200 187110 148000 6 la_output[72]
port 549 nsew signal output
rlabel metal2 s 189630 147200 189686 148000 6 la_output[73]
port 550 nsew signal output
rlabel metal2 s 192206 147200 192262 148000 6 la_output[74]
port 551 nsew signal output
rlabel metal2 s 194782 147200 194838 148000 6 la_output[75]
port 552 nsew signal output
rlabel metal2 s 197358 147200 197414 148000 6 la_output[76]
port 553 nsew signal output
rlabel metal2 s 199934 147200 199990 148000 6 la_output[77]
port 554 nsew signal output
rlabel metal2 s 202510 147200 202566 148000 6 la_output[78]
port 555 nsew signal output
rlabel metal2 s 205086 147200 205142 148000 6 la_output[79]
port 556 nsew signal output
rlabel metal2 s 20166 147200 20222 148000 6 la_output[7]
port 557 nsew signal output
rlabel metal2 s 207662 147200 207718 148000 6 la_output[80]
port 558 nsew signal output
rlabel metal2 s 210238 147200 210294 148000 6 la_output[81]
port 559 nsew signal output
rlabel metal2 s 212814 147200 212870 148000 6 la_output[82]
port 560 nsew signal output
rlabel metal2 s 215390 147200 215446 148000 6 la_output[83]
port 561 nsew signal output
rlabel metal2 s 217874 147200 217930 148000 6 la_output[84]
port 562 nsew signal output
rlabel metal2 s 220450 147200 220506 148000 6 la_output[85]
port 563 nsew signal output
rlabel metal2 s 223026 147200 223082 148000 6 la_output[86]
port 564 nsew signal output
rlabel metal2 s 225602 147200 225658 148000 6 la_output[87]
port 565 nsew signal output
rlabel metal2 s 228178 147200 228234 148000 6 la_output[88]
port 566 nsew signal output
rlabel metal2 s 230754 147200 230810 148000 6 la_output[89]
port 567 nsew signal output
rlabel metal2 s 22742 147200 22798 148000 6 la_output[8]
port 568 nsew signal output
rlabel metal2 s 233330 147200 233386 148000 6 la_output[90]
port 569 nsew signal output
rlabel metal2 s 235906 147200 235962 148000 6 la_output[91]
port 570 nsew signal output
rlabel metal2 s 238482 147200 238538 148000 6 la_output[92]
port 571 nsew signal output
rlabel metal2 s 241058 147200 241114 148000 6 la_output[93]
port 572 nsew signal output
rlabel metal2 s 243634 147200 243690 148000 6 la_output[94]
port 573 nsew signal output
rlabel metal2 s 246210 147200 246266 148000 6 la_output[95]
port 574 nsew signal output
rlabel metal2 s 248694 147200 248750 148000 6 la_output[96]
port 575 nsew signal output
rlabel metal2 s 251270 147200 251326 148000 6 la_output[97]
port 576 nsew signal output
rlabel metal2 s 253846 147200 253902 148000 6 la_output[98]
port 577 nsew signal output
rlabel metal2 s 256422 147200 256478 148000 6 la_output[99]
port 578 nsew signal output
rlabel metal2 s 25318 147200 25374 148000 6 la_output[9]
port 579 nsew signal output
rlabel metal3 s 0 62432 800 62552 6 mem_addr[0]
port 580 nsew signal output
rlabel metal3 s 0 64336 800 64456 6 mem_addr[1]
port 581 nsew signal output
rlabel metal3 s 0 66240 800 66360 6 mem_addr[2]
port 582 nsew signal output
rlabel metal3 s 0 68144 800 68264 6 mem_addr[3]
port 583 nsew signal output
rlabel metal3 s 0 70048 800 70168 6 mem_addr[4]
port 584 nsew signal output
rlabel metal3 s 0 71952 800 72072 6 mem_addr[5]
port 585 nsew signal output
rlabel metal3 s 0 73856 800 73976 6 mem_addr[6]
port 586 nsew signal output
rlabel metal3 s 0 75896 800 76016 6 mem_addr[7]
port 587 nsew signal output
rlabel metal3 s 0 85416 800 85536 6 mem_ena
port 588 nsew signal output
rlabel metal3 s 0 87320 800 87440 6 mem_rdata[0]
port 589 nsew signal input
rlabel metal3 s 0 106632 800 106752 6 mem_rdata[10]
port 590 nsew signal input
rlabel metal3 s 0 108536 800 108656 6 mem_rdata[11]
port 591 nsew signal input
rlabel metal3 s 0 110440 800 110560 6 mem_rdata[12]
port 592 nsew signal input
rlabel metal3 s 0 112344 800 112464 6 mem_rdata[13]
port 593 nsew signal input
rlabel metal3 s 0 114248 800 114368 6 mem_rdata[14]
port 594 nsew signal input
rlabel metal3 s 0 116152 800 116272 6 mem_rdata[15]
port 595 nsew signal input
rlabel metal3 s 0 118056 800 118176 6 mem_rdata[16]
port 596 nsew signal input
rlabel metal3 s 0 120096 800 120216 6 mem_rdata[17]
port 597 nsew signal input
rlabel metal3 s 0 122000 800 122120 6 mem_rdata[18]
port 598 nsew signal input
rlabel metal3 s 0 123904 800 124024 6 mem_rdata[19]
port 599 nsew signal input
rlabel metal3 s 0 89224 800 89344 6 mem_rdata[1]
port 600 nsew signal input
rlabel metal3 s 0 125808 800 125928 6 mem_rdata[20]
port 601 nsew signal input
rlabel metal3 s 0 127712 800 127832 6 mem_rdata[21]
port 602 nsew signal input
rlabel metal3 s 0 129616 800 129736 6 mem_rdata[22]
port 603 nsew signal input
rlabel metal3 s 0 131520 800 131640 6 mem_rdata[23]
port 604 nsew signal input
rlabel metal3 s 0 133424 800 133544 6 mem_rdata[24]
port 605 nsew signal input
rlabel metal3 s 0 135464 800 135584 6 mem_rdata[25]
port 606 nsew signal input
rlabel metal3 s 0 137368 800 137488 6 mem_rdata[26]
port 607 nsew signal input
rlabel metal3 s 0 139272 800 139392 6 mem_rdata[27]
port 608 nsew signal input
rlabel metal3 s 0 141176 800 141296 6 mem_rdata[28]
port 609 nsew signal input
rlabel metal3 s 0 143080 800 143200 6 mem_rdata[29]
port 610 nsew signal input
rlabel metal3 s 0 91264 800 91384 6 mem_rdata[2]
port 611 nsew signal input
rlabel metal3 s 0 144984 800 145104 6 mem_rdata[30]
port 612 nsew signal input
rlabel metal3 s 0 146888 800 147008 6 mem_rdata[31]
port 613 nsew signal input
rlabel metal3 s 0 93168 800 93288 6 mem_rdata[3]
port 614 nsew signal input
rlabel metal3 s 0 95072 800 95192 6 mem_rdata[4]
port 615 nsew signal input
rlabel metal3 s 0 96976 800 97096 6 mem_rdata[5]
port 616 nsew signal input
rlabel metal3 s 0 98880 800 99000 6 mem_rdata[6]
port 617 nsew signal input
rlabel metal3 s 0 100784 800 100904 6 mem_rdata[7]
port 618 nsew signal input
rlabel metal3 s 0 102688 800 102808 6 mem_rdata[8]
port 619 nsew signal input
rlabel metal3 s 0 104728 800 104848 6 mem_rdata[9]
port 620 nsew signal input
rlabel metal3 s 0 960 800 1080 6 mem_wdata[0]
port 621 nsew signal output
rlabel metal3 s 0 20136 800 20256 6 mem_wdata[10]
port 622 nsew signal output
rlabel metal3 s 0 22040 800 22160 6 mem_wdata[11]
port 623 nsew signal output
rlabel metal3 s 0 23944 800 24064 6 mem_wdata[12]
port 624 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 mem_wdata[13]
port 625 nsew signal output
rlabel metal3 s 0 27752 800 27872 6 mem_wdata[14]
port 626 nsew signal output
rlabel metal3 s 0 29656 800 29776 6 mem_wdata[15]
port 627 nsew signal output
rlabel metal3 s 0 31696 800 31816 6 mem_wdata[16]
port 628 nsew signal output
rlabel metal3 s 0 33600 800 33720 6 mem_wdata[17]
port 629 nsew signal output
rlabel metal3 s 0 35504 800 35624 6 mem_wdata[18]
port 630 nsew signal output
rlabel metal3 s 0 37408 800 37528 6 mem_wdata[19]
port 631 nsew signal output
rlabel metal3 s 0 2864 800 2984 6 mem_wdata[1]
port 632 nsew signal output
rlabel metal3 s 0 39312 800 39432 6 mem_wdata[20]
port 633 nsew signal output
rlabel metal3 s 0 41216 800 41336 6 mem_wdata[21]
port 634 nsew signal output
rlabel metal3 s 0 43120 800 43240 6 mem_wdata[22]
port 635 nsew signal output
rlabel metal3 s 0 45024 800 45144 6 mem_wdata[23]
port 636 nsew signal output
rlabel metal3 s 0 47064 800 47184 6 mem_wdata[24]
port 637 nsew signal output
rlabel metal3 s 0 48968 800 49088 6 mem_wdata[25]
port 638 nsew signal output
rlabel metal3 s 0 50872 800 50992 6 mem_wdata[26]
port 639 nsew signal output
rlabel metal3 s 0 52776 800 52896 6 mem_wdata[27]
port 640 nsew signal output
rlabel metal3 s 0 54680 800 54800 6 mem_wdata[28]
port 641 nsew signal output
rlabel metal3 s 0 56584 800 56704 6 mem_wdata[29]
port 642 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 mem_wdata[2]
port 643 nsew signal output
rlabel metal3 s 0 58488 800 58608 6 mem_wdata[30]
port 644 nsew signal output
rlabel metal3 s 0 60528 800 60648 6 mem_wdata[31]
port 645 nsew signal output
rlabel metal3 s 0 6672 800 6792 6 mem_wdata[3]
port 646 nsew signal output
rlabel metal3 s 0 8576 800 8696 6 mem_wdata[4]
port 647 nsew signal output
rlabel metal3 s 0 10480 800 10600 6 mem_wdata[5]
port 648 nsew signal output
rlabel metal3 s 0 12384 800 12504 6 mem_wdata[6]
port 649 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 mem_wdata[7]
port 650 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 mem_wdata[8]
port 651 nsew signal output
rlabel metal3 s 0 18232 800 18352 6 mem_wdata[9]
port 652 nsew signal output
rlabel metal3 s 0 77800 800 77920 6 mem_wen[0]
port 653 nsew signal output
rlabel metal3 s 0 79704 800 79824 6 mem_wen[1]
port 654 nsew signal output
rlabel metal3 s 0 81608 800 81728 6 mem_wen[2]
port 655 nsew signal output
rlabel metal3 s 0 83512 800 83632 6 mem_wen[3]
port 656 nsew signal output
rlabel metal2 s 329010 147200 329066 148000 6 mprj_ack_i
port 657 nsew signal input
rlabel metal2 s 332230 147200 332286 148000 6 mprj_adr_o[0]
port 658 nsew signal output
rlabel metal2 s 354034 147200 354090 148000 6 mprj_adr_o[10]
port 659 nsew signal output
rlabel metal2 s 355966 147200 356022 148000 6 mprj_adr_o[11]
port 660 nsew signal output
rlabel metal2 s 357898 147200 357954 148000 6 mprj_adr_o[12]
port 661 nsew signal output
rlabel metal2 s 359830 147200 359886 148000 6 mprj_adr_o[13]
port 662 nsew signal output
rlabel metal2 s 361762 147200 361818 148000 6 mprj_adr_o[14]
port 663 nsew signal output
rlabel metal2 s 363694 147200 363750 148000 6 mprj_adr_o[15]
port 664 nsew signal output
rlabel metal2 s 365626 147200 365682 148000 6 mprj_adr_o[16]
port 665 nsew signal output
rlabel metal2 s 367558 147200 367614 148000 6 mprj_adr_o[17]
port 666 nsew signal output
rlabel metal2 s 369490 147200 369546 148000 6 mprj_adr_o[18]
port 667 nsew signal output
rlabel metal2 s 371330 147200 371386 148000 6 mprj_adr_o[19]
port 668 nsew signal output
rlabel metal2 s 334806 147200 334862 148000 6 mprj_adr_o[1]
port 669 nsew signal output
rlabel metal2 s 373262 147200 373318 148000 6 mprj_adr_o[20]
port 670 nsew signal output
rlabel metal2 s 375194 147200 375250 148000 6 mprj_adr_o[21]
port 671 nsew signal output
rlabel metal2 s 377126 147200 377182 148000 6 mprj_adr_o[22]
port 672 nsew signal output
rlabel metal2 s 379058 147200 379114 148000 6 mprj_adr_o[23]
port 673 nsew signal output
rlabel metal2 s 380990 147200 381046 148000 6 mprj_adr_o[24]
port 674 nsew signal output
rlabel metal2 s 382922 147200 382978 148000 6 mprj_adr_o[25]
port 675 nsew signal output
rlabel metal2 s 384854 147200 384910 148000 6 mprj_adr_o[26]
port 676 nsew signal output
rlabel metal2 s 386786 147200 386842 148000 6 mprj_adr_o[27]
port 677 nsew signal output
rlabel metal2 s 388718 147200 388774 148000 6 mprj_adr_o[28]
port 678 nsew signal output
rlabel metal2 s 390650 147200 390706 148000 6 mprj_adr_o[29]
port 679 nsew signal output
rlabel metal2 s 337382 147200 337438 148000 6 mprj_adr_o[2]
port 680 nsew signal output
rlabel metal2 s 392582 147200 392638 148000 6 mprj_adr_o[30]
port 681 nsew signal output
rlabel metal2 s 394514 147200 394570 148000 6 mprj_adr_o[31]
port 682 nsew signal output
rlabel metal2 s 339866 147200 339922 148000 6 mprj_adr_o[3]
port 683 nsew signal output
rlabel metal2 s 342442 147200 342498 148000 6 mprj_adr_o[4]
port 684 nsew signal output
rlabel metal2 s 344374 147200 344430 148000 6 mprj_adr_o[5]
port 685 nsew signal output
rlabel metal2 s 346306 147200 346362 148000 6 mprj_adr_o[6]
port 686 nsew signal output
rlabel metal2 s 348238 147200 348294 148000 6 mprj_adr_o[7]
port 687 nsew signal output
rlabel metal2 s 350170 147200 350226 148000 6 mprj_adr_o[8]
port 688 nsew signal output
rlabel metal2 s 352102 147200 352158 148000 6 mprj_adr_o[9]
port 689 nsew signal output
rlabel metal2 s 329654 147200 329710 148000 6 mprj_cyc_o
port 690 nsew signal output
rlabel metal2 s 332874 147200 332930 148000 6 mprj_dat_i[0]
port 691 nsew signal input
rlabel metal2 s 354678 147200 354734 148000 6 mprj_dat_i[10]
port 692 nsew signal input
rlabel metal2 s 356610 147200 356666 148000 6 mprj_dat_i[11]
port 693 nsew signal input
rlabel metal2 s 358542 147200 358598 148000 6 mprj_dat_i[12]
port 694 nsew signal input
rlabel metal2 s 360474 147200 360530 148000 6 mprj_dat_i[13]
port 695 nsew signal input
rlabel metal2 s 362406 147200 362462 148000 6 mprj_dat_i[14]
port 696 nsew signal input
rlabel metal2 s 364338 147200 364394 148000 6 mprj_dat_i[15]
port 697 nsew signal input
rlabel metal2 s 366270 147200 366326 148000 6 mprj_dat_i[16]
port 698 nsew signal input
rlabel metal2 s 368202 147200 368258 148000 6 mprj_dat_i[17]
port 699 nsew signal input
rlabel metal2 s 370042 147200 370098 148000 6 mprj_dat_i[18]
port 700 nsew signal input
rlabel metal2 s 371974 147200 372030 148000 6 mprj_dat_i[19]
port 701 nsew signal input
rlabel metal2 s 335450 147200 335506 148000 6 mprj_dat_i[1]
port 702 nsew signal input
rlabel metal2 s 373906 147200 373962 148000 6 mprj_dat_i[20]
port 703 nsew signal input
rlabel metal2 s 375838 147200 375894 148000 6 mprj_dat_i[21]
port 704 nsew signal input
rlabel metal2 s 377770 147200 377826 148000 6 mprj_dat_i[22]
port 705 nsew signal input
rlabel metal2 s 379702 147200 379758 148000 6 mprj_dat_i[23]
port 706 nsew signal input
rlabel metal2 s 381634 147200 381690 148000 6 mprj_dat_i[24]
port 707 nsew signal input
rlabel metal2 s 383566 147200 383622 148000 6 mprj_dat_i[25]
port 708 nsew signal input
rlabel metal2 s 385498 147200 385554 148000 6 mprj_dat_i[26]
port 709 nsew signal input
rlabel metal2 s 387430 147200 387486 148000 6 mprj_dat_i[27]
port 710 nsew signal input
rlabel metal2 s 389362 147200 389418 148000 6 mprj_dat_i[28]
port 711 nsew signal input
rlabel metal2 s 391294 147200 391350 148000 6 mprj_dat_i[29]
port 712 nsew signal input
rlabel metal2 s 338026 147200 338082 148000 6 mprj_dat_i[2]
port 713 nsew signal input
rlabel metal2 s 393226 147200 393282 148000 6 mprj_dat_i[30]
port 714 nsew signal input
rlabel metal2 s 395158 147200 395214 148000 6 mprj_dat_i[31]
port 715 nsew signal input
rlabel metal2 s 340510 147200 340566 148000 6 mprj_dat_i[3]
port 716 nsew signal input
rlabel metal2 s 343086 147200 343142 148000 6 mprj_dat_i[4]
port 717 nsew signal input
rlabel metal2 s 345018 147200 345074 148000 6 mprj_dat_i[5]
port 718 nsew signal input
rlabel metal2 s 346950 147200 347006 148000 6 mprj_dat_i[6]
port 719 nsew signal input
rlabel metal2 s 348882 147200 348938 148000 6 mprj_dat_i[7]
port 720 nsew signal input
rlabel metal2 s 350814 147200 350870 148000 6 mprj_dat_i[8]
port 721 nsew signal input
rlabel metal2 s 352746 147200 352802 148000 6 mprj_dat_i[9]
port 722 nsew signal input
rlabel metal2 s 333518 147200 333574 148000 6 mprj_dat_o[0]
port 723 nsew signal output
rlabel metal2 s 355322 147200 355378 148000 6 mprj_dat_o[10]
port 724 nsew signal output
rlabel metal2 s 357254 147200 357310 148000 6 mprj_dat_o[11]
port 725 nsew signal output
rlabel metal2 s 359186 147200 359242 148000 6 mprj_dat_o[12]
port 726 nsew signal output
rlabel metal2 s 361118 147200 361174 148000 6 mprj_dat_o[13]
port 727 nsew signal output
rlabel metal2 s 363050 147200 363106 148000 6 mprj_dat_o[14]
port 728 nsew signal output
rlabel metal2 s 364982 147200 365038 148000 6 mprj_dat_o[15]
port 729 nsew signal output
rlabel metal2 s 366914 147200 366970 148000 6 mprj_dat_o[16]
port 730 nsew signal output
rlabel metal2 s 368846 147200 368902 148000 6 mprj_dat_o[17]
port 731 nsew signal output
rlabel metal2 s 370686 147200 370742 148000 6 mprj_dat_o[18]
port 732 nsew signal output
rlabel metal2 s 372618 147200 372674 148000 6 mprj_dat_o[19]
port 733 nsew signal output
rlabel metal2 s 336094 147200 336150 148000 6 mprj_dat_o[1]
port 734 nsew signal output
rlabel metal2 s 374550 147200 374606 148000 6 mprj_dat_o[20]
port 735 nsew signal output
rlabel metal2 s 376482 147200 376538 148000 6 mprj_dat_o[21]
port 736 nsew signal output
rlabel metal2 s 378414 147200 378470 148000 6 mprj_dat_o[22]
port 737 nsew signal output
rlabel metal2 s 380346 147200 380402 148000 6 mprj_dat_o[23]
port 738 nsew signal output
rlabel metal2 s 382278 147200 382334 148000 6 mprj_dat_o[24]
port 739 nsew signal output
rlabel metal2 s 384210 147200 384266 148000 6 mprj_dat_o[25]
port 740 nsew signal output
rlabel metal2 s 386142 147200 386198 148000 6 mprj_dat_o[26]
port 741 nsew signal output
rlabel metal2 s 388074 147200 388130 148000 6 mprj_dat_o[27]
port 742 nsew signal output
rlabel metal2 s 390006 147200 390062 148000 6 mprj_dat_o[28]
port 743 nsew signal output
rlabel metal2 s 391938 147200 391994 148000 6 mprj_dat_o[29]
port 744 nsew signal output
rlabel metal2 s 338670 147200 338726 148000 6 mprj_dat_o[2]
port 745 nsew signal output
rlabel metal2 s 393870 147200 393926 148000 6 mprj_dat_o[30]
port 746 nsew signal output
rlabel metal2 s 395802 147200 395858 148000 6 mprj_dat_o[31]
port 747 nsew signal output
rlabel metal2 s 341154 147200 341210 148000 6 mprj_dat_o[3]
port 748 nsew signal output
rlabel metal2 s 343730 147200 343786 148000 6 mprj_dat_o[4]
port 749 nsew signal output
rlabel metal2 s 345662 147200 345718 148000 6 mprj_dat_o[5]
port 750 nsew signal output
rlabel metal2 s 347594 147200 347650 148000 6 mprj_dat_o[6]
port 751 nsew signal output
rlabel metal2 s 349526 147200 349582 148000 6 mprj_dat_o[7]
port 752 nsew signal output
rlabel metal2 s 351458 147200 351514 148000 6 mprj_dat_o[8]
port 753 nsew signal output
rlabel metal2 s 353390 147200 353446 148000 6 mprj_dat_o[9]
port 754 nsew signal output
rlabel metal2 s 334162 147200 334218 148000 6 mprj_sel_o[0]
port 755 nsew signal output
rlabel metal2 s 336738 147200 336794 148000 6 mprj_sel_o[1]
port 756 nsew signal output
rlabel metal2 s 339222 147200 339278 148000 6 mprj_sel_o[2]
port 757 nsew signal output
rlabel metal2 s 341798 147200 341854 148000 6 mprj_sel_o[3]
port 758 nsew signal output
rlabel metal2 s 330298 147200 330354 148000 6 mprj_stb_o
port 759 nsew signal output
rlabel metal2 s 330942 147200 330998 148000 6 mprj_wb_iena
port 760 nsew signal output
rlabel metal2 s 331586 147200 331642 148000 6 mprj_we_o
port 761 nsew signal output
rlabel metal3 s 399200 81472 400000 81592 6 qspi_enabled
port 762 nsew signal output
rlabel metal2 s 74906 0 74962 800 6 resetn
port 763 nsew signal input
rlabel metal3 s 399200 76032 400000 76152 6 ser_rx
port 764 nsew signal input
rlabel metal3 s 399200 77392 400000 77512 6 ser_tx
port 765 nsew signal output
rlabel metal3 s 399200 73176 400000 73296 6 spi_csb
port 766 nsew signal output
rlabel metal3 s 399200 78752 400000 78872 6 spi_enabled
port 767 nsew signal output
rlabel metal3 s 399200 71816 400000 71936 6 spi_sck
port 768 nsew signal output
rlabel metal3 s 399200 74672 400000 74792 6 spi_sdi
port 769 nsew signal input
rlabel metal3 s 399200 70456 400000 70576 6 spi_sdo
port 770 nsew signal output
rlabel metal3 s 399200 69096 400000 69216 6 spi_sdoenb
port 771 nsew signal output
rlabel metal3 s 399200 2048 400000 2168 6 sram_ro_addr[0]
port 772 nsew signal input
rlabel metal3 s 399200 3408 400000 3528 6 sram_ro_addr[1]
port 773 nsew signal input
rlabel metal3 s 399200 4768 400000 4888 6 sram_ro_addr[2]
port 774 nsew signal input
rlabel metal3 s 399200 6128 400000 6248 6 sram_ro_addr[3]
port 775 nsew signal input
rlabel metal3 s 399200 7488 400000 7608 6 sram_ro_addr[4]
port 776 nsew signal input
rlabel metal3 s 399200 8848 400000 8968 6 sram_ro_addr[5]
port 777 nsew signal input
rlabel metal3 s 399200 10208 400000 10328 6 sram_ro_addr[6]
port 778 nsew signal input
rlabel metal3 s 399200 11568 400000 11688 6 sram_ro_addr[7]
port 779 nsew signal input
rlabel metal3 s 399200 12928 400000 13048 6 sram_ro_clk
port 780 nsew signal input
rlabel metal3 s 399200 688 400000 808 6 sram_ro_csb
port 781 nsew signal input
rlabel metal3 s 399200 14288 400000 14408 6 sram_ro_data[0]
port 782 nsew signal output
rlabel metal3 s 399200 28024 400000 28144 6 sram_ro_data[10]
port 783 nsew signal output
rlabel metal3 s 399200 29384 400000 29504 6 sram_ro_data[11]
port 784 nsew signal output
rlabel metal3 s 399200 30744 400000 30864 6 sram_ro_data[12]
port 785 nsew signal output
rlabel metal3 s 399200 32104 400000 32224 6 sram_ro_data[13]
port 786 nsew signal output
rlabel metal3 s 399200 33464 400000 33584 6 sram_ro_data[14]
port 787 nsew signal output
rlabel metal3 s 399200 34824 400000 34944 6 sram_ro_data[15]
port 788 nsew signal output
rlabel metal3 s 399200 36184 400000 36304 6 sram_ro_data[16]
port 789 nsew signal output
rlabel metal3 s 399200 37680 400000 37800 6 sram_ro_data[17]
port 790 nsew signal output
rlabel metal3 s 399200 39040 400000 39160 6 sram_ro_data[18]
port 791 nsew signal output
rlabel metal3 s 399200 40400 400000 40520 6 sram_ro_data[19]
port 792 nsew signal output
rlabel metal3 s 399200 15648 400000 15768 6 sram_ro_data[1]
port 793 nsew signal output
rlabel metal3 s 399200 41760 400000 41880 6 sram_ro_data[20]
port 794 nsew signal output
rlabel metal3 s 399200 43120 400000 43240 6 sram_ro_data[21]
port 795 nsew signal output
rlabel metal3 s 399200 44480 400000 44600 6 sram_ro_data[22]
port 796 nsew signal output
rlabel metal3 s 399200 45840 400000 45960 6 sram_ro_data[23]
port 797 nsew signal output
rlabel metal3 s 399200 47200 400000 47320 6 sram_ro_data[24]
port 798 nsew signal output
rlabel metal3 s 399200 48560 400000 48680 6 sram_ro_data[25]
port 799 nsew signal output
rlabel metal3 s 399200 49920 400000 50040 6 sram_ro_data[26]
port 800 nsew signal output
rlabel metal3 s 399200 51280 400000 51400 6 sram_ro_data[27]
port 801 nsew signal output
rlabel metal3 s 399200 52640 400000 52760 6 sram_ro_data[28]
port 802 nsew signal output
rlabel metal3 s 399200 54000 400000 54120 6 sram_ro_data[29]
port 803 nsew signal output
rlabel metal3 s 399200 17008 400000 17128 6 sram_ro_data[2]
port 804 nsew signal output
rlabel metal3 s 399200 55360 400000 55480 6 sram_ro_data[30]
port 805 nsew signal output
rlabel metal3 s 399200 56856 400000 56976 6 sram_ro_data[31]
port 806 nsew signal output
rlabel metal3 s 399200 18368 400000 18488 6 sram_ro_data[3]
port 807 nsew signal output
rlabel metal3 s 399200 19864 400000 19984 6 sram_ro_data[4]
port 808 nsew signal output
rlabel metal3 s 399200 21224 400000 21344 6 sram_ro_data[5]
port 809 nsew signal output
rlabel metal3 s 399200 22584 400000 22704 6 sram_ro_data[6]
port 810 nsew signal output
rlabel metal3 s 399200 23944 400000 24064 6 sram_ro_data[7]
port 811 nsew signal output
rlabel metal3 s 399200 25304 400000 25424 6 sram_ro_data[8]
port 812 nsew signal output
rlabel metal3 s 399200 26664 400000 26784 6 sram_ro_data[9]
port 813 nsew signal output
rlabel metal3 s 399200 63656 400000 63776 6 trap
port 814 nsew signal output
rlabel metal3 s 399200 80112 400000 80232 6 uart_enabled
port 815 nsew signal output
rlabel metal2 s 396446 147200 396502 148000 6 user_irq_ena[0]
port 816 nsew signal output
rlabel metal2 s 397090 147200 397146 148000 6 user_irq_ena[1]
port 817 nsew signal output
rlabel metal2 s 397734 147200 397790 148000 6 user_irq_ena[2]
port 818 nsew signal output
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 400000 148000
string LEFview TRUE
string GDS_FILE ../gds/mgmt_core.gds
string GDS_END 120940904
string GDS_START 16949608
<< end >>

