magic
tech sky130A
magscale 1 2
timestamp 1637416515
<< metal1 >>
rect 277136 160160 277394 160188
rect 83642 160012 83648 160064
rect 83700 160052 83706 160064
rect 166994 160052 167000 160064
rect 83700 160024 167000 160052
rect 83700 160012 83706 160024
rect 166994 160012 167000 160024
rect 167052 160012 167058 160064
rect 170214 160012 170220 160064
rect 170272 160052 170278 160064
rect 198918 160052 198924 160064
rect 170272 160024 198924 160052
rect 170272 160012 170278 160024
rect 198918 160012 198924 160024
rect 198976 160012 198982 160064
rect 211430 160012 211436 160064
rect 211488 160052 211494 160064
rect 277136 160052 277164 160160
rect 211488 160024 277164 160052
rect 277366 160052 277394 160160
rect 330662 160120 330668 160132
rect 327368 160092 330668 160120
rect 280338 160052 280344 160064
rect 277366 160024 280344 160052
rect 211488 160012 211494 160024
rect 280338 160012 280344 160024
rect 280396 160012 280402 160064
rect 281258 160012 281264 160064
rect 281316 160052 281322 160064
rect 327368 160052 327396 160092
rect 330662 160080 330668 160092
rect 330720 160080 330726 160132
rect 335354 160120 335360 160132
rect 335004 160092 335360 160120
rect 281316 160024 327396 160052
rect 281316 160012 281322 160024
rect 327442 160012 327448 160064
rect 327500 160052 327506 160064
rect 334158 160052 334164 160064
rect 327500 160024 334164 160052
rect 327500 160012 327506 160024
rect 334158 160012 334164 160024
rect 334216 160012 334222 160064
rect 334250 160012 334256 160064
rect 334308 160052 334314 160064
rect 335004 160052 335032 160092
rect 335354 160080 335360 160092
rect 335412 160080 335418 160132
rect 334308 160024 335032 160052
rect 334308 160012 334314 160024
rect 335078 160012 335084 160064
rect 335136 160052 335142 160064
rect 374730 160052 374736 160064
rect 335136 160024 374736 160052
rect 335136 160012 335142 160024
rect 374730 160012 374736 160024
rect 374788 160012 374794 160064
rect 378870 160012 378876 160064
rect 378928 160052 378934 160064
rect 398098 160052 398104 160064
rect 378928 160024 398104 160052
rect 378928 160012 378934 160024
rect 398098 160012 398104 160024
rect 398156 160012 398162 160064
rect 404078 160012 404084 160064
rect 404136 160052 404142 160064
rect 427354 160052 427360 160064
rect 404136 160024 427360 160052
rect 404136 160012 404142 160024
rect 427354 160012 427360 160024
rect 427412 160012 427418 160064
rect 25590 159944 25596 159996
rect 25648 159984 25654 159996
rect 109126 159984 109132 159996
rect 25648 159956 109132 159984
rect 25648 159944 25654 159956
rect 109126 159944 109132 159956
rect 109184 159944 109190 159996
rect 117222 159944 117228 159996
rect 117280 159984 117286 159996
rect 191742 159984 191748 159996
rect 117280 159956 191748 159984
rect 117280 159944 117286 159956
rect 191742 159944 191748 159956
rect 191800 159944 191806 159996
rect 197998 159944 198004 159996
rect 198056 159984 198062 159996
rect 270126 159984 270132 159996
rect 198056 159956 270132 159984
rect 198056 159944 198062 159956
rect 270126 159944 270132 159956
rect 270184 159944 270190 159996
rect 271230 159944 271236 159996
rect 271288 159984 271294 159996
rect 272794 159984 272800 159996
rect 271288 159956 272800 159984
rect 271288 159944 271294 159956
rect 272794 159944 272800 159956
rect 272852 159944 272858 159996
rect 275370 159944 275376 159996
rect 275428 159984 275434 159996
rect 329098 159984 329104 159996
rect 275428 159956 329104 159984
rect 275428 159944 275434 159956
rect 329098 159944 329104 159956
rect 329156 159944 329162 159996
rect 329190 159944 329196 159996
rect 329248 159984 329254 159996
rect 370222 159984 370228 159996
rect 329248 159956 370228 159984
rect 329248 159944 329254 159956
rect 370222 159944 370228 159956
rect 370280 159944 370286 159996
rect 374638 159944 374644 159996
rect 374696 159984 374702 159996
rect 388438 159984 388444 159996
rect 374696 159956 388444 159984
rect 374696 159944 374702 159956
rect 388438 159944 388444 159956
rect 388496 159944 388502 159996
rect 389818 159944 389824 159996
rect 389876 159984 389882 159996
rect 413830 159984 413836 159996
rect 389876 159956 413836 159984
rect 389876 159944 389882 159956
rect 413830 159944 413836 159956
rect 413888 159944 413894 159996
rect 70118 159876 70124 159928
rect 70176 159916 70182 159928
rect 148778 159916 148784 159928
rect 70176 159888 148784 159916
rect 70176 159876 70182 159888
rect 148778 159876 148784 159888
rect 148836 159876 148842 159928
rect 148870 159876 148876 159928
rect 148928 159916 148934 159928
rect 148928 159888 150664 159916
rect 148928 159876 148934 159888
rect 56686 159808 56692 159860
rect 56744 159848 56750 159860
rect 136542 159848 136548 159860
rect 56744 159820 136548 159848
rect 56744 159808 56750 159820
rect 136542 159808 136548 159820
rect 136600 159808 136606 159860
rect 136634 159808 136640 159860
rect 136692 159848 136698 159860
rect 136692 159820 146984 159848
rect 136692 159808 136698 159820
rect 63402 159740 63408 159792
rect 63460 159780 63466 159792
rect 146846 159780 146852 159792
rect 63460 159752 146852 159780
rect 63460 159740 63466 159752
rect 146846 159740 146852 159752
rect 146904 159740 146910 159792
rect 18874 159672 18880 159724
rect 18932 159712 18938 159724
rect 107102 159712 107108 159724
rect 18932 159684 107108 159712
rect 18932 159672 18938 159684
rect 107102 159672 107108 159684
rect 107160 159672 107166 159724
rect 109678 159672 109684 159724
rect 109736 159712 109742 159724
rect 137554 159712 137560 159724
rect 109736 159684 137560 159712
rect 109736 159672 109742 159684
rect 137554 159672 137560 159684
rect 137612 159672 137618 159724
rect 139946 159672 139952 159724
rect 140004 159712 140010 159724
rect 146956 159712 146984 159820
rect 147030 159808 147036 159860
rect 147088 159848 147094 159860
rect 150526 159848 150532 159860
rect 147088 159820 150532 159848
rect 147088 159808 147094 159820
rect 150526 159808 150532 159820
rect 150584 159808 150590 159860
rect 147306 159740 147312 159792
rect 147364 159780 147370 159792
rect 148870 159780 148876 159792
rect 147364 159752 148876 159780
rect 147364 159740 147370 159752
rect 148870 159740 148876 159752
rect 148928 159740 148934 159792
rect 150636 159780 150664 159888
rect 152458 159876 152464 159928
rect 152516 159916 152522 159928
rect 160094 159916 160100 159928
rect 152516 159888 160100 159916
rect 152516 159876 152522 159888
rect 160094 159876 160100 159888
rect 160152 159876 160158 159928
rect 160186 159876 160192 159928
rect 160244 159916 160250 159928
rect 188338 159916 188344 159928
rect 160244 159888 188344 159916
rect 160244 159876 160250 159888
rect 188338 159876 188344 159888
rect 188396 159876 188402 159928
rect 191282 159876 191288 159928
rect 191340 159916 191346 159928
rect 264882 159916 264888 159928
rect 191340 159888 264888 159916
rect 191340 159876 191346 159888
rect 264882 159876 264888 159888
rect 264940 159876 264946 159928
rect 268654 159876 268660 159928
rect 268712 159916 268718 159928
rect 324038 159916 324044 159928
rect 268712 159888 324044 159916
rect 268712 159876 268718 159888
rect 324038 159876 324044 159888
rect 324096 159876 324102 159928
rect 328362 159876 328368 159928
rect 328420 159916 328426 159928
rect 369486 159916 369492 159928
rect 328420 159888 369492 159916
rect 328420 159876 328426 159888
rect 369486 159876 369492 159888
rect 369544 159876 369550 159928
rect 372154 159876 372160 159928
rect 372212 159916 372218 159928
rect 396166 159916 396172 159928
rect 372212 159888 396172 159916
rect 372212 159876 372218 159888
rect 396166 159876 396172 159888
rect 396224 159876 396230 159928
rect 403250 159876 403256 159928
rect 403308 159916 403314 159928
rect 416590 159916 416596 159928
rect 403308 159888 416596 159916
rect 403308 159876 403314 159888
rect 416590 159876 416596 159888
rect 416648 159876 416654 159928
rect 450354 159876 450360 159928
rect 450412 159916 450418 159928
rect 457162 159916 457168 159928
rect 450412 159888 457168 159916
rect 450412 159876 450418 159888
rect 457162 159876 457168 159888
rect 457220 159876 457226 159928
rect 458726 159876 458732 159928
rect 458784 159916 458790 159928
rect 465074 159916 465080 159928
rect 458784 159888 465080 159916
rect 458784 159876 458790 159888
rect 465074 159876 465080 159888
rect 465132 159876 465138 159928
rect 478966 159876 478972 159928
rect 479024 159916 479030 159928
rect 484578 159916 484584 159928
rect 479024 159888 484584 159916
rect 479024 159876 479030 159888
rect 484578 159876 484584 159888
rect 484636 159876 484642 159928
rect 150710 159808 150716 159860
rect 150768 159848 150774 159860
rect 174630 159848 174636 159860
rect 150768 159820 174636 159848
rect 150768 159808 150774 159820
rect 174630 159808 174636 159820
rect 174688 159808 174694 159860
rect 180702 159848 180708 159860
rect 174740 159820 180708 159848
rect 153378 159780 153384 159792
rect 148980 159752 149284 159780
rect 150636 159752 153384 159780
rect 148980 159712 149008 159752
rect 140004 159684 146800 159712
rect 146956 159684 149008 159712
rect 140004 159672 140010 159684
rect 49970 159604 49976 159656
rect 50028 159644 50034 159656
rect 143258 159644 143264 159656
rect 50028 159616 143264 159644
rect 50028 159604 50034 159616
rect 143258 159604 143264 159616
rect 143316 159604 143322 159656
rect 143350 159604 143356 159656
rect 143408 159644 143414 159656
rect 146662 159644 146668 159656
rect 143408 159616 146668 159644
rect 143408 159604 143414 159616
rect 146662 159604 146668 159616
rect 146720 159604 146726 159656
rect 32306 159536 32312 159588
rect 32364 159576 32370 159588
rect 126422 159576 126428 159588
rect 32364 159548 126428 159576
rect 32364 159536 32370 159548
rect 126422 159536 126428 159548
rect 126480 159536 126486 159588
rect 126606 159536 126612 159588
rect 126664 159576 126670 159588
rect 146202 159576 146208 159588
rect 126664 159548 146208 159576
rect 126664 159536 126670 159548
rect 146202 159536 146208 159548
rect 146260 159536 146266 159588
rect 146772 159576 146800 159684
rect 146938 159604 146944 159656
rect 146996 159644 147002 159656
rect 149054 159644 149060 159656
rect 146996 159616 149060 159644
rect 146996 159604 147002 159616
rect 149054 159604 149060 159616
rect 149112 159604 149118 159656
rect 149256 159644 149284 159752
rect 153378 159740 153384 159752
rect 153436 159740 153442 159792
rect 153470 159740 153476 159792
rect 153528 159780 153534 159792
rect 174740 159780 174768 159820
rect 180702 159808 180708 159820
rect 180760 159808 180766 159860
rect 184566 159808 184572 159860
rect 184624 159848 184630 159860
rect 259822 159848 259828 159860
rect 184624 159820 259828 159848
rect 184624 159808 184630 159820
rect 259822 159808 259828 159820
rect 259880 159808 259886 159860
rect 261938 159808 261944 159860
rect 261996 159848 262002 159860
rect 318978 159848 318984 159860
rect 261996 159820 318984 159848
rect 261996 159808 262002 159820
rect 318978 159808 318984 159820
rect 319036 159808 319042 159860
rect 320818 159808 320824 159860
rect 320876 159848 320882 159860
rect 357526 159848 357532 159860
rect 320876 159820 357532 159848
rect 320876 159808 320882 159820
rect 357526 159808 357532 159820
rect 357584 159808 357590 159860
rect 357986 159848 357992 159860
rect 357636 159820 357992 159848
rect 153528 159752 174768 159780
rect 153528 159740 153534 159752
rect 177850 159740 177856 159792
rect 177908 159780 177914 159792
rect 253934 159780 253940 159792
rect 177908 159752 253940 159780
rect 177908 159740 177914 159752
rect 253934 159740 253940 159752
rect 253992 159740 253998 159792
rect 255222 159740 255228 159792
rect 255280 159780 255286 159792
rect 313734 159780 313740 159792
rect 255280 159752 313740 159780
rect 255280 159740 255286 159752
rect 313734 159740 313740 159752
rect 313792 159740 313798 159792
rect 314102 159740 314108 159792
rect 314160 159780 314166 159792
rect 357636 159780 357664 159820
rect 357986 159808 357992 159820
rect 358044 159808 358050 159860
rect 376294 159808 376300 159860
rect 376352 159848 376358 159860
rect 406194 159848 406200 159860
rect 376352 159820 406200 159848
rect 376352 159808 376358 159820
rect 406194 159808 406200 159820
rect 406252 159808 406258 159860
rect 467190 159808 467196 159860
rect 467248 159848 467254 159860
rect 473354 159848 473360 159860
rect 467248 159820 473360 159848
rect 467248 159808 467254 159820
rect 473354 159808 473360 159820
rect 473412 159808 473418 159860
rect 314160 159752 357664 159780
rect 314160 159740 314166 159752
rect 357802 159740 357808 159792
rect 357860 159780 357866 159792
rect 365346 159780 365352 159792
rect 357860 159752 365352 159780
rect 357860 159740 357866 159752
rect 365346 159740 365352 159752
rect 365404 159740 365410 159792
rect 365438 159740 365444 159792
rect 365496 159780 365502 159792
rect 395522 159780 395528 159792
rect 365496 159752 395528 159780
rect 365496 159740 365502 159752
rect 395522 159740 395528 159752
rect 395580 159740 395586 159792
rect 396534 159740 396540 159792
rect 396592 159780 396598 159792
rect 413646 159780 413652 159792
rect 396592 159752 413652 159780
rect 396592 159740 396598 159752
rect 413646 159740 413652 159752
rect 413704 159740 413710 159792
rect 424318 159740 424324 159792
rect 424376 159780 424382 159792
rect 442718 159780 442724 159792
rect 424376 159752 442724 159780
rect 424376 159740 424382 159752
rect 442718 159740 442724 159752
rect 442776 159740 442782 159792
rect 471422 159740 471428 159792
rect 471480 159780 471486 159792
rect 477678 159780 477684 159792
rect 471480 159752 477684 159780
rect 471480 159740 471486 159752
rect 477678 159740 477684 159752
rect 477736 159740 477742 159792
rect 149330 159672 149336 159724
rect 149388 159712 149394 159724
rect 164142 159712 164148 159724
rect 149388 159684 164148 159712
rect 149388 159672 149394 159684
rect 164142 159672 164148 159684
rect 164200 159672 164206 159724
rect 167730 159672 167736 159724
rect 167788 159712 167794 159724
rect 245838 159712 245844 159724
rect 167788 159684 245844 159712
rect 167788 159672 167794 159684
rect 245838 159672 245844 159684
rect 245896 159672 245902 159724
rect 248506 159672 248512 159724
rect 248564 159712 248570 159724
rect 248564 159684 306374 159712
rect 248564 159672 248570 159684
rect 160094 159644 160100 159656
rect 149256 159616 160100 159644
rect 160094 159604 160100 159616
rect 160152 159604 160158 159656
rect 161014 159604 161020 159656
rect 161072 159644 161078 159656
rect 240318 159644 240324 159656
rect 161072 159616 240324 159644
rect 161072 159604 161078 159616
rect 240318 159604 240324 159616
rect 240376 159604 240382 159656
rect 241790 159604 241796 159656
rect 241848 159644 241854 159656
rect 302418 159644 302424 159656
rect 241848 159616 302424 159644
rect 241848 159604 241854 159616
rect 302418 159604 302424 159616
rect 302476 159604 302482 159656
rect 306346 159644 306374 159684
rect 308214 159672 308220 159724
rect 308272 159712 308278 159724
rect 347682 159712 347688 159724
rect 308272 159684 347688 159712
rect 308272 159672 308278 159684
rect 347682 159672 347688 159684
rect 347740 159672 347746 159724
rect 347774 159672 347780 159724
rect 347832 159712 347838 159724
rect 378778 159712 378784 159724
rect 347832 159684 378784 159712
rect 347832 159672 347838 159684
rect 378778 159672 378784 159684
rect 378836 159672 378842 159724
rect 379698 159672 379704 159724
rect 379756 159712 379762 159724
rect 405826 159712 405832 159724
rect 379756 159684 405832 159712
rect 379756 159672 379762 159684
rect 405826 159672 405832 159684
rect 405884 159672 405890 159724
rect 409966 159672 409972 159724
rect 410024 159712 410030 159724
rect 417878 159712 417884 159724
rect 410024 159684 417884 159712
rect 410024 159672 410030 159684
rect 417878 159672 417884 159684
rect 417936 159672 417942 159724
rect 420914 159672 420920 159724
rect 420972 159712 420978 159724
rect 440326 159712 440332 159724
rect 420972 159684 440332 159712
rect 420972 159672 420978 159684
rect 440326 159672 440332 159684
rect 440384 159672 440390 159724
rect 308582 159644 308588 159656
rect 306346 159616 308588 159644
rect 308582 159604 308588 159616
rect 308640 159604 308646 159656
rect 309042 159604 309048 159656
rect 309100 159644 309106 159656
rect 354858 159644 354864 159656
rect 309100 159616 354864 159644
rect 309100 159604 309106 159616
rect 354858 159604 354864 159616
rect 354916 159604 354922 159656
rect 355226 159604 355232 159656
rect 355284 159644 355290 159656
rect 362954 159644 362960 159656
rect 355284 159616 362960 159644
rect 355284 159604 355290 159616
rect 362954 159604 362960 159616
rect 363012 159604 363018 159656
rect 369578 159604 369584 159656
rect 369636 159644 369642 159656
rect 401042 159644 401048 159656
rect 369636 159616 401048 159644
rect 369636 159604 369642 159616
rect 401042 159604 401048 159616
rect 401100 159604 401106 159656
rect 414198 159604 414204 159656
rect 414256 159644 414262 159656
rect 435082 159644 435088 159656
rect 414256 159616 435088 159644
rect 414256 159604 414262 159616
rect 435082 159604 435088 159616
rect 435140 159604 435146 159656
rect 459646 159604 459652 159656
rect 459704 159644 459710 159656
rect 466454 159644 466460 159656
rect 459704 159616 466460 159644
rect 459704 159604 459710 159616
rect 466454 159604 466460 159616
rect 466512 159604 466518 159656
rect 468018 159604 468024 159656
rect 468076 159644 468082 159656
rect 476022 159644 476028 159656
rect 468076 159616 476028 159644
rect 468076 159604 468082 159616
rect 476022 159604 476028 159616
rect 476080 159604 476086 159656
rect 157150 159576 157156 159588
rect 146772 159548 157156 159576
rect 157150 159536 157156 159548
rect 157208 159536 157214 159588
rect 157610 159536 157616 159588
rect 157668 159576 157674 159588
rect 239306 159576 239312 159588
rect 157668 159548 239312 159576
rect 157668 159536 157674 159548
rect 239306 159536 239312 159548
rect 239364 159536 239370 159588
rect 250990 159536 250996 159588
rect 251048 159576 251054 159588
rect 310606 159576 310612 159588
rect 251048 159548 310612 159576
rect 251048 159536 251054 159548
rect 310606 159536 310612 159548
rect 310664 159536 310670 159588
rect 315758 159536 315764 159588
rect 315816 159576 315822 159588
rect 358906 159576 358912 159588
rect 315816 159548 358912 159576
rect 315816 159536 315822 159548
rect 358906 159536 358912 159548
rect 358964 159536 358970 159588
rect 362862 159536 362868 159588
rect 362920 159576 362926 159588
rect 394786 159576 394792 159588
rect 362920 159548 394792 159576
rect 362920 159536 362926 159548
rect 394786 159536 394792 159548
rect 394844 159536 394850 159588
rect 399018 159536 399024 159588
rect 399076 159576 399082 159588
rect 408494 159576 408500 159588
rect 399076 159548 408500 159576
rect 399076 159536 399082 159548
rect 408494 159536 408500 159548
rect 408552 159536 408558 159588
rect 410794 159536 410800 159588
rect 410852 159576 410858 159588
rect 432506 159576 432512 159588
rect 410852 159548 432512 159576
rect 410852 159536 410858 159548
rect 432506 159536 432512 159548
rect 432564 159536 432570 159588
rect 448698 159536 448704 159588
rect 448756 159576 448762 159588
rect 456058 159576 456064 159588
rect 448756 159548 456064 159576
rect 448756 159536 448762 159548
rect 456058 159536 456064 159548
rect 456116 159536 456122 159588
rect 460474 159536 460480 159588
rect 460532 159576 460538 159588
rect 466638 159576 466644 159588
rect 460532 159548 466644 159576
rect 460532 159536 460538 159548
rect 466638 159536 466644 159548
rect 466696 159536 466702 159588
rect 470502 159536 470508 159588
rect 470560 159576 470566 159588
rect 476114 159576 476120 159588
rect 470560 159548 476120 159576
rect 470560 159536 470566 159548
rect 476114 159536 476120 159548
rect 476172 159536 476178 159588
rect 479794 159536 479800 159588
rect 479852 159576 479858 159588
rect 485222 159576 485228 159588
rect 479852 159548 485228 159576
rect 479852 159536 479858 159548
rect 485222 159536 485228 159548
rect 485280 159536 485286 159588
rect 43254 159468 43260 159520
rect 43312 159508 43318 159520
rect 137370 159508 137376 159520
rect 43312 159480 137376 159508
rect 43312 159468 43318 159480
rect 137370 159468 137376 159480
rect 137428 159468 137434 159520
rect 137462 159468 137468 159520
rect 137520 159508 137526 159520
rect 146754 159508 146760 159520
rect 137520 159480 146760 159508
rect 137520 159468 137526 159480
rect 146754 159468 146760 159480
rect 146812 159468 146818 159520
rect 225046 159508 225052 159520
rect 147048 159480 225052 159508
rect 36538 159400 36544 159452
rect 36596 159440 36602 159452
rect 135162 159440 135168 159452
rect 36596 159412 135168 159440
rect 36596 159400 36602 159412
rect 135162 159400 135168 159412
rect 135220 159400 135226 159452
rect 136542 159400 136548 159452
rect 136600 159440 136606 159452
rect 144086 159440 144092 159452
rect 136600 159412 144092 159440
rect 136600 159400 136606 159412
rect 144086 159400 144092 159412
rect 144144 159400 144150 159452
rect 144178 159400 144184 159452
rect 144236 159440 144242 159452
rect 147048 159440 147076 159480
rect 225046 159468 225052 159480
rect 225104 159468 225110 159520
rect 231670 159468 231676 159520
rect 231728 159508 231734 159520
rect 295518 159508 295524 159520
rect 231728 159480 295524 159508
rect 231728 159468 231734 159480
rect 295518 159468 295524 159480
rect 295576 159468 295582 159520
rect 295610 159468 295616 159520
rect 295668 159508 295674 159520
rect 339218 159508 339224 159520
rect 295668 159480 339224 159508
rect 295668 159468 295674 159480
rect 339218 159468 339224 159480
rect 339276 159468 339282 159520
rect 339310 159468 339316 159520
rect 339368 159508 339374 159520
rect 349798 159508 349804 159520
rect 339368 159480 349804 159508
rect 339368 159468 339374 159480
rect 349798 159468 349804 159480
rect 349856 159468 349862 159520
rect 354214 159508 354220 159520
rect 349908 159480 354220 159508
rect 144236 159412 147076 159440
rect 144236 159400 144242 159412
rect 147214 159400 147220 159452
rect 147272 159440 147278 159452
rect 150434 159440 150440 159452
rect 147272 159412 150440 159440
rect 147272 159400 147278 159412
rect 150434 159400 150440 159412
rect 150492 159400 150498 159452
rect 150894 159400 150900 159452
rect 150952 159440 150958 159452
rect 234154 159440 234160 159452
rect 150952 159412 234160 159440
rect 150952 159400 150958 159412
rect 234154 159400 234160 159412
rect 234212 159400 234218 159452
rect 234982 159400 234988 159452
rect 235040 159440 235046 159452
rect 298002 159440 298008 159452
rect 235040 159412 298008 159440
rect 235040 159400 235046 159412
rect 298002 159400 298008 159412
rect 298060 159400 298066 159452
rect 301498 159400 301504 159452
rect 301556 159440 301562 159452
rect 347958 159440 347964 159452
rect 301556 159412 347964 159440
rect 301556 159400 301562 159412
rect 347958 159400 347964 159412
rect 348016 159400 348022 159452
rect 348050 159400 348056 159452
rect 348108 159440 348114 159452
rect 349908 159440 349936 159480
rect 354214 159468 354220 159480
rect 354272 159468 354278 159520
rect 358630 159468 358636 159520
rect 358688 159508 358694 159520
rect 392762 159508 392768 159520
rect 358688 159480 392768 159508
rect 358688 159468 358694 159480
rect 392762 159468 392768 159480
rect 392820 159468 392826 159520
rect 407482 159468 407488 159520
rect 407540 159508 407546 159520
rect 429930 159508 429936 159520
rect 407540 159480 429936 159508
rect 407540 159468 407546 159480
rect 429930 159468 429936 159480
rect 429988 159468 429994 159520
rect 449526 159468 449532 159520
rect 449584 159508 449590 159520
rect 455782 159508 455788 159520
rect 449584 159480 455788 159508
rect 449584 159468 449590 159480
rect 455782 159468 455788 159480
rect 455840 159468 455846 159520
rect 457070 159468 457076 159520
rect 457128 159508 457134 159520
rect 464154 159508 464160 159520
rect 457128 159480 464160 159508
rect 457128 159468 457134 159480
rect 464154 159468 464160 159480
rect 464212 159468 464218 159520
rect 468846 159468 468852 159520
rect 468904 159508 468910 159520
rect 474826 159508 474832 159520
rect 468904 159480 474832 159508
rect 468904 159468 468910 159480
rect 474826 159468 474832 159480
rect 474884 159468 474890 159520
rect 477310 159468 477316 159520
rect 477368 159508 477374 159520
rect 483290 159508 483296 159520
rect 477368 159480 483296 159508
rect 477368 159468 477374 159480
rect 483290 159468 483296 159480
rect 483348 159468 483354 159520
rect 518066 159468 518072 159520
rect 518124 159508 518130 159520
rect 522666 159508 522672 159520
rect 518124 159480 522672 159508
rect 518124 159468 518130 159480
rect 522666 159468 522672 159480
rect 522724 159468 522730 159520
rect 348108 159412 349936 159440
rect 348108 159400 348114 159412
rect 351086 159400 351092 159452
rect 351144 159440 351150 159452
rect 355594 159440 355600 159452
rect 351144 159412 355600 159440
rect 351144 159400 351150 159412
rect 355594 159400 355600 159412
rect 355652 159400 355658 159452
rect 356146 159400 356152 159452
rect 356204 159440 356210 159452
rect 390830 159440 390836 159452
rect 356204 159412 390836 159440
rect 356204 159400 356210 159412
rect 390830 159400 390836 159412
rect 390888 159400 390894 159452
rect 427630 159400 427636 159452
rect 427688 159440 427694 159452
rect 445386 159440 445392 159452
rect 427688 159412 445392 159440
rect 427688 159400 427694 159412
rect 445386 159400 445392 159412
rect 445444 159400 445450 159452
rect 451182 159400 451188 159452
rect 451240 159440 451246 159452
rect 456794 159440 456800 159452
rect 451240 159412 456800 159440
rect 451240 159400 451246 159412
rect 456794 159400 456800 159412
rect 456852 159400 456858 159452
rect 6270 159332 6276 159384
rect 6328 159372 6334 159384
rect 122650 159372 122656 159384
rect 6328 159344 122656 159372
rect 6328 159332 6334 159344
rect 122650 159332 122656 159344
rect 122708 159332 122714 159384
rect 123110 159332 123116 159384
rect 123168 159372 123174 159384
rect 146846 159372 146852 159384
rect 123168 159344 146852 159372
rect 123168 159332 123174 159344
rect 146846 159332 146852 159344
rect 146904 159332 146910 159384
rect 146938 159332 146944 159384
rect 146996 159372 147002 159384
rect 223574 159372 223580 159384
rect 146996 159344 223580 159372
rect 146996 159332 147002 159344
rect 223574 159332 223580 159344
rect 223632 159332 223638 159384
rect 224954 159332 224960 159384
rect 225012 159372 225018 159384
rect 290642 159372 290648 159384
rect 225012 159344 290648 159372
rect 225012 159332 225018 159344
rect 290642 159332 290648 159344
rect 290700 159332 290706 159384
rect 294782 159332 294788 159384
rect 294840 159372 294846 159384
rect 294840 159344 338528 159372
rect 294840 159332 294846 159344
rect 76926 159264 76932 159316
rect 76984 159304 76990 159316
rect 152458 159304 152464 159316
rect 76984 159276 152464 159304
rect 76984 159264 76990 159276
rect 152458 159264 152464 159276
rect 152516 159264 152522 159316
rect 163498 159264 163504 159316
rect 163556 159304 163562 159316
rect 196986 159304 196992 159316
rect 163556 159276 196992 159304
rect 163556 159264 163562 159276
rect 196986 159264 196992 159276
rect 197044 159264 197050 159316
rect 201402 159264 201408 159316
rect 201460 159304 201466 159316
rect 212626 159304 212632 159316
rect 201460 159276 212632 159304
rect 201460 159264 201466 159276
rect 212626 159264 212632 159276
rect 212684 159264 212690 159316
rect 214006 159264 214012 159316
rect 214064 159304 214070 159316
rect 281534 159304 281540 159316
rect 214064 159276 281540 159304
rect 214064 159264 214070 159276
rect 281534 159264 281540 159276
rect 281592 159264 281598 159316
rect 282086 159264 282092 159316
rect 282144 159304 282150 159316
rect 327442 159304 327448 159316
rect 282144 159276 327448 159304
rect 282144 159264 282150 159276
rect 327442 159264 327448 159276
rect 327500 159264 327506 159316
rect 327534 159264 327540 159316
rect 327592 159304 327598 159316
rect 330570 159304 330576 159316
rect 327592 159276 330576 159304
rect 327592 159264 327598 159276
rect 330570 159264 330576 159276
rect 330628 159264 330634 159316
rect 330662 159264 330668 159316
rect 330720 159304 330726 159316
rect 333698 159304 333704 159316
rect 330720 159276 333704 159304
rect 330720 159264 330726 159276
rect 333698 159264 333704 159276
rect 333756 159264 333762 159316
rect 335354 159264 335360 159316
rect 335412 159304 335418 159316
rect 338298 159304 338304 159316
rect 335412 159276 338304 159304
rect 335412 159264 335418 159276
rect 338298 159264 338304 159276
rect 338356 159264 338362 159316
rect 93670 159196 93676 159248
rect 93728 159236 93734 159248
rect 93728 159208 171134 159236
rect 93728 159196 93734 159208
rect 86954 159128 86960 159180
rect 87012 159168 87018 159180
rect 169754 159168 169760 159180
rect 87012 159140 169760 159168
rect 87012 159128 87018 159140
rect 169754 159128 169760 159140
rect 169812 159128 169818 159180
rect 171106 159168 171134 159208
rect 180334 159196 180340 159248
rect 180392 159236 180398 159248
rect 183554 159236 183560 159248
rect 180392 159208 183560 159236
rect 180392 159196 180398 159208
rect 183554 159196 183560 159208
rect 183612 159196 183618 159248
rect 187050 159196 187056 159248
rect 187108 159236 187114 159248
rect 216674 159236 216680 159248
rect 187108 159208 216680 159236
rect 187108 159196 187114 159208
rect 216674 159196 216680 159208
rect 216732 159196 216738 159248
rect 218238 159196 218244 159248
rect 218296 159236 218302 159248
rect 285398 159236 285404 159248
rect 218296 159208 285404 159236
rect 218296 159196 218302 159208
rect 285398 159196 285404 159208
rect 285456 159196 285462 159248
rect 287974 159196 287980 159248
rect 288032 159236 288038 159248
rect 338390 159236 338396 159248
rect 288032 159208 338396 159236
rect 288032 159196 288038 159208
rect 338390 159196 338396 159208
rect 338448 159196 338454 159248
rect 338500 159236 338528 159344
rect 338666 159332 338672 159384
rect 338724 159372 338730 159384
rect 339494 159372 339500 159384
rect 338724 159344 339500 159372
rect 338724 159332 338730 159344
rect 339494 159332 339500 159344
rect 339552 159332 339558 159384
rect 339586 159332 339592 159384
rect 339644 159372 339650 159384
rect 342438 159372 342444 159384
rect 339644 159344 342444 159372
rect 339644 159332 339650 159344
rect 342438 159332 342444 159344
rect 342496 159332 342502 159384
rect 346026 159332 346032 159384
rect 346084 159372 346090 159384
rect 382826 159372 382832 159384
rect 346084 159344 382832 159372
rect 346084 159332 346090 159344
rect 382826 159332 382832 159344
rect 382884 159332 382890 159384
rect 392302 159332 392308 159384
rect 392360 159372 392366 159384
rect 403434 159372 403440 159384
rect 392360 159344 403440 159372
rect 392360 159332 392366 159344
rect 403434 159332 403440 159344
rect 403492 159332 403498 159384
rect 417510 159332 417516 159384
rect 417568 159372 417574 159384
rect 437658 159372 437664 159384
rect 417568 159344 437664 159372
rect 417568 159332 417574 159344
rect 437658 159332 437664 159344
rect 437716 159332 437722 159384
rect 447870 159332 447876 159384
rect 447928 159372 447934 159384
rect 447928 159344 451274 159372
rect 447928 159332 447934 159344
rect 338574 159264 338580 159316
rect 338632 159304 338638 159316
rect 374086 159304 374092 159316
rect 338632 159276 374092 159304
rect 338632 159264 338638 159276
rect 374086 159264 374092 159276
rect 374144 159264 374150 159316
rect 378042 159264 378048 159316
rect 378100 159304 378106 159316
rect 388346 159304 388352 159316
rect 378100 159276 388352 159304
rect 378100 159264 378106 159276
rect 388346 159264 388352 159276
rect 388404 159264 388410 159316
rect 388990 159264 388996 159316
rect 389048 159304 389054 159316
rect 403894 159304 403900 159316
rect 389048 159276 403900 159304
rect 389048 159264 389054 159276
rect 403894 159264 403900 159276
rect 403952 159264 403958 159316
rect 451246 159304 451274 159344
rect 453758 159332 453764 159384
rect 453816 159372 453822 159384
rect 459646 159372 459652 159384
rect 453816 159344 459652 159372
rect 453816 159332 453822 159344
rect 459646 159332 459652 159344
rect 459704 159332 459710 159384
rect 469674 159332 469680 159384
rect 469732 159372 469738 159384
rect 477402 159372 477408 159384
rect 469732 159344 477408 159372
rect 469732 159332 469738 159344
rect 477402 159332 477408 159344
rect 477460 159332 477466 159384
rect 478138 159332 478144 159384
rect 478196 159372 478202 159384
rect 483934 159372 483940 159384
rect 478196 159344 483940 159372
rect 478196 159332 478202 159344
rect 483934 159332 483940 159344
rect 483992 159332 483998 159384
rect 518710 159332 518716 159384
rect 518768 159372 518774 159384
rect 523494 159372 523500 159384
rect 518768 159344 523500 159372
rect 518768 159332 518774 159344
rect 523494 159332 523500 159344
rect 523552 159332 523558 159384
rect 456886 159304 456892 159316
rect 451246 159276 456892 159304
rect 456886 159264 456892 159276
rect 456944 159264 456950 159316
rect 457898 159264 457904 159316
rect 457956 159304 457962 159316
rect 464522 159304 464528 159316
rect 457956 159276 464528 159304
rect 457956 159264 457962 159276
rect 464522 159264 464528 159276
rect 464580 159264 464586 159316
rect 342346 159236 342352 159248
rect 338500 159208 342352 159236
rect 342346 159196 342352 159208
rect 342404 159196 342410 159248
rect 342714 159196 342720 159248
rect 342772 159236 342778 159248
rect 343818 159236 343824 159248
rect 342772 159208 343824 159236
rect 342772 159196 342778 159208
rect 343818 159196 343824 159208
rect 343876 159196 343882 159248
rect 349798 159196 349804 159248
rect 349856 159236 349862 159248
rect 377950 159236 377956 159248
rect 349856 159208 377956 159236
rect 349856 159196 349862 159208
rect 377950 159196 377956 159208
rect 378008 159196 378014 159248
rect 385586 159196 385592 159248
rect 385644 159236 385650 159248
rect 399846 159236 399852 159248
rect 385644 159208 399852 159236
rect 385644 159196 385650 159208
rect 399846 159196 399852 159208
rect 399904 159196 399910 159248
rect 461302 159196 461308 159248
rect 461360 159236 461366 159248
rect 468018 159236 468024 159248
rect 461360 159208 468024 159236
rect 461360 159196 461366 159208
rect 468018 159196 468024 159208
rect 468076 159196 468082 159248
rect 176654 159168 176660 159180
rect 171106 159140 176660 159168
rect 176654 159128 176660 159140
rect 176712 159128 176718 159180
rect 181438 159128 181444 159180
rect 181496 159168 181502 159180
rect 193122 159168 193128 159180
rect 181496 159140 183232 159168
rect 181496 159128 181502 159140
rect 100478 159060 100484 159112
rect 100536 159100 100542 159112
rect 183094 159100 183100 159112
rect 100536 159072 183100 159100
rect 100536 159060 100542 159072
rect 183094 159060 183100 159072
rect 183152 159060 183158 159112
rect 183204 159100 183232 159140
rect 183480 159140 193128 159168
rect 183480 159100 183508 159140
rect 193122 159128 193128 159140
rect 193180 159128 193186 159180
rect 193766 159128 193772 159180
rect 193824 159168 193830 159180
rect 220630 159168 220636 159180
rect 193824 159140 220636 159168
rect 193824 159128 193830 159140
rect 220630 159128 220636 159140
rect 220688 159128 220694 159180
rect 224126 159128 224132 159180
rect 224184 159168 224190 159180
rect 288342 159168 288348 159180
rect 224184 159140 288348 159168
rect 224184 159128 224190 159140
rect 288342 159128 288348 159140
rect 288400 159128 288406 159180
rect 288894 159128 288900 159180
rect 288952 159168 288958 159180
rect 339402 159168 339408 159180
rect 288952 159140 339408 159168
rect 288952 159128 288958 159140
rect 339402 159128 339408 159140
rect 339460 159128 339466 159180
rect 341886 159128 341892 159180
rect 341944 159168 341950 159180
rect 378226 159168 378232 159180
rect 341944 159140 378232 159168
rect 341944 159128 341950 159140
rect 378226 159128 378232 159140
rect 378284 159128 378290 159180
rect 395706 159128 395712 159180
rect 395764 159168 395770 159180
rect 405366 159168 405372 159180
rect 395764 159140 405372 159168
rect 395764 159128 395770 159140
rect 405366 159128 405372 159140
rect 405424 159128 405430 159180
rect 462130 159128 462136 159180
rect 462188 159168 462194 159180
rect 467926 159168 467932 159180
rect 462188 159140 467932 159168
rect 462188 159128 462194 159140
rect 467926 159128 467932 159140
rect 467984 159128 467990 159180
rect 183204 159072 183508 159100
rect 183738 159060 183744 159112
rect 183796 159100 183802 159112
rect 203794 159100 203800 159112
rect 183796 159072 203800 159100
rect 183796 159060 183802 159072
rect 203794 159060 203800 159072
rect 203852 159060 203858 159112
rect 203886 159060 203892 159112
rect 203944 159100 203950 159112
rect 210510 159100 210516 159112
rect 203944 159072 210516 159100
rect 203944 159060 203950 159072
rect 210510 159060 210516 159072
rect 210568 159060 210574 159112
rect 210602 159060 210608 159112
rect 210660 159100 210666 159112
rect 215294 159100 215300 159112
rect 210660 159072 215300 159100
rect 210660 159060 210666 159072
rect 215294 159060 215300 159072
rect 215352 159060 215358 159112
rect 220722 159060 220728 159112
rect 220780 159100 220786 159112
rect 278682 159100 278688 159112
rect 220780 159072 278688 159100
rect 220780 159060 220786 159072
rect 278682 159060 278688 159072
rect 278740 159060 278746 159112
rect 278774 159060 278780 159112
rect 278832 159100 278838 159112
rect 279878 159100 279884 159112
rect 278832 159072 279884 159100
rect 278832 159060 278838 159072
rect 279878 159060 279884 159072
rect 279936 159060 279942 159112
rect 280062 159060 280068 159112
rect 280120 159100 280126 159112
rect 282914 159100 282920 159112
rect 280120 159072 282920 159100
rect 280120 159060 280126 159072
rect 282914 159060 282920 159072
rect 282972 159060 282978 159112
rect 283006 159060 283012 159112
rect 283064 159100 283070 159112
rect 284202 159100 284208 159112
rect 283064 159072 284208 159100
rect 283064 159060 283070 159072
rect 284202 159060 284208 159072
rect 284260 159060 284266 159112
rect 284662 159060 284668 159112
rect 284720 159100 284726 159112
rect 285858 159100 285864 159112
rect 284720 159072 285864 159100
rect 284720 159060 284726 159072
rect 285858 159060 285864 159072
rect 285916 159060 285922 159112
rect 302326 159060 302332 159112
rect 302384 159100 302390 159112
rect 349706 159100 349712 159112
rect 302384 159072 349712 159100
rect 302384 159060 302390 159072
rect 349706 159060 349712 159072
rect 349764 159060 349770 159112
rect 351914 159060 351920 159112
rect 351972 159100 351978 159112
rect 385494 159100 385500 159112
rect 351972 159072 385500 159100
rect 351972 159060 351978 159072
rect 385494 159060 385500 159072
rect 385552 159060 385558 159112
rect 386414 159060 386420 159112
rect 386472 159100 386478 159112
rect 387702 159100 387708 159112
rect 386472 159072 387708 159100
rect 386472 159060 386478 159072
rect 387702 159060 387708 159072
rect 387760 159060 387766 159112
rect 412542 159060 412548 159112
rect 412600 159100 412606 159112
rect 413922 159100 413928 159112
rect 412600 159072 413928 159100
rect 412600 159060 412606 159072
rect 413922 159060 413928 159072
rect 413980 159060 413986 159112
rect 462958 159060 462964 159112
rect 463016 159100 463022 159112
rect 469214 159100 469220 159112
rect 463016 159072 469220 159100
rect 463016 159060 463022 159072
rect 469214 159060 469220 159072
rect 469272 159060 469278 159112
rect 472250 159060 472256 159112
rect 472308 159100 472314 159112
rect 479426 159100 479432 159112
rect 472308 159072 479432 159100
rect 472308 159060 472314 159072
rect 479426 159060 479432 159072
rect 479484 159060 479490 159112
rect 107194 158992 107200 159044
rect 107252 159032 107258 159044
rect 107252 159004 181576 159032
rect 107252 158992 107258 159004
rect 73522 158924 73528 158976
rect 73580 158964 73586 158976
rect 107562 158964 107568 158976
rect 73580 158936 107568 158964
rect 73580 158924 73586 158936
rect 107562 158924 107568 158936
rect 107620 158924 107626 158976
rect 119798 158924 119804 158976
rect 119856 158964 119862 158976
rect 126606 158964 126612 158976
rect 119856 158936 126612 158964
rect 119856 158924 119862 158936
rect 126606 158924 126612 158936
rect 126664 158924 126670 158976
rect 181438 158964 181444 158976
rect 126808 158936 181444 158964
rect 96246 158856 96252 158908
rect 96304 158896 96310 158908
rect 120534 158896 120540 158908
rect 96304 158868 120540 158896
rect 96304 158856 96310 158868
rect 120534 158856 120540 158868
rect 120592 158856 120598 158908
rect 120626 158856 120632 158908
rect 120684 158896 120690 158908
rect 121178 158896 121184 158908
rect 120684 158868 121184 158896
rect 120684 158856 120690 158868
rect 121178 158856 121184 158868
rect 121236 158856 121242 158908
rect 124030 158856 124036 158908
rect 124088 158896 124094 158908
rect 126808 158896 126836 158936
rect 181438 158924 181444 158936
rect 181496 158924 181502 158976
rect 181548 158964 181576 159004
rect 183646 158992 183652 159044
rect 183704 159032 183710 159044
rect 183704 159004 195284 159032
rect 183704 158992 183710 159004
rect 185578 158964 185584 158976
rect 181548 158936 185584 158964
rect 185578 158924 185584 158936
rect 185636 158924 185642 158976
rect 127802 158896 127808 158908
rect 124088 158868 126836 158896
rect 126900 158868 127808 158896
rect 124088 158856 124094 158868
rect 125502 158828 125508 158840
rect 103486 158800 125508 158828
rect 102962 158720 102968 158772
rect 103020 158760 103026 158772
rect 103486 158760 103514 158800
rect 125502 158788 125508 158800
rect 125560 158788 125566 158840
rect 126900 158828 126928 158868
rect 127802 158856 127808 158868
rect 127860 158856 127866 158908
rect 130746 158856 130752 158908
rect 130804 158896 130810 158908
rect 195146 158896 195152 158908
rect 130804 158868 195152 158896
rect 130804 158856 130810 158868
rect 195146 158856 195152 158868
rect 195204 158856 195210 158908
rect 195256 158896 195284 159004
rect 200086 159004 200620 159032
rect 197170 158924 197176 158976
rect 197228 158964 197234 158976
rect 200086 158964 200114 159004
rect 197228 158936 200114 158964
rect 200592 158964 200620 159004
rect 200666 158992 200672 159044
rect 200724 159032 200730 159044
rect 227714 159032 227720 159044
rect 200724 159004 227720 159032
rect 200724 158992 200730 159004
rect 227714 158992 227720 159004
rect 227772 158992 227778 159044
rect 230842 158992 230848 159044
rect 230900 159032 230906 159044
rect 295150 159032 295156 159044
rect 230900 159004 295156 159032
rect 230900 158992 230906 159004
rect 295150 158992 295156 159004
rect 295208 158992 295214 159044
rect 299474 159032 299480 159044
rect 296824 159004 299480 159032
rect 200592 158936 214604 158964
rect 197228 158924 197234 158936
rect 200390 158896 200396 158908
rect 195256 158868 200396 158896
rect 200390 158856 200396 158868
rect 200448 158856 200454 158908
rect 203794 158856 203800 158908
rect 203852 158896 203858 158908
rect 204898 158896 204904 158908
rect 203852 158868 204904 158896
rect 203852 158856 203858 158868
rect 204898 158856 204904 158868
rect 204956 158856 204962 158908
rect 210510 158856 210516 158908
rect 210568 158896 210574 158908
rect 213730 158896 213736 158908
rect 210568 158868 213736 158896
rect 210568 158856 210574 158868
rect 213730 158856 213736 158868
rect 213788 158856 213794 158908
rect 126440 158800 126928 158828
rect 103020 158732 103514 158760
rect 103020 158720 103026 158732
rect 106366 158720 106372 158772
rect 106424 158760 106430 158772
rect 126440 158760 126468 158800
rect 127342 158788 127348 158840
rect 127400 158828 127406 158840
rect 130838 158828 130844 158840
rect 127400 158800 130844 158828
rect 127400 158788 127406 158800
rect 130838 158788 130844 158800
rect 130896 158788 130902 158840
rect 133230 158788 133236 158840
rect 133288 158828 133294 158840
rect 133288 158800 137324 158828
rect 133288 158788 133294 158800
rect 106424 158732 126468 158760
rect 106424 158720 106430 158732
rect 126514 158720 126520 158772
rect 126572 158760 126578 158772
rect 137186 158760 137192 158772
rect 126572 158732 137192 158760
rect 126572 158720 126578 158732
rect 137186 158720 137192 158732
rect 137244 158720 137250 158772
rect 137296 158760 137324 158800
rect 137370 158788 137376 158840
rect 137428 158828 137434 158840
rect 147306 158828 147312 158840
rect 137428 158800 147312 158828
rect 137428 158788 137434 158800
rect 147306 158788 147312 158800
rect 147364 158788 147370 158840
rect 147582 158788 147588 158840
rect 147640 158828 147646 158840
rect 149054 158828 149060 158840
rect 147640 158800 149060 158828
rect 147640 158788 147646 158800
rect 149054 158788 149060 158800
rect 149112 158788 149118 158840
rect 149146 158788 149152 158840
rect 149204 158828 149210 158840
rect 156046 158828 156052 158840
rect 149204 158800 156052 158828
rect 149204 158788 149210 158800
rect 156046 158788 156052 158800
rect 156104 158788 156110 158840
rect 156782 158788 156788 158840
rect 156840 158828 156846 158840
rect 194502 158828 194508 158840
rect 156840 158800 194508 158828
rect 156840 158788 156846 158800
rect 194502 158788 194508 158800
rect 194560 158788 194566 158840
rect 194686 158788 194692 158840
rect 194744 158828 194750 158840
rect 203702 158828 203708 158840
rect 194744 158800 203708 158828
rect 194744 158788 194750 158800
rect 203702 158788 203708 158800
rect 203760 158788 203766 158840
rect 208118 158788 208124 158840
rect 208176 158828 208182 158840
rect 211982 158828 211988 158840
rect 208176 158800 211988 158828
rect 208176 158788 208182 158800
rect 211982 158788 211988 158800
rect 212040 158788 212046 158840
rect 214576 158828 214604 158936
rect 217318 158924 217324 158976
rect 217376 158964 217382 158976
rect 220446 158964 220452 158976
rect 217376 158936 220452 158964
rect 217376 158924 217382 158936
rect 220446 158924 220452 158936
rect 220504 158924 220510 158976
rect 238386 158924 238392 158976
rect 238444 158964 238450 158976
rect 242434 158964 242440 158976
rect 238444 158936 242440 158964
rect 238444 158924 238450 158936
rect 242434 158924 242440 158936
rect 242492 158924 242498 158976
rect 296824 158964 296852 159004
rect 299474 158992 299480 159004
rect 299532 158992 299538 159044
rect 307386 158992 307392 159044
rect 307444 159032 307450 159044
rect 353202 159032 353208 159044
rect 307444 159004 353208 159032
rect 307444 158992 307450 159004
rect 353202 158992 353208 159004
rect 353260 158992 353266 159044
rect 355594 158992 355600 159044
rect 355652 159032 355658 159044
rect 382550 159032 382556 159044
rect 355652 159004 382556 159032
rect 355652 158992 355658 159004
rect 382550 158992 382556 159004
rect 382608 158992 382614 159044
rect 383102 158992 383108 159044
rect 383160 159032 383166 159044
rect 411438 159032 411444 159044
rect 383160 159004 411444 159032
rect 383160 158992 383166 159004
rect 411438 158992 411444 159004
rect 411496 158992 411502 159044
rect 455414 158992 455420 159044
rect 455472 159032 455478 159044
rect 463326 159032 463332 159044
rect 455472 159004 463332 159032
rect 455472 158992 455478 159004
rect 463326 158992 463332 159004
rect 463384 158992 463390 159044
rect 473906 158992 473912 159044
rect 473964 159032 473970 159044
rect 480254 159032 480260 159044
rect 473964 159004 480260 159032
rect 473964 158992 473970 159004
rect 480254 158992 480260 159004
rect 480312 158992 480318 159044
rect 480622 158992 480628 159044
rect 480680 159032 480686 159044
rect 485866 159032 485872 159044
rect 480680 159004 485872 159032
rect 480680 158992 480686 159004
rect 485866 158992 485872 159004
rect 485924 158992 485930 159044
rect 507118 158992 507124 159044
rect 507176 159032 507182 159044
rect 508406 159032 508412 159044
rect 507176 159004 508412 159032
rect 507176 158992 507182 159004
rect 508406 158992 508412 159004
rect 508464 158992 508470 159044
rect 305362 158964 305368 158976
rect 248386 158936 296852 158964
rect 298020 158936 305368 158964
rect 214742 158856 214748 158908
rect 214800 158896 214806 158908
rect 248386 158896 248414 158936
rect 298020 158896 298048 158936
rect 305362 158924 305368 158936
rect 305420 158924 305426 158976
rect 310698 158924 310704 158976
rect 310756 158964 310762 158976
rect 313182 158964 313188 158976
rect 310756 158936 313188 158964
rect 310756 158924 310762 158936
rect 313182 158924 313188 158936
rect 313240 158924 313246 158976
rect 314930 158924 314936 158976
rect 314988 158964 314994 158976
rect 357434 158964 357440 158976
rect 314988 158936 357440 158964
rect 314988 158924 314994 158936
rect 357434 158924 357440 158936
rect 357492 158924 357498 158976
rect 357526 158924 357532 158976
rect 357584 158964 357590 158976
rect 363506 158964 363512 158976
rect 357584 158936 363512 158964
rect 357584 158924 357590 158936
rect 363506 158924 363512 158936
rect 363564 158924 363570 158976
rect 365162 158964 365168 158976
rect 364306 158936 365168 158964
rect 214800 158868 229094 158896
rect 214800 158856 214806 158868
rect 214576 158800 214788 158828
rect 158714 158760 158720 158772
rect 137296 158732 158720 158760
rect 158714 158720 158720 158732
rect 158772 158720 158778 158772
rect 171134 158720 171140 158772
rect 171192 158760 171198 158772
rect 172606 158760 172612 158772
rect 171192 158732 172612 158760
rect 171192 158720 171198 158732
rect 172606 158720 172612 158732
rect 172664 158720 172670 158772
rect 173618 158720 173624 158772
rect 173676 158760 173682 158772
rect 197354 158760 197360 158772
rect 173676 158732 197360 158760
rect 173676 158720 173682 158732
rect 197354 158720 197360 158732
rect 197412 158720 197418 158772
rect 207290 158720 207296 158772
rect 207348 158760 207354 158772
rect 214558 158760 214564 158772
rect 207348 158732 214564 158760
rect 207348 158720 207354 158732
rect 214558 158720 214564 158732
rect 214616 158720 214622 158772
rect 214760 158760 214788 158800
rect 214834 158788 214840 158840
rect 214892 158828 214898 158840
rect 221458 158828 221464 158840
rect 214892 158800 221464 158828
rect 214892 158788 214898 158800
rect 221458 158788 221464 158800
rect 221516 158788 221522 158840
rect 221550 158788 221556 158840
rect 221608 158828 221614 158840
rect 224770 158828 224776 158840
rect 221608 158800 224776 158828
rect 221608 158788 221614 158800
rect 224770 158788 224776 158800
rect 224828 158788 224834 158840
rect 229066 158828 229094 158868
rect 238726 158868 248414 158896
rect 258046 158868 298048 158896
rect 231302 158828 231308 158840
rect 229066 158800 231308 158828
rect 231302 158788 231308 158800
rect 231360 158788 231366 158840
rect 237558 158788 237564 158840
rect 237616 158828 237622 158840
rect 238726 158828 238754 158868
rect 237616 158800 238754 158828
rect 237616 158788 237622 158800
rect 244274 158788 244280 158840
rect 244332 158828 244338 158840
rect 258046 158828 258074 158868
rect 298094 158856 298100 158908
rect 298152 158896 298158 158908
rect 300302 158896 300308 158908
rect 298152 158868 300308 158896
rect 298152 158856 298158 158868
rect 300302 158856 300308 158868
rect 300360 158856 300366 158908
rect 305638 158856 305644 158908
rect 305696 158896 305702 158908
rect 307294 158896 307300 158908
rect 305696 158868 307300 158896
rect 305696 158856 305702 158868
rect 307294 158856 307300 158868
rect 307352 158856 307358 158908
rect 312446 158856 312452 158908
rect 312504 158896 312510 158908
rect 313458 158896 313464 158908
rect 312504 158868 313464 158896
rect 312504 158856 312510 158868
rect 313458 158856 313464 158868
rect 313516 158856 313522 158908
rect 364306 158896 364334 158936
rect 365162 158924 365168 158936
rect 365220 158924 365226 158976
rect 365346 158924 365352 158976
rect 365404 158964 365410 158976
rect 365404 158936 373994 158964
rect 365404 158924 365410 158936
rect 329668 158868 364334 158896
rect 373966 158896 373994 158936
rect 378686 158924 378692 158976
rect 378744 158964 378750 158976
rect 386230 158964 386236 158976
rect 378744 158936 386236 158964
rect 378744 158924 378750 158936
rect 386230 158924 386236 158936
rect 386288 158924 386294 158976
rect 391474 158924 391480 158976
rect 391532 158964 391538 158976
rect 394326 158964 394332 158976
rect 391532 158936 394332 158964
rect 391532 158924 391538 158936
rect 394326 158924 394332 158936
rect 394384 158924 394390 158976
rect 409138 158924 409144 158976
rect 409196 158964 409202 158976
rect 410886 158964 410892 158976
rect 409196 158936 410892 158964
rect 409196 158924 409202 158936
rect 410886 158924 410892 158936
rect 410944 158924 410950 158976
rect 416682 158924 416688 158976
rect 416740 158964 416746 158976
rect 419534 158964 419540 158976
rect 416740 158936 419540 158964
rect 416740 158924 416746 158936
rect 419534 158924 419540 158936
rect 419592 158924 419598 158976
rect 420086 158924 420092 158976
rect 420144 158964 420150 158976
rect 423582 158964 423588 158976
rect 420144 158936 423588 158964
rect 420144 158924 420150 158936
rect 423582 158924 423588 158936
rect 423640 158924 423646 158976
rect 454586 158924 454592 158976
rect 454644 158964 454650 158976
rect 461854 158964 461860 158976
rect 454644 158936 461860 158964
rect 454644 158924 454650 158936
rect 461854 158924 461860 158936
rect 461912 158924 461918 158976
rect 466362 158924 466368 158976
rect 466420 158964 466426 158976
rect 472526 158964 472532 158976
rect 466420 158936 472532 158964
rect 466420 158924 466426 158936
rect 472526 158924 472532 158936
rect 472584 158924 472590 158976
rect 475562 158924 475568 158976
rect 475620 158964 475626 158976
rect 482002 158964 482008 158976
rect 475620 158936 482008 158964
rect 475620 158924 475626 158936
rect 482002 158924 482008 158936
rect 482060 158924 482066 158976
rect 373966 158868 383654 158896
rect 244332 158800 258074 158828
rect 244332 158788 244338 158800
rect 261110 158788 261116 158840
rect 261168 158828 261174 158840
rect 317138 158828 317144 158840
rect 261168 158800 317144 158828
rect 261168 158788 261174 158800
rect 317138 158788 317144 158800
rect 317196 158788 317202 158840
rect 317414 158788 317420 158840
rect 317472 158828 317478 158840
rect 318426 158828 318432 158840
rect 317472 158800 318432 158828
rect 317472 158788 317478 158800
rect 318426 158788 318432 158800
rect 318484 158788 318490 158840
rect 319162 158788 319168 158840
rect 319220 158828 319226 158840
rect 321554 158828 321560 158840
rect 319220 158800 321560 158828
rect 319220 158788 319226 158800
rect 321554 158788 321560 158800
rect 321612 158788 321618 158840
rect 322474 158788 322480 158840
rect 322532 158828 322538 158840
rect 329668 158828 329696 158868
rect 355226 158828 355232 158840
rect 322532 158800 329696 158828
rect 330496 158800 355232 158828
rect 322532 158788 322538 158800
rect 222102 158760 222108 158772
rect 214760 158732 222108 158760
rect 222102 158720 222108 158732
rect 222160 158720 222166 158772
rect 240870 158720 240876 158772
rect 240928 158760 240934 158772
rect 243354 158760 243360 158772
rect 240928 158732 243360 158760
rect 240928 158720 240934 158732
rect 243354 158720 243360 158732
rect 243412 158720 243418 158772
rect 254394 158720 254400 158772
rect 254452 158760 254458 158772
rect 255406 158760 255412 158772
rect 254452 158732 255412 158760
rect 254452 158720 254458 158732
rect 255406 158720 255412 158732
rect 255464 158720 255470 158772
rect 258534 158720 258540 158772
rect 258592 158760 258598 158772
rect 261018 158760 261024 158772
rect 258592 158732 261024 158760
rect 258592 158720 258598 158732
rect 261018 158720 261024 158732
rect 261076 158720 261082 158772
rect 264422 158720 264428 158772
rect 264480 158760 264486 158772
rect 267642 158760 267648 158772
rect 264480 158732 267648 158760
rect 264480 158720 264486 158732
rect 267642 158720 267648 158732
rect 267700 158720 267706 158772
rect 267826 158720 267832 158772
rect 267884 158760 267890 158772
rect 320266 158760 320272 158772
rect 267884 158732 320272 158760
rect 267884 158720 267890 158732
rect 320266 158720 320272 158732
rect 320324 158720 320330 158772
rect 321646 158720 321652 158772
rect 321704 158760 321710 158772
rect 330496 158760 330524 158800
rect 355226 158788 355232 158800
rect 355284 158788 355290 158840
rect 360166 158800 361252 158828
rect 321704 158732 330524 158760
rect 321704 158720 321710 158732
rect 330570 158720 330576 158772
rect 330628 158760 330634 158772
rect 360166 158760 360194 158800
rect 330628 158732 360194 158760
rect 361224 158760 361252 158800
rect 361298 158788 361304 158840
rect 361356 158828 361362 158840
rect 383626 158828 383654 158868
rect 384758 158856 384764 158908
rect 384816 158896 384822 158908
rect 389634 158896 389640 158908
rect 384816 158868 389640 158896
rect 384816 158856 384822 158868
rect 389634 158856 389640 158868
rect 389692 158856 389698 158908
rect 446122 158856 446128 158908
rect 446180 158896 446186 158908
rect 453942 158896 453948 158908
rect 446180 158868 453948 158896
rect 446180 158856 446186 158868
rect 453942 158856 453948 158868
rect 454000 158856 454006 158908
rect 456242 158856 456248 158908
rect 456300 158896 456306 158908
rect 462958 158896 462964 158908
rect 456300 158868 462964 158896
rect 456300 158856 456306 158868
rect 462958 158856 462964 158868
rect 463016 158856 463022 158908
rect 463786 158856 463792 158908
rect 463844 158896 463850 158908
rect 471238 158896 471244 158908
rect 463844 158868 471244 158896
rect 463844 158856 463850 158868
rect 471238 158856 471244 158868
rect 471296 158856 471302 158908
rect 474734 158856 474740 158908
rect 474792 158896 474798 158908
rect 481358 158896 481364 158908
rect 474792 158868 481364 158896
rect 474792 158856 474798 158868
rect 481358 158856 481364 158868
rect 481416 158856 481422 158908
rect 481450 158856 481456 158908
rect 481508 158896 481514 158908
rect 486418 158896 486424 158908
rect 481508 158868 486424 158896
rect 481508 158856 481514 158868
rect 486418 158856 486424 158868
rect 486476 158856 486482 158908
rect 508406 158856 508412 158908
rect 508464 158896 508470 158908
rect 510062 158896 510068 158908
rect 508464 158868 510068 158896
rect 508464 158856 508470 158868
rect 510062 158856 510068 158868
rect 510120 158856 510126 158908
rect 384942 158828 384948 158840
rect 361356 158800 378824 158828
rect 383626 158800 384948 158828
rect 361356 158788 361362 158800
rect 367186 158760 367192 158772
rect 361224 158732 367192 158760
rect 330628 158720 330634 158732
rect 367186 158720 367192 158732
rect 367244 158720 367250 158772
rect 367922 158720 367928 158772
rect 367980 158760 367986 158772
rect 378686 158760 378692 158772
rect 367980 158732 378692 158760
rect 367980 158720 367986 158732
rect 378686 158720 378692 158732
rect 378744 158720 378750 158772
rect 378796 158760 378824 158800
rect 384942 158788 384948 158800
rect 385000 158788 385006 158840
rect 404906 158788 404912 158840
rect 404964 158828 404970 158840
rect 405642 158828 405648 158840
rect 404964 158800 405648 158828
rect 404964 158788 404970 158800
rect 405642 158788 405648 158800
rect 405700 158788 405706 158840
rect 452010 158788 452016 158840
rect 452068 158828 452074 158840
rect 458174 158828 458180 158840
rect 452068 158800 458180 158828
rect 452068 158788 452074 158800
rect 458174 158788 458180 158800
rect 458232 158788 458238 158840
rect 464614 158788 464620 158840
rect 464672 158828 464678 158840
rect 471606 158828 471612 158840
rect 464672 158800 471612 158828
rect 464672 158788 464678 158800
rect 471606 158788 471612 158800
rect 471664 158788 471670 158840
rect 476390 158788 476396 158840
rect 476448 158828 476454 158840
rect 481634 158828 481640 158840
rect 476448 158800 481640 158828
rect 476448 158788 476454 158800
rect 481634 158788 481640 158800
rect 481692 158788 481698 158840
rect 499942 158788 499948 158840
rect 500000 158828 500006 158840
rect 500586 158828 500592 158840
rect 500000 158800 500592 158828
rect 500000 158788 500006 158800
rect 500586 158788 500592 158800
rect 500644 158788 500650 158840
rect 506290 158788 506296 158840
rect 506348 158828 506354 158840
rect 507578 158828 507584 158840
rect 506348 158800 507584 158828
rect 506348 158788 506354 158800
rect 507578 158788 507584 158800
rect 507636 158788 507642 158840
rect 385310 158760 385316 158772
rect 378796 158732 385316 158760
rect 385310 158720 385316 158732
rect 385368 158720 385374 158772
rect 388070 158720 388076 158772
rect 388128 158760 388134 158772
rect 390370 158760 390376 158772
rect 388128 158732 390376 158760
rect 388128 158720 388134 158732
rect 390370 158720 390376 158732
rect 390428 158720 390434 158772
rect 405734 158720 405740 158772
rect 405792 158760 405798 158772
rect 409138 158760 409144 158772
rect 405792 158732 409144 158760
rect 405792 158720 405798 158732
rect 409138 158720 409144 158732
rect 409196 158720 409202 158772
rect 413370 158720 413376 158772
rect 413428 158760 413434 158772
rect 419626 158760 419632 158772
rect 413428 158732 419632 158760
rect 413428 158720 413434 158732
rect 419626 158720 419632 158732
rect 419684 158720 419690 158772
rect 435174 158720 435180 158772
rect 435232 158760 435238 158772
rect 435818 158760 435824 158772
rect 435232 158732 435824 158760
rect 435232 158720 435238 158732
rect 435818 158720 435824 158732
rect 435876 158720 435882 158772
rect 452838 158720 452844 158772
rect 452896 158760 452902 158772
rect 459554 158760 459560 158772
rect 452896 158732 459560 158760
rect 452896 158720 452902 158732
rect 459554 158720 459560 158732
rect 459612 158720 459618 158772
rect 465534 158720 465540 158772
rect 465592 158760 465598 158772
rect 472434 158760 472440 158772
rect 465592 158732 472440 158760
rect 465592 158720 465598 158732
rect 472434 158720 472440 158732
rect 472492 158720 472498 158772
rect 473078 158720 473084 158772
rect 473136 158760 473142 158772
rect 478966 158760 478972 158772
rect 473136 158732 478972 158760
rect 473136 158720 473142 158732
rect 478966 158720 478972 158732
rect 479024 158720 479030 158772
rect 482278 158720 482284 158772
rect 482336 158760 482342 158772
rect 487246 158760 487252 158772
rect 482336 158732 487252 158760
rect 482336 158720 482342 158732
rect 487246 158720 487252 158732
rect 487304 158720 487310 158772
rect 504450 158720 504456 158772
rect 504508 158760 504514 158772
rect 505002 158760 505008 158772
rect 504508 158732 505008 158760
rect 504508 158720 504514 158732
rect 505002 158720 505008 158732
rect 505060 158720 505066 158772
rect 505830 158720 505836 158772
rect 505888 158760 505894 158772
rect 506474 158760 506480 158772
rect 505888 158732 506480 158760
rect 505888 158720 505894 158732
rect 506474 158720 506480 158732
rect 506532 158720 506538 158772
rect 509694 158720 509700 158772
rect 509752 158760 509758 158772
rect 511718 158760 511724 158772
rect 509752 158732 511724 158760
rect 509752 158720 509758 158732
rect 511718 158720 511724 158732
rect 511776 158720 511782 158772
rect 514938 158720 514944 158772
rect 514996 158760 515002 158772
rect 518526 158760 518532 158772
rect 514996 158732 518532 158760
rect 514996 158720 515002 158732
rect 518526 158720 518532 158732
rect 518584 158720 518590 158772
rect 81066 158652 81072 158704
rect 81124 158692 81130 158704
rect 180794 158692 180800 158704
rect 81124 158664 180800 158692
rect 81124 158652 81130 158664
rect 180794 158652 180800 158664
rect 180852 158652 180858 158704
rect 180886 158652 180892 158704
rect 180944 158692 180950 158704
rect 181898 158692 181904 158704
rect 180944 158664 181904 158692
rect 180944 158652 180950 158664
rect 181898 158652 181904 158664
rect 181956 158652 181962 158704
rect 181990 158652 181996 158704
rect 182048 158692 182054 158704
rect 256786 158692 256792 158704
rect 182048 158664 256792 158692
rect 182048 158652 182054 158664
rect 256786 158652 256792 158664
rect 256844 158652 256850 158704
rect 67634 158584 67640 158636
rect 67692 158624 67698 158636
rect 170306 158624 170312 158636
rect 67692 158596 170312 158624
rect 67692 158584 67698 158596
rect 170306 158584 170312 158596
rect 170364 158584 170370 158636
rect 171962 158584 171968 158636
rect 172020 158624 172026 158636
rect 250070 158624 250076 158636
rect 172020 158596 250076 158624
rect 172020 158584 172026 158596
rect 250070 158584 250076 158596
rect 250128 158584 250134 158636
rect 71038 158516 71044 158568
rect 71096 158556 71102 158568
rect 172698 158556 172704 158568
rect 71096 158528 172704 158556
rect 71096 158516 71102 158528
rect 172698 158516 172704 158528
rect 172756 158516 172762 158568
rect 178678 158516 178684 158568
rect 178736 158556 178742 158568
rect 255314 158556 255320 158568
rect 178736 158528 255320 158556
rect 178736 158516 178742 158528
rect 255314 158516 255320 158528
rect 255372 158516 255378 158568
rect 74350 158448 74356 158500
rect 74408 158488 74414 158500
rect 175182 158488 175188 158500
rect 74408 158460 175188 158488
rect 74408 158448 74414 158460
rect 175182 158448 175188 158460
rect 175240 158448 175246 158500
rect 175274 158448 175280 158500
rect 175332 158488 175338 158500
rect 252554 158488 252560 158500
rect 175332 158460 252560 158488
rect 175332 158448 175338 158460
rect 252554 158448 252560 158460
rect 252612 158448 252618 158500
rect 64230 158380 64236 158432
rect 64288 158420 64294 158432
rect 167546 158420 167552 158432
rect 64288 158392 167552 158420
rect 64288 158380 64294 158392
rect 167546 158380 167552 158392
rect 167604 158380 167610 158432
rect 168558 158380 168564 158432
rect 168616 158420 168622 158432
rect 247586 158420 247592 158432
rect 168616 158392 247592 158420
rect 168616 158380 168622 158392
rect 247586 158380 247592 158392
rect 247644 158380 247650 158432
rect 60918 158312 60924 158364
rect 60976 158352 60982 158364
rect 164326 158352 164332 158364
rect 60976 158324 164332 158352
rect 60976 158312 60982 158324
rect 164326 158312 164332 158324
rect 164384 158312 164390 158364
rect 165246 158312 165252 158364
rect 165304 158352 165310 158364
rect 245010 158352 245016 158364
rect 165304 158324 245016 158352
rect 165304 158312 165310 158324
rect 245010 158312 245016 158324
rect 245068 158312 245074 158364
rect 54202 158244 54208 158296
rect 54260 158284 54266 158296
rect 160278 158284 160284 158296
rect 54260 158256 160284 158284
rect 54260 158244 54266 158256
rect 160278 158244 160284 158256
rect 160336 158244 160342 158296
rect 161842 158244 161848 158296
rect 161900 158284 161906 158296
rect 242066 158284 242072 158296
rect 161900 158256 242072 158284
rect 161900 158244 161906 158256
rect 242066 158244 242072 158256
rect 242124 158244 242130 158296
rect 50798 158176 50804 158228
rect 50856 158216 50862 158228
rect 157702 158216 157708 158228
rect 50856 158188 157708 158216
rect 50856 158176 50862 158188
rect 157702 158176 157708 158188
rect 157760 158176 157766 158228
rect 158438 158176 158444 158228
rect 158496 158216 158502 158228
rect 238846 158216 238852 158228
rect 158496 158188 238852 158216
rect 158496 158176 158502 158188
rect 238846 158176 238852 158188
rect 238904 158176 238910 158228
rect 256878 158176 256884 158228
rect 256936 158216 256942 158228
rect 315022 158216 315028 158228
rect 256936 158188 315028 158216
rect 256936 158176 256942 158188
rect 315022 158176 315028 158188
rect 315080 158176 315086 158228
rect 47486 158108 47492 158160
rect 47544 158148 47550 158160
rect 155034 158148 155040 158160
rect 47544 158120 155040 158148
rect 47544 158108 47550 158120
rect 155034 158108 155040 158120
rect 155092 158108 155098 158160
rect 155126 158108 155132 158160
rect 155184 158148 155190 158160
rect 237374 158148 237380 158160
rect 155184 158120 237380 158148
rect 155184 158108 155190 158120
rect 237374 158108 237380 158120
rect 237432 158108 237438 158160
rect 246758 158108 246764 158160
rect 246816 158148 246822 158160
rect 306926 158148 306932 158160
rect 246816 158120 306932 158148
rect 246816 158108 246822 158120
rect 306926 158108 306932 158120
rect 306984 158108 306990 158160
rect 37366 158040 37372 158092
rect 37424 158080 37430 158092
rect 146386 158080 146392 158092
rect 37424 158052 146392 158080
rect 37424 158040 37430 158052
rect 146386 158040 146392 158052
rect 146444 158040 146450 158092
rect 148410 158040 148416 158092
rect 148468 158080 148474 158092
rect 231854 158080 231860 158092
rect 148468 158052 231860 158080
rect 148468 158040 148474 158052
rect 231854 158040 231860 158052
rect 231912 158040 231918 158092
rect 233326 158040 233332 158092
rect 233384 158080 233390 158092
rect 297082 158080 297088 158092
rect 233384 158052 297088 158080
rect 233384 158040 233390 158052
rect 297082 158040 297088 158052
rect 297140 158040 297146 158092
rect 300670 158040 300676 158092
rect 300728 158080 300734 158092
rect 348418 158080 348424 158092
rect 300728 158052 348424 158080
rect 300728 158040 300734 158052
rect 348418 158040 348424 158052
rect 348476 158040 348482 158092
rect 382 157972 388 158024
rect 440 158012 446 158024
rect 118878 158012 118884 158024
rect 440 157984 118884 158012
rect 440 157972 446 157984
rect 118878 157972 118884 157984
rect 118936 157972 118942 158024
rect 131574 157972 131580 158024
rect 131632 158012 131638 158024
rect 218238 158012 218244 158024
rect 131632 157984 218244 158012
rect 131632 157972 131638 157984
rect 218238 157972 218244 157984
rect 218296 157972 218302 158024
rect 240042 157972 240048 158024
rect 240100 158012 240106 158024
rect 302234 158012 302240 158024
rect 240100 157984 302240 158012
rect 240100 157972 240106 157984
rect 302234 157972 302240 157984
rect 302292 157972 302298 158024
rect 77754 157904 77760 157956
rect 77812 157944 77818 157956
rect 77812 157916 176056 157944
rect 77812 157904 77818 157916
rect 84470 157836 84476 157888
rect 84528 157876 84534 157888
rect 175918 157876 175924 157888
rect 84528 157848 175924 157876
rect 84528 157836 84534 157848
rect 175918 157836 175924 157848
rect 175976 157836 175982 157888
rect 176028 157876 176056 157916
rect 176194 157904 176200 157956
rect 176252 157944 176258 157956
rect 182266 157944 182272 157956
rect 176252 157916 182272 157944
rect 176252 157904 176258 157916
rect 182266 157904 182272 157916
rect 182324 157904 182330 157956
rect 185394 157904 185400 157956
rect 185452 157944 185458 157956
rect 259454 157944 259460 157956
rect 185452 157916 259460 157944
rect 185452 157904 185458 157916
rect 259454 157904 259460 157916
rect 259512 157904 259518 157956
rect 178034 157876 178040 157888
rect 176028 157848 178040 157876
rect 178034 157836 178040 157848
rect 178092 157836 178098 157888
rect 181530 157836 181536 157888
rect 181588 157876 181594 157888
rect 188522 157876 188528 157888
rect 181588 157848 188528 157876
rect 181588 157836 181594 157848
rect 188522 157836 188528 157848
rect 188580 157836 188586 157888
rect 188798 157836 188804 157888
rect 188856 157876 188862 157888
rect 263042 157876 263048 157888
rect 188856 157848 263048 157876
rect 188856 157836 188862 157848
rect 263042 157836 263048 157848
rect 263100 157836 263106 157888
rect 87782 157768 87788 157820
rect 87840 157808 87846 157820
rect 181622 157808 181628 157820
rect 87840 157780 181628 157808
rect 87840 157768 87846 157780
rect 181622 157768 181628 157780
rect 181680 157768 181686 157820
rect 181806 157768 181812 157820
rect 181864 157808 181870 157820
rect 190638 157808 190644 157820
rect 181864 157780 190644 157808
rect 181864 157768 181870 157780
rect 190638 157768 190644 157780
rect 190696 157768 190702 157820
rect 195514 157768 195520 157820
rect 195572 157808 195578 157820
rect 267734 157808 267740 157820
rect 195572 157780 267740 157808
rect 195572 157768 195578 157780
rect 267734 157768 267740 157780
rect 267792 157768 267798 157820
rect 91186 157700 91192 157752
rect 91244 157740 91250 157752
rect 181254 157740 181260 157752
rect 91244 157712 181260 157740
rect 91244 157700 91250 157712
rect 181254 157700 181260 157712
rect 181312 157700 181318 157752
rect 181898 157700 181904 157752
rect 181956 157740 181962 157752
rect 181956 157712 186314 157740
rect 181956 157700 181962 157712
rect 94590 157632 94596 157684
rect 94648 157672 94654 157684
rect 181530 157672 181536 157684
rect 94648 157644 181536 157672
rect 94648 157632 94654 157644
rect 181530 157632 181536 157644
rect 181588 157632 181594 157684
rect 181714 157632 181720 157684
rect 181772 157672 181778 157684
rect 185394 157672 185400 157684
rect 181772 157644 185400 157672
rect 181772 157632 181778 157644
rect 185394 157632 185400 157644
rect 185452 157632 185458 157684
rect 186286 157672 186314 157712
rect 190454 157700 190460 157752
rect 190512 157740 190518 157752
rect 263778 157740 263784 157752
rect 190512 157712 263784 157740
rect 190512 157700 190518 157712
rect 263778 157700 263784 157712
rect 263836 157700 263842 157752
rect 236086 157672 236092 157684
rect 186286 157644 236092 157672
rect 236086 157632 236092 157644
rect 236144 157632 236150 157684
rect 97902 157564 97908 157616
rect 97960 157604 97966 157616
rect 193214 157604 193220 157616
rect 97960 157576 193220 157604
rect 97960 157564 97966 157576
rect 193214 157564 193220 157576
rect 193272 157564 193278 157616
rect 197354 157564 197360 157616
rect 197412 157604 197418 157616
rect 251450 157604 251456 157616
rect 197412 157576 251456 157604
rect 197412 157564 197418 157576
rect 251450 157564 251456 157576
rect 251508 157564 251514 157616
rect 111334 157496 111340 157548
rect 111392 157536 111398 157548
rect 203426 157536 203432 157548
rect 111392 157508 203432 157536
rect 111392 157496 111398 157508
rect 203426 157496 203432 157508
rect 203484 157496 203490 157548
rect 204898 157496 204904 157548
rect 204956 157536 204962 157548
rect 258074 157536 258080 157548
rect 204956 157508 258080 157536
rect 204956 157496 204962 157508
rect 258074 157496 258080 157508
rect 258132 157496 258138 157548
rect 114738 157428 114744 157480
rect 114796 157468 114802 157480
rect 206554 157468 206560 157480
rect 114796 157440 206560 157468
rect 114796 157428 114802 157440
rect 206554 157428 206560 157440
rect 206612 157428 206618 157480
rect 141694 157360 141700 157412
rect 141752 157400 141758 157412
rect 227070 157400 227076 157412
rect 141752 157372 227076 157400
rect 141752 157360 141758 157372
rect 227070 157360 227076 157372
rect 227128 157360 227134 157412
rect 55858 157292 55864 157344
rect 55916 157332 55922 157344
rect 161566 157332 161572 157344
rect 55916 157304 161572 157332
rect 55916 157292 55922 157304
rect 161566 157292 161572 157304
rect 161624 157292 161630 157344
rect 204898 157332 204904 157344
rect 171106 157304 204904 157332
rect 52454 157224 52460 157276
rect 52512 157264 52518 157276
rect 158990 157264 158996 157276
rect 52512 157236 158996 157264
rect 52512 157224 52518 157236
rect 158990 157224 158996 157236
rect 159048 157224 159054 157276
rect 160094 157224 160100 157276
rect 160152 157264 160158 157276
rect 171106 157264 171134 157304
rect 204898 157292 204904 157304
rect 204956 157292 204962 157344
rect 204990 157292 204996 157344
rect 205048 157332 205054 157344
rect 273254 157332 273260 157344
rect 205048 157304 273260 157332
rect 205048 157292 205054 157304
rect 273254 157292 273260 157304
rect 273312 157292 273318 157344
rect 160152 157236 171134 157264
rect 160152 157224 160158 157236
rect 192110 157224 192116 157276
rect 192168 157264 192174 157276
rect 265158 157264 265164 157276
rect 192168 157236 265164 157264
rect 192168 157224 192174 157236
rect 265158 157224 265164 157236
rect 265216 157224 265222 157276
rect 290550 157224 290556 157276
rect 290608 157264 290614 157276
rect 339954 157264 339960 157276
rect 290608 157236 339960 157264
rect 290608 157224 290614 157236
rect 339954 157224 339960 157236
rect 340012 157224 340018 157276
rect 45738 157156 45744 157208
rect 45796 157196 45802 157208
rect 153746 157196 153752 157208
rect 45796 157168 153752 157196
rect 45796 157156 45802 157168
rect 153746 157156 153752 157168
rect 153804 157156 153810 157208
rect 166902 157156 166908 157208
rect 166960 157196 166966 157208
rect 246298 157196 246304 157208
rect 166960 157168 246304 157196
rect 166960 157156 166966 157168
rect 246298 157156 246304 157168
rect 246356 157156 246362 157208
rect 280430 157156 280436 157208
rect 280488 157196 280494 157208
rect 332686 157196 332692 157208
rect 280488 157168 332692 157196
rect 280488 157156 280494 157168
rect 332686 157156 332692 157168
rect 332744 157156 332750 157208
rect 39022 157088 39028 157140
rect 39080 157128 39086 157140
rect 143718 157128 143724 157140
rect 39080 157100 143724 157128
rect 39080 157088 39086 157100
rect 143718 157088 143724 157100
rect 143776 157088 143782 157140
rect 145466 157128 145472 157140
rect 143828 157100 145472 157128
rect 35710 157020 35716 157072
rect 35768 157060 35774 157072
rect 143828 157060 143856 157100
rect 145466 157088 145472 157100
rect 145524 157088 145530 157140
rect 151722 157088 151728 157140
rect 151780 157128 151786 157140
rect 234798 157128 234804 157140
rect 151780 157100 234804 157128
rect 151780 157088 151786 157100
rect 234798 157088 234804 157100
rect 234856 157088 234862 157140
rect 273714 157088 273720 157140
rect 273772 157128 273778 157140
rect 327902 157128 327908 157140
rect 273772 157100 327908 157128
rect 273772 157088 273778 157100
rect 327902 157088 327908 157100
rect 327960 157088 327966 157140
rect 35768 157032 143856 157060
rect 35768 157020 35774 157032
rect 145282 157020 145288 157072
rect 145340 157060 145346 157072
rect 229646 157060 229652 157072
rect 145340 157032 229652 157060
rect 145340 157020 145346 157032
rect 229646 157020 229652 157032
rect 229704 157020 229710 157072
rect 277118 157020 277124 157072
rect 277176 157060 277182 157072
rect 330478 157060 330484 157072
rect 277176 157032 330484 157060
rect 277176 157020 277182 157032
rect 330478 157020 330484 157032
rect 330536 157020 330542 157072
rect 24762 156952 24768 157004
rect 24820 156992 24826 157004
rect 137186 156992 137192 157004
rect 24820 156964 137192 156992
rect 24820 156952 24826 156964
rect 137186 156952 137192 156964
rect 137244 156952 137250 157004
rect 139118 156952 139124 157004
rect 139176 156992 139182 157004
rect 225138 156992 225144 157004
rect 139176 156964 225144 156992
rect 139176 156952 139182 156964
rect 225138 156952 225144 156964
rect 225196 156952 225202 157004
rect 270310 156952 270316 157004
rect 270368 156992 270374 157004
rect 325326 156992 325332 157004
rect 270368 156964 325332 156992
rect 270368 156952 270374 156964
rect 325326 156952 325332 156964
rect 325384 156952 325390 157004
rect 18046 156884 18052 156936
rect 18104 156924 18110 156936
rect 132494 156924 132500 156936
rect 18104 156896 132500 156924
rect 18104 156884 18110 156896
rect 132494 156884 132500 156896
rect 132552 156884 132558 156936
rect 134886 156884 134892 156936
rect 134944 156924 134950 156936
rect 213822 156924 213828 156936
rect 134944 156896 213828 156924
rect 134944 156884 134950 156896
rect 213822 156884 213828 156896
rect 213880 156884 213886 156936
rect 213914 156884 213920 156936
rect 213972 156924 213978 156936
rect 223114 156924 223120 156936
rect 213972 156896 223120 156924
rect 213972 156884 213978 156896
rect 223114 156884 223120 156896
rect 223172 156884 223178 156936
rect 226610 156884 226616 156936
rect 226668 156924 226674 156936
rect 291930 156924 291936 156936
rect 226668 156896 291936 156924
rect 226668 156884 226674 156896
rect 291930 156884 291936 156896
rect 291988 156884 291994 156936
rect 21358 156816 21364 156868
rect 21416 156856 21422 156868
rect 135254 156856 135260 156868
rect 21416 156828 135260 156856
rect 21416 156816 21422 156828
rect 135254 156816 135260 156828
rect 135312 156816 135318 156868
rect 135806 156816 135812 156868
rect 135864 156856 135870 156868
rect 222562 156856 222568 156868
rect 135864 156828 222568 156856
rect 135864 156816 135870 156828
rect 222562 156816 222568 156828
rect 222620 156816 222626 156868
rect 230014 156816 230020 156868
rect 230072 156856 230078 156868
rect 294046 156856 294052 156868
rect 230072 156828 294052 156856
rect 230072 156816 230078 156828
rect 294046 156816 294052 156828
rect 294104 156816 294110 156868
rect 297266 156816 297272 156868
rect 297324 156856 297330 156868
rect 345842 156856 345848 156868
rect 297324 156828 345848 156856
rect 297324 156816 297330 156828
rect 345842 156816 345848 156828
rect 345900 156816 345906 156868
rect 11238 156748 11244 156800
rect 11296 156788 11302 156800
rect 127526 156788 127532 156800
rect 11296 156760 127532 156788
rect 11296 156748 11302 156760
rect 127526 156748 127532 156760
rect 127584 156748 127590 156800
rect 128170 156748 128176 156800
rect 128228 156788 128234 156800
rect 216766 156788 216772 156800
rect 128228 156760 216772 156788
rect 128228 156748 128234 156760
rect 216766 156748 216772 156760
rect 216824 156748 216830 156800
rect 219894 156748 219900 156800
rect 219952 156788 219958 156800
rect 285674 156788 285680 156800
rect 219952 156760 285680 156788
rect 219952 156748 219958 156760
rect 285674 156748 285680 156760
rect 285732 156748 285738 156800
rect 287146 156748 287152 156800
rect 287204 156788 287210 156800
rect 338114 156788 338120 156800
rect 287204 156760 338120 156788
rect 287204 156748 287210 156760
rect 338114 156748 338120 156760
rect 338172 156748 338178 156800
rect 14642 156680 14648 156732
rect 14700 156720 14706 156732
rect 130102 156720 130108 156732
rect 14700 156692 130108 156720
rect 14700 156680 14706 156692
rect 130102 156680 130108 156692
rect 130160 156680 130166 156732
rect 132402 156680 132408 156732
rect 132460 156720 132466 156732
rect 219986 156720 219992 156732
rect 132460 156692 219992 156720
rect 132460 156680 132466 156692
rect 219986 156680 219992 156692
rect 220044 156680 220050 156732
rect 223206 156680 223212 156732
rect 223264 156720 223270 156732
rect 289354 156720 289360 156732
rect 223264 156692 289360 156720
rect 223264 156680 223270 156692
rect 289354 156680 289360 156692
rect 289412 156680 289418 156732
rect 293862 156680 293868 156732
rect 293920 156720 293926 156732
rect 343266 156720 343272 156732
rect 293920 156692 343272 156720
rect 293920 156680 293926 156692
rect 343266 156680 343272 156692
rect 343324 156680 343330 156732
rect 344370 156680 344376 156732
rect 344428 156720 344434 156732
rect 381814 156720 381820 156732
rect 344428 156692 381820 156720
rect 344428 156680 344434 156692
rect 381814 156680 381820 156692
rect 381872 156680 381878 156732
rect 2038 156612 2044 156664
rect 2096 156652 2102 156664
rect 120442 156652 120448 156664
rect 2096 156624 120448 156652
rect 2096 156612 2102 156624
rect 120442 156612 120448 156624
rect 120500 156612 120506 156664
rect 121454 156612 121460 156664
rect 121512 156652 121518 156664
rect 201310 156652 201316 156664
rect 121512 156624 201316 156652
rect 121512 156612 121518 156624
rect 201310 156612 201316 156624
rect 201368 156612 201374 156664
rect 219894 156652 219900 156664
rect 201420 156624 219900 156652
rect 143718 156544 143724 156596
rect 143776 156584 143782 156596
rect 147674 156584 147680 156596
rect 143776 156556 147680 156584
rect 143776 156544 143782 156556
rect 147674 156544 147680 156556
rect 147732 156544 147738 156596
rect 158714 156544 158720 156596
rect 158772 156584 158778 156596
rect 201420 156584 201448 156624
rect 219894 156612 219900 156624
rect 219952 156612 219958 156664
rect 220078 156612 220084 156664
rect 220136 156652 220142 156664
rect 281626 156652 281632 156664
rect 220136 156624 281632 156652
rect 220136 156612 220142 156624
rect 281626 156612 281632 156624
rect 281684 156612 281690 156664
rect 283834 156612 283840 156664
rect 283892 156652 283898 156664
rect 335538 156652 335544 156664
rect 283892 156624 335544 156652
rect 283892 156612 283898 156624
rect 335538 156612 335544 156624
rect 335596 156612 335602 156664
rect 337654 156612 337660 156664
rect 337712 156652 337718 156664
rect 375558 156652 375564 156664
rect 337712 156624 375564 156652
rect 337712 156612 337718 156624
rect 375558 156612 375564 156624
rect 375616 156612 375622 156664
rect 270494 156584 270500 156596
rect 158772 156556 201448 156584
rect 201512 156556 270500 156584
rect 158772 156544 158778 156556
rect 72694 156476 72700 156528
rect 72752 156516 72758 156528
rect 174446 156516 174452 156528
rect 72752 156488 174452 156516
rect 72752 156476 72758 156488
rect 174446 156476 174452 156488
rect 174504 156476 174510 156528
rect 174630 156476 174636 156528
rect 174688 156516 174694 156528
rect 174688 156488 180794 156516
rect 174688 156476 174694 156488
rect 79410 156408 79416 156460
rect 79468 156448 79474 156460
rect 179598 156448 179604 156460
rect 79468 156420 179604 156448
rect 79468 156408 79474 156420
rect 179598 156408 179604 156420
rect 179656 156408 179662 156460
rect 180766 156448 180794 156488
rect 198826 156476 198832 156528
rect 198884 156516 198890 156528
rect 201512 156516 201540 156556
rect 270494 156544 270500 156556
rect 270552 156544 270558 156596
rect 198884 156488 201540 156516
rect 198884 156476 198890 156488
rect 204898 156476 204904 156528
rect 204956 156516 204962 156528
rect 213914 156516 213920 156528
rect 204956 156488 213920 156516
rect 204956 156476 204962 156488
rect 213914 156476 213920 156488
rect 213972 156476 213978 156528
rect 214558 156476 214564 156528
rect 214616 156516 214622 156528
rect 273898 156516 273904 156528
rect 214616 156488 273904 156516
rect 214616 156476 214622 156488
rect 273898 156476 273904 156488
rect 273956 156476 273962 156528
rect 180766 156420 196388 156448
rect 92842 156340 92848 156392
rect 92900 156380 92906 156392
rect 189810 156380 189816 156392
rect 92900 156352 189816 156380
rect 92900 156340 92906 156352
rect 189810 156340 189816 156352
rect 189868 156340 189874 156392
rect 101306 156272 101312 156324
rect 101364 156312 101370 156324
rect 196250 156312 196256 156324
rect 101364 156284 196256 156312
rect 101364 156272 101370 156284
rect 196250 156272 196256 156284
rect 196308 156272 196314 156324
rect 196360 156312 196388 156420
rect 201310 156408 201316 156460
rect 201368 156448 201374 156460
rect 211614 156448 211620 156460
rect 201368 156420 211620 156448
rect 201368 156408 201374 156420
rect 211614 156408 211620 156420
rect 211672 156408 211678 156460
rect 279050 156448 279056 156460
rect 211724 156420 279056 156448
rect 202230 156340 202236 156392
rect 202288 156380 202294 156392
rect 204990 156380 204996 156392
rect 202288 156352 204996 156380
rect 202288 156340 202294 156352
rect 204990 156340 204996 156352
rect 205048 156340 205054 156392
rect 209774 156340 209780 156392
rect 209832 156380 209838 156392
rect 211724 156380 211752 156420
rect 279050 156408 279056 156420
rect 279108 156408 279114 156460
rect 209832 156352 211752 156380
rect 212506 156352 216444 156380
rect 209832 156340 209838 156352
rect 212506 156312 212534 156352
rect 196360 156284 212534 156312
rect 216416 156312 216444 156352
rect 216490 156340 216496 156392
rect 216548 156380 216554 156392
rect 283098 156380 283104 156392
rect 216548 156352 283104 156380
rect 216548 156340 216554 156352
rect 283098 156340 283104 156352
rect 283156 156340 283162 156392
rect 230934 156312 230940 156324
rect 216416 156284 230940 156312
rect 230934 156272 230940 156284
rect 230992 156272 230998 156324
rect 108022 156204 108028 156256
rect 108080 156244 108086 156256
rect 200298 156244 200304 156256
rect 108080 156216 200304 156244
rect 108080 156204 108086 156216
rect 200298 156204 200304 156216
rect 200356 156204 200362 156256
rect 203058 156204 203064 156256
rect 203116 156244 203122 156256
rect 214558 156244 214564 156256
rect 203116 156216 214564 156244
rect 203116 156204 203122 156216
rect 214558 156204 214564 156216
rect 214616 156204 214622 156256
rect 222102 156204 222108 156256
rect 222160 156244 222166 156256
rect 269206 156244 269212 156256
rect 222160 156216 269212 156244
rect 222160 156204 222166 156216
rect 269206 156204 269212 156216
rect 269264 156204 269270 156256
rect 118142 156136 118148 156188
rect 118200 156176 118206 156188
rect 209130 156176 209136 156188
rect 118200 156148 209136 156176
rect 118200 156136 118206 156148
rect 209130 156136 209136 156148
rect 209188 156136 209194 156188
rect 213178 156136 213184 156188
rect 213236 156176 213242 156188
rect 220078 156176 220084 156188
rect 213236 156148 220084 156176
rect 213236 156136 213242 156148
rect 220078 156136 220084 156148
rect 220136 156136 220142 156188
rect 220630 156136 220636 156188
rect 220688 156176 220694 156188
rect 266906 156176 266912 156188
rect 220688 156148 266912 156176
rect 220688 156136 220694 156148
rect 266906 156136 266912 156148
rect 266964 156136 266970 156188
rect 124858 156068 124864 156120
rect 124916 156108 124922 156120
rect 213914 156108 213920 156120
rect 124916 156080 213920 156108
rect 124916 156068 124922 156080
rect 213914 156068 213920 156080
rect 213972 156068 213978 156120
rect 219894 156068 219900 156120
rect 219952 156108 219958 156120
rect 220538 156108 220544 156120
rect 219952 156080 220544 156108
rect 219952 156068 219958 156080
rect 220538 156068 220544 156080
rect 220596 156068 220602 156120
rect 227714 156068 227720 156120
rect 227772 156108 227778 156120
rect 272058 156108 272064 156120
rect 227772 156080 272064 156108
rect 227772 156068 227778 156080
rect 272058 156068 272064 156080
rect 272116 156068 272122 156120
rect 138290 156000 138296 156052
rect 138348 156040 138354 156052
rect 224494 156040 224500 156052
rect 138348 156012 224500 156040
rect 138348 156000 138354 156012
rect 224494 156000 224500 156012
rect 224552 156000 224558 156052
rect 59262 155932 59268 155984
rect 59320 155972 59326 155984
rect 164142 155972 164148 155984
rect 59320 155944 164148 155972
rect 59320 155932 59326 155944
rect 164142 155932 164148 155944
rect 164200 155932 164206 155984
rect 164234 155932 164240 155984
rect 164292 155972 164298 155984
rect 228358 155972 228364 155984
rect 164292 155944 228364 155972
rect 164292 155932 164298 155944
rect 228358 155932 228364 155944
rect 228416 155932 228422 155984
rect 60090 155864 60096 155916
rect 60148 155904 60154 155916
rect 85482 155904 85488 155916
rect 60148 155876 85488 155904
rect 60148 155864 60154 155876
rect 85482 155864 85488 155876
rect 85540 155864 85546 155916
rect 88702 155864 88708 155916
rect 88760 155904 88766 155916
rect 186774 155904 186780 155916
rect 88760 155876 186780 155904
rect 88760 155864 88766 155876
rect 186774 155864 186780 155876
rect 186832 155864 186838 155916
rect 189626 155864 189632 155916
rect 189684 155904 189690 155916
rect 263686 155904 263692 155916
rect 189684 155876 263692 155904
rect 189684 155864 189690 155876
rect 263686 155864 263692 155876
rect 263744 155864 263750 155916
rect 303154 155864 303160 155916
rect 303212 155904 303218 155916
rect 350350 155904 350356 155916
rect 303212 155876 350356 155904
rect 303212 155864 303218 155876
rect 350350 155864 350356 155876
rect 350408 155864 350414 155916
rect 12158 155796 12164 155848
rect 12216 155836 12222 155848
rect 109678 155836 109684 155848
rect 12216 155808 109684 155836
rect 12216 155796 12222 155808
rect 109678 155796 109684 155808
rect 109736 155796 109742 155848
rect 112254 155796 112260 155848
rect 112312 155836 112318 155848
rect 204622 155836 204628 155848
rect 112312 155808 204628 155836
rect 112312 155796 112318 155808
rect 204622 155796 204628 155808
rect 204680 155796 204686 155848
rect 206462 155796 206468 155848
rect 206520 155836 206526 155848
rect 276014 155836 276020 155848
rect 206520 155808 276020 155836
rect 206520 155796 206526 155808
rect 276014 155796 276020 155808
rect 276072 155796 276078 155848
rect 293034 155796 293040 155848
rect 293092 155836 293098 155848
rect 342622 155836 342628 155848
rect 293092 155808 342628 155836
rect 293092 155796 293098 155808
rect 342622 155796 342628 155808
rect 342680 155796 342686 155848
rect 53374 155728 53380 155780
rect 53432 155768 53438 155780
rect 76742 155768 76748 155780
rect 53432 155740 76748 155768
rect 53432 155728 53438 155740
rect 76742 155728 76748 155740
rect 76800 155728 76806 155780
rect 81894 155728 81900 155780
rect 81952 155768 81958 155780
rect 181438 155768 181444 155780
rect 81952 155740 181444 155768
rect 81952 155728 81958 155740
rect 181438 155728 181444 155740
rect 181496 155728 181502 155780
rect 186222 155728 186228 155780
rect 186280 155768 186286 155780
rect 260834 155768 260840 155780
rect 186280 155740 260840 155768
rect 186280 155728 186286 155740
rect 260834 155728 260840 155740
rect 260892 155728 260898 155780
rect 296438 155728 296444 155780
rect 296496 155768 296502 155780
rect 345198 155768 345204 155780
rect 296496 155740 345204 155768
rect 296496 155728 296502 155740
rect 345198 155728 345204 155740
rect 345256 155728 345262 155780
rect 33134 155660 33140 155712
rect 33192 155700 33198 155712
rect 59998 155700 60004 155712
rect 33192 155672 60004 155700
rect 33192 155660 33198 155672
rect 59998 155660 60004 155672
rect 60056 155660 60062 155712
rect 71866 155660 71872 155712
rect 71924 155700 71930 155712
rect 173066 155700 173072 155712
rect 71924 155672 173072 155700
rect 71924 155660 71930 155672
rect 173066 155660 173072 155672
rect 173124 155660 173130 155712
rect 176286 155660 176292 155712
rect 176344 155700 176350 155712
rect 176344 155672 176516 155700
rect 176344 155660 176350 155672
rect 46566 155592 46572 155644
rect 46624 155632 46630 155644
rect 75086 155632 75092 155644
rect 46624 155604 75092 155632
rect 46624 155592 46630 155604
rect 75086 155592 75092 155604
rect 75144 155592 75150 155644
rect 75178 155592 75184 155644
rect 75236 155632 75242 155644
rect 176378 155632 176384 155644
rect 75236 155604 176384 155632
rect 75236 155592 75242 155604
rect 176378 155592 176384 155604
rect 176436 155592 176442 155644
rect 176488 155632 176516 155672
rect 177114 155660 177120 155712
rect 177172 155700 177178 155712
rect 254026 155700 254032 155712
rect 177172 155672 254032 155700
rect 177172 155660 177178 155672
rect 254026 155660 254032 155672
rect 254084 155660 254090 155712
rect 289722 155660 289728 155712
rect 289780 155700 289786 155712
rect 339586 155700 339592 155712
rect 289780 155672 339592 155700
rect 289780 155660 289786 155672
rect 339586 155660 339592 155672
rect 339644 155660 339650 155712
rect 253382 155632 253388 155644
rect 176488 155604 253388 155632
rect 253382 155592 253388 155604
rect 253440 155592 253446 155644
rect 266998 155592 267004 155644
rect 267056 155632 267062 155644
rect 322106 155632 322112 155644
rect 267056 155604 322112 155632
rect 267056 155592 267062 155604
rect 322106 155592 322112 155604
rect 322164 155592 322170 155644
rect 39850 155524 39856 155576
rect 39908 155564 39914 155576
rect 71774 155564 71780 155576
rect 39908 155536 71780 155564
rect 39908 155524 39914 155536
rect 71774 155524 71780 155536
rect 71832 155524 71838 155576
rect 78582 155524 78588 155576
rect 78640 155564 78646 155576
rect 178954 155564 178960 155576
rect 78640 155536 178960 155564
rect 78640 155524 78646 155536
rect 178954 155524 178960 155536
rect 179012 155524 179018 155576
rect 179506 155524 179512 155576
rect 179564 155564 179570 155576
rect 255866 155564 255872 155576
rect 179564 155536 255872 155564
rect 179564 155524 179570 155536
rect 255866 155524 255872 155536
rect 255924 155524 255930 155576
rect 263594 155524 263600 155576
rect 263652 155564 263658 155576
rect 320174 155564 320180 155576
rect 263652 155536 320180 155564
rect 263652 155524 263658 155536
rect 320174 155524 320180 155536
rect 320232 155524 320238 155576
rect 340966 155524 340972 155576
rect 341024 155564 341030 155576
rect 378134 155564 378140 155576
rect 341024 155536 378140 155564
rect 341024 155524 341030 155536
rect 378134 155524 378140 155536
rect 378192 155524 378198 155576
rect 28902 155456 28908 155508
rect 28960 155496 28966 155508
rect 56226 155496 56232 155508
rect 28960 155468 56232 155496
rect 28960 155456 28966 155468
rect 56226 155456 56232 155468
rect 56284 155456 56290 155508
rect 62574 155456 62580 155508
rect 62632 155496 62638 155508
rect 165614 155496 165620 155508
rect 62632 155468 165620 155496
rect 62632 155456 62638 155468
rect 165614 155456 165620 155468
rect 165672 155456 165678 155508
rect 169386 155456 169392 155508
rect 169444 155496 169450 155508
rect 247126 155496 247132 155508
rect 169444 155468 247132 155496
rect 169444 155456 169450 155468
rect 247126 155456 247132 155468
rect 247184 155456 247190 155508
rect 260282 155456 260288 155508
rect 260340 155496 260346 155508
rect 317598 155496 317604 155508
rect 260340 155468 317604 155496
rect 260340 155456 260346 155468
rect 317598 155456 317604 155468
rect 317656 155456 317662 155508
rect 333422 155456 333428 155508
rect 333480 155496 333486 155508
rect 373442 155496 373448 155508
rect 333480 155468 373448 155496
rect 333480 155456 333486 155468
rect 373442 155456 373448 155468
rect 373500 155456 373506 155508
rect 7926 155388 7932 155440
rect 7984 155428 7990 155440
rect 122006 155428 122012 155440
rect 7984 155400 122012 155428
rect 7984 155388 7990 155400
rect 122006 155388 122012 155400
rect 122064 155388 122070 155440
rect 125594 155428 125600 155440
rect 122116 155400 125600 155428
rect 4522 155320 4528 155372
rect 4580 155360 4586 155372
rect 121914 155360 121920 155372
rect 4580 155332 121920 155360
rect 4580 155320 4586 155332
rect 121914 155320 121920 155332
rect 121972 155320 121978 155372
rect 8754 155252 8760 155304
rect 8812 155292 8818 155304
rect 122116 155292 122144 155400
rect 125594 155388 125600 155400
rect 125652 155388 125658 155440
rect 134058 155388 134064 155440
rect 134116 155428 134122 155440
rect 137462 155428 137468 155440
rect 134116 155400 137468 155428
rect 134116 155388 134122 155400
rect 137462 155388 137468 155400
rect 137520 155388 137526 155440
rect 142522 155388 142528 155440
rect 142580 155428 142586 155440
rect 227714 155428 227720 155440
rect 142580 155400 227720 155428
rect 142580 155388 142586 155400
rect 227714 155388 227720 155400
rect 227772 155388 227778 155440
rect 250162 155388 250168 155440
rect 250220 155428 250226 155440
rect 309870 155428 309876 155440
rect 250220 155400 309876 155428
rect 250220 155388 250226 155400
rect 309870 155388 309876 155400
rect 309928 155388 309934 155440
rect 330110 155388 330116 155440
rect 330168 155428 330174 155440
rect 369854 155428 369860 155440
rect 330168 155400 369860 155428
rect 330168 155388 330174 155400
rect 369854 155388 369860 155400
rect 369912 155388 369918 155440
rect 122282 155320 122288 155372
rect 122340 155360 122346 155372
rect 211246 155360 211252 155372
rect 122340 155332 211252 155360
rect 122340 155320 122346 155332
rect 211246 155320 211252 155332
rect 211304 155320 211310 155372
rect 213822 155320 213828 155372
rect 213880 155360 213886 155372
rect 213880 155332 214972 155360
rect 213880 155320 213886 155332
rect 8812 155264 122144 155292
rect 8812 155252 8818 155264
rect 125686 155252 125692 155304
rect 125744 155292 125750 155304
rect 214834 155292 214840 155304
rect 125744 155264 214840 155292
rect 125744 155252 125750 155264
rect 214834 155252 214840 155264
rect 214892 155252 214898 155304
rect 214944 155292 214972 155332
rect 216674 155320 216680 155372
rect 216732 155360 216738 155372
rect 261386 155360 261392 155372
rect 216732 155332 261392 155360
rect 216732 155320 216738 155332
rect 261386 155320 261392 155332
rect 261444 155320 261450 155372
rect 263594 155320 263600 155372
rect 263652 155360 263658 155372
rect 263778 155360 263784 155372
rect 263652 155332 263784 155360
rect 263652 155320 263658 155332
rect 263778 155320 263784 155332
rect 263836 155320 263842 155372
rect 316586 155320 316592 155372
rect 316644 155360 316650 155372
rect 360654 155360 360660 155372
rect 316644 155332 360660 155360
rect 316644 155320 316650 155332
rect 360654 155320 360660 155332
rect 360712 155320 360718 155372
rect 221918 155292 221924 155304
rect 214944 155264 221924 155292
rect 221918 155252 221924 155264
rect 221976 155252 221982 155304
rect 243446 155252 243452 155304
rect 243504 155292 243510 155304
rect 304718 155292 304724 155304
rect 243504 155264 304724 155292
rect 243504 155252 243510 155264
rect 304718 155252 304724 155264
rect 304776 155252 304782 155304
rect 309962 155252 309968 155304
rect 310020 155292 310026 155304
rect 354674 155292 354680 155304
rect 310020 155264 354680 155292
rect 310020 155252 310026 155264
rect 354674 155252 354680 155264
rect 354732 155252 354738 155304
rect 373810 155252 373816 155304
rect 373868 155292 373874 155304
rect 403158 155292 403164 155304
rect 373868 155264 403164 155292
rect 373868 155252 373874 155264
rect 403158 155252 403164 155264
rect 403216 155252 403222 155304
rect 5350 155184 5356 155236
rect 5408 155224 5414 155236
rect 123018 155224 123024 155236
rect 5408 155196 123024 155224
rect 5408 155184 5414 155196
rect 123018 155184 123024 155196
rect 123076 155184 123082 155236
rect 128998 155184 129004 155236
rect 129056 155224 129062 155236
rect 217410 155224 217416 155236
rect 129056 155196 217416 155224
rect 129056 155184 129062 155196
rect 217410 155184 217416 155196
rect 217468 155184 217474 155236
rect 236730 155184 236736 155236
rect 236788 155224 236794 155236
rect 299658 155224 299664 155236
rect 236788 155196 299664 155224
rect 236788 155184 236794 155196
rect 299658 155184 299664 155196
rect 299716 155184 299722 155236
rect 299750 155184 299756 155236
rect 299808 155224 299814 155236
rect 347774 155224 347780 155236
rect 299808 155196 347780 155224
rect 299808 155184 299814 155196
rect 347774 155184 347780 155196
rect 347832 155184 347838 155236
rect 367094 155184 367100 155236
rect 367152 155224 367158 155236
rect 399110 155224 399116 155236
rect 367152 155196 399116 155224
rect 367152 155184 367158 155196
rect 399110 155184 399116 155196
rect 399168 155184 399174 155236
rect 401594 155184 401600 155236
rect 401652 155224 401658 155236
rect 425514 155224 425520 155236
rect 401652 155196 425520 155224
rect 401652 155184 401658 155196
rect 425514 155184 425520 155196
rect 425572 155184 425578 155236
rect 86126 155116 86132 155168
rect 86184 155156 86190 155168
rect 183554 155156 183560 155168
rect 86184 155128 183560 155156
rect 86184 155116 86190 155128
rect 183554 155116 183560 155128
rect 183612 155116 183618 155168
rect 186682 155116 186688 155168
rect 186740 155156 186746 155168
rect 186740 155128 192892 155156
rect 186740 155116 186746 155128
rect 95418 155048 95424 155100
rect 95476 155088 95482 155100
rect 186314 155088 186320 155100
rect 95476 155060 186320 155088
rect 95476 155048 95482 155060
rect 186314 155048 186320 155060
rect 186372 155048 186378 155100
rect 186498 155048 186504 155100
rect 186556 155088 186562 155100
rect 191742 155088 191748 155100
rect 186556 155060 191748 155088
rect 186556 155048 186562 155060
rect 191742 155048 191748 155060
rect 191800 155048 191806 155100
rect 192864 155088 192892 155128
rect 192938 155116 192944 155168
rect 192996 155156 193002 155168
rect 266078 155156 266084 155168
rect 192996 155128 266084 155156
rect 192996 155116 193002 155128
rect 266078 155116 266084 155128
rect 266136 155116 266142 155168
rect 306558 155116 306564 155168
rect 306616 155156 306622 155168
rect 352926 155156 352932 155168
rect 306616 155128 352932 155156
rect 306616 155116 306622 155128
rect 352926 155116 352932 155128
rect 352984 155116 352990 155168
rect 194962 155088 194968 155100
rect 192864 155060 194968 155088
rect 194962 155048 194968 155060
rect 195020 155048 195026 155100
rect 196342 155048 196348 155100
rect 196400 155088 196406 155100
rect 268838 155088 268844 155100
rect 196400 155060 268844 155088
rect 196400 155048 196406 155060
rect 268838 155048 268844 155060
rect 268896 155048 268902 155100
rect 98730 154980 98736 155032
rect 98788 155020 98794 155032
rect 186222 155020 186228 155032
rect 98788 154992 186228 155020
rect 98788 154980 98794 154992
rect 186222 154980 186228 154992
rect 186280 154980 186286 155032
rect 186590 154980 186596 155032
rect 186648 155020 186654 155032
rect 194318 155020 194324 155032
rect 186648 154992 194324 155020
rect 186648 154980 186654 154992
rect 194318 154980 194324 154992
rect 194376 154980 194382 155032
rect 199654 154980 199660 155032
rect 199712 155020 199718 155032
rect 271414 155020 271420 155032
rect 199712 154992 271420 155020
rect 199712 154980 199718 154992
rect 271414 154980 271420 154992
rect 271472 154980 271478 155032
rect 80238 154912 80244 154964
rect 80296 154952 80302 154964
rect 86862 154952 86868 154964
rect 80296 154924 86868 154952
rect 80296 154912 80302 154924
rect 86862 154912 86868 154924
rect 86920 154912 86926 154964
rect 99558 154912 99564 154964
rect 99616 154952 99622 154964
rect 186314 154952 186320 154964
rect 99616 154924 186320 154952
rect 99616 154912 99622 154924
rect 186314 154912 186320 154924
rect 186372 154912 186378 154964
rect 188338 154912 188344 154964
rect 188396 154952 188402 154964
rect 240686 154952 240692 154964
rect 188396 154924 240692 154952
rect 188396 154912 188402 154924
rect 240686 154912 240692 154924
rect 240744 154912 240750 154964
rect 253566 154912 253572 154964
rect 253624 154952 253630 154964
rect 312446 154952 312452 154964
rect 253624 154924 312452 154952
rect 253624 154912 253630 154924
rect 312446 154912 312452 154924
rect 312504 154912 312510 154964
rect 107102 154844 107108 154896
rect 107160 154884 107166 154896
rect 133322 154884 133328 154896
rect 107160 154856 133328 154884
rect 107160 154844 107166 154856
rect 133322 154844 133328 154856
rect 133380 154844 133386 154896
rect 145834 154844 145840 154896
rect 145892 154884 145898 154896
rect 229186 154884 229192 154896
rect 145892 154856 229192 154884
rect 145892 154844 145898 154856
rect 229186 154844 229192 154856
rect 229244 154844 229250 154896
rect 231302 154844 231308 154896
rect 231360 154884 231366 154896
rect 277118 154884 277124 154896
rect 231360 154856 277124 154884
rect 231360 154844 231366 154856
rect 277118 154844 277124 154856
rect 277176 154844 277182 154896
rect 110506 154776 110512 154828
rect 110564 154816 110570 154828
rect 128354 154816 128360 154828
rect 110564 154788 128360 154816
rect 110564 154776 110570 154788
rect 128354 154776 128360 154788
rect 128412 154776 128418 154828
rect 149238 154776 149244 154828
rect 149296 154816 149302 154828
rect 232866 154816 232872 154828
rect 149296 154788 232872 154816
rect 149296 154776 149302 154788
rect 232866 154776 232872 154788
rect 232924 154776 232930 154828
rect 122006 154708 122012 154760
rect 122064 154748 122070 154760
rect 124950 154748 124956 154760
rect 122064 154720 124956 154748
rect 122064 154708 122070 154720
rect 124950 154708 124956 154720
rect 125008 154708 125014 154760
rect 155954 154708 155960 154760
rect 156012 154748 156018 154760
rect 238018 154748 238024 154760
rect 156012 154720 238024 154748
rect 156012 154708 156018 154720
rect 238018 154708 238024 154720
rect 238076 154708 238082 154760
rect 118970 154640 118976 154692
rect 119028 154680 119034 154692
rect 124398 154680 124404 154692
rect 119028 154652 124404 154680
rect 119028 154640 119034 154652
rect 124398 154640 124404 154652
rect 124456 154640 124462 154692
rect 146202 154640 146208 154692
rect 146260 154680 146266 154692
rect 146260 154652 150756 154680
rect 146260 154640 146266 154652
rect 121914 154572 121920 154624
rect 121972 154612 121978 154624
rect 122374 154612 122380 154624
rect 121972 154584 122380 154612
rect 121972 154572 121978 154584
rect 122374 154572 122380 154584
rect 122432 154572 122438 154624
rect 44910 154504 44916 154556
rect 44968 154544 44974 154556
rect 146478 154544 146484 154556
rect 44968 154516 146484 154544
rect 44968 154504 44974 154516
rect 146478 154504 146484 154516
rect 146536 154504 146542 154556
rect 150618 154544 150624 154556
rect 146680 154516 150624 154544
rect 41598 154436 41604 154488
rect 41656 154476 41662 154488
rect 146680 154476 146708 154516
rect 150618 154504 150624 154516
rect 150676 154504 150682 154556
rect 150728 154544 150756 154652
rect 162670 154640 162676 154692
rect 162728 154680 162734 154692
rect 243078 154680 243084 154692
rect 162728 154652 243084 154680
rect 162728 154640 162734 154652
rect 243078 154640 243084 154652
rect 243136 154640 243142 154692
rect 159358 154572 159364 154624
rect 159416 154612 159422 154624
rect 240134 154612 240140 154624
rect 159416 154584 240140 154612
rect 159416 154572 159422 154584
rect 240134 154572 240140 154584
rect 240192 154572 240198 154624
rect 156782 154544 156788 154556
rect 150728 154516 156788 154544
rect 156782 154504 156788 154516
rect 156840 154504 156846 154556
rect 157334 154504 157340 154556
rect 157392 154544 157398 154556
rect 225782 154544 225788 154556
rect 157392 154516 225788 154544
rect 157392 154504 157398 154516
rect 225782 154504 225788 154516
rect 225840 154504 225846 154556
rect 232498 154504 232504 154556
rect 232556 154544 232562 154556
rect 296438 154544 296444 154556
rect 232556 154516 296444 154544
rect 232556 154504 232562 154516
rect 296438 154504 296444 154516
rect 296496 154504 296502 154556
rect 357342 154504 357348 154556
rect 357400 154544 357406 154556
rect 391474 154544 391480 154556
rect 357400 154516 391480 154544
rect 357400 154504 357406 154516
rect 391474 154504 391480 154516
rect 391532 154504 391538 154556
rect 185118 154476 185124 154488
rect 41656 154448 146708 154476
rect 146772 154448 185124 154476
rect 41656 154436 41662 154448
rect 34790 154368 34796 154420
rect 34848 154408 34854 154420
rect 145374 154408 145380 154420
rect 34848 154380 145380 154408
rect 34848 154368 34854 154380
rect 145374 154368 145380 154380
rect 145432 154368 145438 154420
rect 38470 154300 38476 154352
rect 38528 154340 38534 154352
rect 145098 154340 145104 154352
rect 38528 154312 145104 154340
rect 38528 154300 38534 154312
rect 145098 154300 145104 154312
rect 145156 154300 145162 154352
rect 30650 154232 30656 154284
rect 30708 154272 30714 154284
rect 137094 154272 137100 154284
rect 30708 154244 137100 154272
rect 30708 154232 30714 154244
rect 137094 154232 137100 154244
rect 137152 154232 137158 154284
rect 146772 154272 146800 154448
rect 185118 154436 185124 154448
rect 185176 154436 185182 154488
rect 191282 154436 191288 154488
rect 191340 154476 191346 154488
rect 200114 154476 200120 154488
rect 191340 154448 200120 154476
rect 191340 154436 191346 154448
rect 200114 154436 200120 154448
rect 200172 154436 200178 154488
rect 225874 154436 225880 154488
rect 225932 154476 225938 154488
rect 291286 154476 291292 154488
rect 225932 154448 291292 154476
rect 225932 154436 225938 154448
rect 291286 154436 291292 154448
rect 291344 154436 291350 154488
rect 353662 154436 353668 154488
rect 353720 154476 353726 154488
rect 388898 154476 388904 154488
rect 353720 154448 388904 154476
rect 353720 154436 353726 154448
rect 388898 154436 388904 154448
rect 388956 154436 388962 154488
rect 400766 154436 400772 154488
rect 400824 154476 400830 154488
rect 424870 154476 424876 154488
rect 400824 154448 424876 154476
rect 400824 154436 400830 154448
rect 424870 154436 424876 154448
rect 424928 154436 424934 154488
rect 188430 154408 188436 154420
rect 137204 154244 146800 154272
rect 146864 154380 188436 154408
rect 23934 154164 23940 154216
rect 23992 154204 23998 154216
rect 137002 154204 137008 154216
rect 23992 154176 137008 154204
rect 23992 154164 23998 154176
rect 137002 154164 137008 154176
rect 137060 154164 137066 154216
rect 13814 154096 13820 154148
rect 13872 154136 13878 154148
rect 13872 154108 120764 154136
rect 13872 154096 13878 154108
rect 10410 154028 10416 154080
rect 10468 154068 10474 154080
rect 120626 154068 120632 154080
rect 10468 154040 120632 154068
rect 10468 154028 10474 154040
rect 120626 154028 120632 154040
rect 120684 154028 120690 154080
rect 120736 154068 120764 154108
rect 121546 154096 121552 154148
rect 121604 154136 121610 154148
rect 137204 154136 137232 154244
rect 146864 154204 146892 154380
rect 188430 154368 188436 154380
rect 188488 154368 188494 154420
rect 191466 154368 191472 154420
rect 191524 154408 191530 154420
rect 202690 154408 202696 154420
rect 191524 154380 202696 154408
rect 191524 154368 191530 154380
rect 202690 154368 202696 154380
rect 202748 154368 202754 154420
rect 208946 154368 208952 154420
rect 209004 154408 209010 154420
rect 278406 154408 278412 154420
rect 209004 154380 278412 154408
rect 209004 154368 209010 154380
rect 278406 154368 278412 154380
rect 278464 154368 278470 154420
rect 279970 154368 279976 154420
rect 280028 154408 280034 154420
rect 332410 154408 332416 154420
rect 280028 154380 332416 154408
rect 280028 154368 280034 154380
rect 332410 154368 332416 154380
rect 332468 154368 332474 154420
rect 350258 154368 350264 154420
rect 350316 154408 350322 154420
rect 386322 154408 386328 154420
rect 350316 154380 386328 154408
rect 350316 154368 350322 154380
rect 386322 154368 386328 154380
rect 386380 154368 386386 154420
rect 398190 154368 398196 154420
rect 398248 154408 398254 154420
rect 423030 154408 423036 154420
rect 398248 154380 423036 154408
rect 398248 154368 398254 154380
rect 423030 154368 423036 154380
rect 423088 154368 423094 154420
rect 146938 154300 146944 154352
rect 146996 154340 147002 154352
rect 191282 154340 191288 154352
rect 146996 154312 191288 154340
rect 146996 154300 147002 154312
rect 191282 154300 191288 154312
rect 191340 154300 191346 154352
rect 191374 154300 191380 154352
rect 191432 154340 191438 154352
rect 202046 154340 202052 154352
rect 191432 154312 202052 154340
rect 191432 154300 191438 154312
rect 202046 154300 202052 154312
rect 202104 154300 202110 154352
rect 205542 154300 205548 154352
rect 205600 154340 205606 154352
rect 275830 154340 275836 154352
rect 205600 154312 275836 154340
rect 205600 154300 205606 154312
rect 275830 154300 275836 154312
rect 275888 154300 275894 154352
rect 276198 154300 276204 154352
rect 276256 154340 276262 154352
rect 329834 154340 329840 154352
rect 276256 154312 329840 154340
rect 276256 154300 276262 154312
rect 329834 154300 329840 154312
rect 329892 154300 329898 154352
rect 346854 154300 346860 154352
rect 346912 154340 346918 154352
rect 383746 154340 383752 154352
rect 346912 154312 383752 154340
rect 346912 154300 346918 154312
rect 383746 154300 383752 154312
rect 383804 154300 383810 154352
rect 390646 154300 390652 154352
rect 390704 154340 390710 154352
rect 417142 154340 417148 154352
rect 390704 154312 417148 154340
rect 390704 154300 390710 154312
rect 417142 154300 417148 154312
rect 417200 154300 417206 154352
rect 185210 154272 185216 154284
rect 121604 154108 137232 154136
rect 137296 154176 146892 154204
rect 146956 154244 185216 154272
rect 121604 154096 121610 154108
rect 129458 154068 129464 154080
rect 120736 154040 129464 154068
rect 129458 154028 129464 154040
rect 129516 154028 129522 154080
rect 129550 154028 129556 154080
rect 129608 154068 129614 154080
rect 137296 154068 137324 154176
rect 146846 154136 146852 154148
rect 129608 154040 137324 154068
rect 137388 154108 146852 154136
rect 129608 154028 129614 154040
rect 7098 153960 7104 154012
rect 7156 154000 7162 154012
rect 118602 154000 118608 154012
rect 7156 153972 118608 154000
rect 7156 153960 7162 153972
rect 118602 153960 118608 153972
rect 118660 153960 118666 154012
rect 118694 153960 118700 154012
rect 118752 154000 118758 154012
rect 124306 154000 124312 154012
rect 118752 153972 120488 154000
rect 118752 153960 118758 153972
rect 1210 153892 1216 153944
rect 1268 153932 1274 153944
rect 119798 153932 119804 153944
rect 1268 153904 119804 153932
rect 1268 153892 1274 153904
rect 119798 153892 119804 153904
rect 119856 153892 119862 153944
rect 120460 153932 120488 153972
rect 120644 153972 124312 154000
rect 120644 153932 120672 153972
rect 124306 153960 124312 153972
rect 124364 153960 124370 154012
rect 124398 153960 124404 154012
rect 124456 154000 124462 154012
rect 124456 153972 127020 154000
rect 124456 153960 124462 153972
rect 120460 153904 120672 153932
rect 120718 153892 120724 153944
rect 120776 153932 120782 153944
rect 126882 153932 126888 153944
rect 120776 153904 126888 153932
rect 120776 153892 120782 153904
rect 126882 153892 126888 153904
rect 126940 153892 126946 153944
rect 126992 153932 127020 153972
rect 127802 153960 127808 154012
rect 127860 154000 127866 154012
rect 137388 154000 137416 154108
rect 146846 154096 146852 154108
rect 146904 154096 146910 154148
rect 137554 154028 137560 154080
rect 137612 154068 137618 154080
rect 146956 154068 146984 154244
rect 185210 154232 185216 154244
rect 185268 154232 185274 154284
rect 185302 154232 185308 154284
rect 185360 154272 185366 154284
rect 258534 154272 258540 154284
rect 185360 154244 258540 154272
rect 185360 154232 185366 154244
rect 258534 154232 258540 154244
rect 258592 154232 258598 154284
rect 266170 154232 266176 154284
rect 266228 154272 266234 154284
rect 322014 154272 322020 154284
rect 266228 154244 322020 154272
rect 266228 154232 266234 154244
rect 322014 154232 322020 154244
rect 322072 154232 322078 154284
rect 343542 154232 343548 154284
rect 343600 154272 343606 154284
rect 381170 154272 381176 154284
rect 343600 154244 381176 154272
rect 343600 154232 343606 154244
rect 381170 154232 381176 154244
rect 381228 154232 381234 154284
rect 393958 154232 393964 154284
rect 394016 154272 394022 154284
rect 419718 154272 419724 154284
rect 394016 154244 419724 154272
rect 394016 154232 394022 154244
rect 419718 154232 419724 154244
rect 419776 154232 419782 154284
rect 147122 154164 147128 154216
rect 147180 154204 147186 154216
rect 156598 154204 156604 154216
rect 147180 154176 156604 154204
rect 147180 154164 147186 154176
rect 156598 154164 156604 154176
rect 156656 154164 156662 154216
rect 156690 154164 156696 154216
rect 156748 154204 156754 154216
rect 163498 154204 163504 154216
rect 156748 154176 163504 154204
rect 156748 154164 156754 154176
rect 163498 154164 163504 154176
rect 163556 154164 163562 154216
rect 165062 154164 165068 154216
rect 165120 154204 165126 154216
rect 168650 154204 168656 154216
rect 165120 154176 168656 154204
rect 165120 154164 165126 154176
rect 168650 154164 168656 154176
rect 168708 154164 168714 154216
rect 172790 154164 172796 154216
rect 172848 154204 172854 154216
rect 250806 154204 250812 154216
rect 172848 154176 250812 154204
rect 172848 154164 172854 154176
rect 250806 154164 250812 154176
rect 250864 154164 250870 154216
rect 252646 154164 252652 154216
rect 252704 154204 252710 154216
rect 311710 154204 311716 154216
rect 252704 154176 311716 154204
rect 252704 154164 252710 154176
rect 311710 154164 311716 154176
rect 311768 154164 311774 154216
rect 326706 154164 326712 154216
rect 326764 154204 326770 154216
rect 368290 154204 368296 154216
rect 326764 154176 368296 154204
rect 326764 154164 326770 154176
rect 368290 154164 368296 154176
rect 368348 154164 368354 154216
rect 387610 154164 387616 154216
rect 387668 154204 387674 154216
rect 414566 154204 414572 154216
rect 387668 154176 414572 154204
rect 387668 154164 387674 154176
rect 414566 154164 414572 154176
rect 414624 154164 414630 154216
rect 147030 154096 147036 154148
rect 147088 154136 147094 154148
rect 153194 154136 153200 154148
rect 147088 154108 153200 154136
rect 147088 154096 147094 154108
rect 153194 154096 153200 154108
rect 153252 154096 153258 154148
rect 153378 154096 153384 154148
rect 153436 154136 153442 154148
rect 166258 154136 166264 154148
rect 153436 154108 166264 154136
rect 153436 154096 153442 154108
rect 166258 154096 166264 154108
rect 166316 154096 166322 154148
rect 166350 154096 166356 154148
rect 166408 154136 166414 154148
rect 245654 154136 245660 154148
rect 166408 154108 245660 154136
rect 166408 154096 166414 154108
rect 245654 154096 245660 154108
rect 245712 154096 245718 154148
rect 245930 154096 245936 154148
rect 245988 154136 245994 154148
rect 306650 154136 306656 154148
rect 245988 154108 306656 154136
rect 245988 154096 245994 154108
rect 306650 154096 306656 154108
rect 306708 154096 306714 154148
rect 323302 154096 323308 154148
rect 323360 154136 323366 154148
rect 365714 154136 365720 154148
rect 323360 154108 365720 154136
rect 323360 154096 323366 154108
rect 365714 154096 365720 154108
rect 365772 154096 365778 154148
rect 383930 154096 383936 154148
rect 383988 154136 383994 154148
rect 411990 154136 411996 154148
rect 383988 154108 411996 154136
rect 383988 154096 383994 154108
rect 411990 154096 411996 154108
rect 412048 154096 412054 154148
rect 137612 154040 146984 154068
rect 137612 154028 137618 154040
rect 152642 154028 152648 154080
rect 152700 154068 152706 154080
rect 235442 154068 235448 154080
rect 152700 154040 235448 154068
rect 152700 154028 152706 154040
rect 235442 154028 235448 154040
rect 235500 154028 235506 154080
rect 242618 154028 242624 154080
rect 242676 154068 242682 154080
rect 304074 154068 304080 154080
rect 242676 154040 304080 154068
rect 242676 154028 242682 154040
rect 304074 154028 304080 154040
rect 304132 154028 304138 154080
rect 319990 154028 319996 154080
rect 320048 154068 320054 154080
rect 363230 154068 363236 154080
rect 320048 154040 363236 154068
rect 320048 154028 320054 154040
rect 363230 154028 363236 154040
rect 363288 154028 363294 154080
rect 370406 154028 370412 154080
rect 370464 154068 370470 154080
rect 401686 154068 401692 154080
rect 370464 154040 401692 154068
rect 370464 154028 370470 154040
rect 401686 154028 401692 154040
rect 401744 154028 401750 154080
rect 127860 153972 137416 154000
rect 127860 153960 127866 153972
rect 137646 153960 137652 154012
rect 137704 154000 137710 154012
rect 142338 154000 142344 154012
rect 137704 153972 142344 154000
rect 137704 153960 137710 153972
rect 142338 153960 142344 153972
rect 142396 153960 142402 154012
rect 145098 153960 145104 154012
rect 145156 154000 145162 154012
rect 148134 154000 148140 154012
rect 145156 153972 148140 154000
rect 145156 153960 145162 153972
rect 148134 153960 148140 153972
rect 148192 153960 148198 154012
rect 150342 153960 150348 154012
rect 150400 154000 150406 154012
rect 233510 154000 233516 154012
rect 150400 153972 233516 154000
rect 150400 153960 150406 153972
rect 233510 153960 233516 153972
rect 233568 153960 233574 154012
rect 235902 153960 235908 154012
rect 235960 154000 235966 154012
rect 299014 154000 299020 154012
rect 235960 153972 299020 154000
rect 235960 153960 235966 153972
rect 299014 153960 299020 153972
rect 299072 153960 299078 154012
rect 313274 153960 313280 154012
rect 313332 154000 313338 154012
rect 357894 154000 357900 154012
rect 313332 153972 357900 154000
rect 313332 153960 313338 153972
rect 357894 153960 357900 153972
rect 357952 153960 357958 154012
rect 363690 153960 363696 154012
rect 363748 154000 363754 154012
rect 396534 154000 396540 154012
rect 363748 153972 396540 154000
rect 363748 153960 363754 153972
rect 396534 153960 396540 153972
rect 396592 153960 396598 154012
rect 397362 153960 397368 154012
rect 397420 154000 397426 154012
rect 422294 154000 422300 154012
rect 397420 153972 422300 154000
rect 397420 153960 397426 153972
rect 422294 153960 422300 153972
rect 422352 153960 422358 154012
rect 209774 153932 209780 153944
rect 126992 153904 209780 153932
rect 209774 153892 209780 153904
rect 209832 153892 209838 153944
rect 215662 153892 215668 153944
rect 215720 153932 215726 153944
rect 283650 153932 283656 153944
rect 215720 153904 283656 153932
rect 215720 153892 215726 153904
rect 283650 153892 283656 153904
rect 283708 153892 283714 153944
rect 284202 153892 284208 153944
rect 284260 153932 284266 153944
rect 334894 153932 334900 153944
rect 284260 153904 334900 153932
rect 284260 153892 284266 153904
rect 334894 153892 334900 153904
rect 334952 153892 334958 153944
rect 336826 153892 336832 153944
rect 336884 153932 336890 153944
rect 336884 153904 337608 153932
rect 336884 153892 336890 153904
rect 3970 153824 3976 153876
rect 4028 153864 4034 153876
rect 113818 153864 113824 153876
rect 4028 153836 113824 153864
rect 4028 153824 4034 153836
rect 113818 153824 113824 153836
rect 113876 153824 113882 153876
rect 115566 153824 115572 153876
rect 115624 153864 115630 153876
rect 118510 153864 118516 153876
rect 115624 153836 118516 153864
rect 115624 153824 115630 153836
rect 118510 153824 118516 153836
rect 118568 153824 118574 153876
rect 118602 153824 118608 153876
rect 118660 153864 118666 153876
rect 118694 153864 118700 153876
rect 118660 153836 118700 153864
rect 118660 153824 118666 153836
rect 118694 153824 118700 153836
rect 118752 153824 118758 153876
rect 125502 153824 125508 153876
rect 125560 153864 125566 153876
rect 129550 153864 129556 153876
rect 125560 153836 129556 153864
rect 125560 153824 125566 153836
rect 129550 153824 129556 153836
rect 129608 153824 129614 153876
rect 129918 153824 129924 153876
rect 129976 153864 129982 153876
rect 218054 153864 218060 153876
rect 129976 153836 218060 153864
rect 129976 153824 129982 153836
rect 218054 153824 218060 153836
rect 218112 153824 218118 153876
rect 219342 153824 219348 153876
rect 219400 153864 219406 153876
rect 286134 153864 286140 153876
rect 219400 153836 286140 153864
rect 219400 153824 219406 153836
rect 286134 153824 286140 153836
rect 286192 153824 286198 153876
rect 286318 153824 286324 153876
rect 286376 153864 286382 153876
rect 337470 153864 337476 153876
rect 286376 153836 337476 153864
rect 286376 153824 286382 153836
rect 337470 153824 337476 153836
rect 337528 153824 337534 153876
rect 337580 153864 337608 153904
rect 340138 153892 340144 153944
rect 340196 153932 340202 153944
rect 378594 153932 378600 153944
rect 340196 153904 378600 153932
rect 340196 153892 340202 153904
rect 378594 153892 378600 153904
rect 378652 153892 378658 153944
rect 380802 153892 380808 153944
rect 380860 153932 380866 153944
rect 409414 153932 409420 153944
rect 380860 153904 409420 153932
rect 380860 153892 380866 153904
rect 409414 153892 409420 153904
rect 409472 153892 409478 153944
rect 376018 153864 376024 153876
rect 337580 153836 376024 153864
rect 376018 153824 376024 153836
rect 376076 153824 376082 153876
rect 377214 153824 377220 153876
rect 377272 153864 377278 153876
rect 406838 153864 406844 153876
rect 377272 153836 406844 153864
rect 377272 153824 377278 153836
rect 406838 153824 406844 153836
rect 406896 153824 406902 153876
rect 48314 153756 48320 153808
rect 48372 153796 48378 153808
rect 155770 153796 155776 153808
rect 48372 153768 155776 153796
rect 48372 153756 48378 153768
rect 155770 153756 155776 153768
rect 155828 153756 155834 153808
rect 156598 153756 156604 153808
rect 156656 153796 156662 153808
rect 212902 153796 212908 153808
rect 156656 153768 212908 153796
rect 156656 153756 156662 153768
rect 212902 153756 212908 153768
rect 212960 153756 212966 153808
rect 222378 153756 222384 153808
rect 222436 153796 222442 153808
rect 288710 153796 288716 153808
rect 222436 153768 288716 153796
rect 222436 153756 222442 153768
rect 288710 153756 288716 153768
rect 288768 153756 288774 153808
rect 360378 153756 360384 153808
rect 360436 153796 360442 153808
rect 394050 153796 394056 153808
rect 360436 153768 394056 153796
rect 360436 153756 360442 153768
rect 394050 153756 394056 153768
rect 394108 153756 394114 153808
rect 58342 153688 58348 153740
rect 58400 153728 58406 153740
rect 156690 153728 156696 153740
rect 58400 153700 156696 153728
rect 58400 153688 58406 153700
rect 156690 153688 156696 153700
rect 156748 153688 156754 153740
rect 156782 153688 156788 153740
rect 156840 153728 156846 153740
rect 210418 153728 210424 153740
rect 156840 153700 210424 153728
rect 156840 153688 156846 153700
rect 210418 153688 210424 153700
rect 210476 153688 210482 153740
rect 229094 153688 229100 153740
rect 229152 153728 229158 153740
rect 293862 153728 293868 153740
rect 229152 153700 293868 153728
rect 229152 153688 229158 153700
rect 293862 153688 293868 153700
rect 293920 153688 293926 153740
rect 65150 153620 65156 153672
rect 65208 153660 65214 153672
rect 165062 153660 165068 153672
rect 65208 153632 165068 153660
rect 65208 153620 65214 153632
rect 165062 153620 165068 153632
rect 165120 153620 165126 153672
rect 166258 153620 166264 153672
rect 166316 153660 166322 153672
rect 215478 153660 215484 153672
rect 166316 153632 215484 153660
rect 166316 153620 166322 153632
rect 215478 153620 215484 153632
rect 215536 153620 215542 153672
rect 239214 153620 239220 153672
rect 239272 153660 239278 153672
rect 301590 153660 301596 153672
rect 239272 153632 301596 153660
rect 239272 153620 239278 153632
rect 301590 153620 301596 153632
rect 301648 153620 301654 153672
rect 82814 153552 82820 153604
rect 82872 153592 82878 153604
rect 182082 153592 182088 153604
rect 82872 153564 182088 153592
rect 82872 153552 82878 153564
rect 182082 153552 182088 153564
rect 182140 153552 182146 153604
rect 182910 153552 182916 153604
rect 182968 153592 182974 153604
rect 185026 153592 185032 153604
rect 182968 153564 185032 153592
rect 182968 153552 182974 153564
rect 185026 153552 185032 153564
rect 185084 153552 185090 153604
rect 185118 153552 185124 153604
rect 185176 153592 185182 153604
rect 188338 153592 188344 153604
rect 185176 153564 188344 153592
rect 185176 153552 185182 153564
rect 188338 153552 188344 153564
rect 188396 153552 188402 153604
rect 188430 153552 188436 153604
rect 188488 153592 188494 153604
rect 197538 153592 197544 153604
rect 188488 153564 197544 153592
rect 188488 153552 188494 153564
rect 197538 153552 197544 153564
rect 197596 153552 197602 153604
rect 198918 153552 198924 153604
rect 198976 153592 198982 153604
rect 248874 153592 248880 153604
rect 198976 153564 248880 153592
rect 198976 153552 198982 153564
rect 248874 153552 248880 153564
rect 248932 153552 248938 153604
rect 249702 153552 249708 153604
rect 249760 153592 249766 153604
rect 309226 153592 309232 153604
rect 249760 153564 309232 153592
rect 249760 153552 249766 153564
rect 309226 153552 309232 153564
rect 309284 153552 309290 153604
rect 102134 153484 102140 153536
rect 102192 153524 102198 153536
rect 196894 153524 196900 153536
rect 102192 153496 196900 153524
rect 102192 153484 102198 153496
rect 196894 153484 196900 153496
rect 196952 153484 196958 153536
rect 196986 153484 196992 153536
rect 197044 153524 197050 153536
rect 199378 153524 199384 153536
rect 197044 153496 199384 153524
rect 197044 153484 197050 153496
rect 199378 153484 199384 153496
rect 199436 153484 199442 153536
rect 199488 153496 200114 153524
rect 108850 153416 108856 153468
rect 108908 153456 108914 153468
rect 191374 153456 191380 153468
rect 108908 153428 191380 153456
rect 108908 153416 108914 153428
rect 191374 153416 191380 153428
rect 191432 153416 191438 153468
rect 194502 153416 194508 153468
rect 194560 153456 194566 153468
rect 199488 153456 199516 153496
rect 194560 153428 199516 153456
rect 200086 153456 200114 153496
rect 200390 153484 200396 153536
rect 200448 153524 200454 153536
rect 256510 153524 256516 153536
rect 200448 153496 256516 153524
rect 200448 153484 200454 153496
rect 256510 153484 256516 153496
rect 256568 153484 256574 153536
rect 314378 153524 314384 153536
rect 258046 153496 314384 153524
rect 238662 153456 238668 153468
rect 200086 153428 238668 153456
rect 194560 153416 194566 153428
rect 238662 153416 238668 153428
rect 238720 153416 238726 153468
rect 105446 153348 105452 153400
rect 105504 153388 105510 153400
rect 199470 153388 199476 153400
rect 105504 153360 199476 153388
rect 105504 153348 105510 153360
rect 199470 153348 199476 153360
rect 199528 153348 199534 153400
rect 199562 153348 199568 153400
rect 199620 153388 199626 153400
rect 243722 153388 243728 153400
rect 199620 153360 243728 153388
rect 199620 153348 199626 153360
rect 243722 153348 243728 153360
rect 243780 153348 243786 153400
rect 256050 153348 256056 153400
rect 256108 153388 256114 153400
rect 258046 153388 258074 153496
rect 314378 153484 314384 153496
rect 314436 153484 314442 153536
rect 262766 153416 262772 153468
rect 262824 153456 262830 153468
rect 319530 153456 319536 153468
rect 262824 153428 319536 153456
rect 262824 153416 262830 153428
rect 319530 153416 319536 153428
rect 319588 153416 319594 153468
rect 256108 153360 258074 153388
rect 256108 153348 256114 153360
rect 259546 153348 259552 153400
rect 259604 153388 259610 153400
rect 316954 153388 316960 153400
rect 259604 153360 316960 153388
rect 259604 153348 259610 153360
rect 316954 153348 316960 153360
rect 317012 153348 317018 153400
rect 113818 153280 113824 153332
rect 113876 153320 113882 153332
rect 118418 153320 118424 153332
rect 113876 153292 118424 153320
rect 113876 153280 113882 153292
rect 118418 153280 118424 153292
rect 118476 153280 118482 153332
rect 120718 153280 120724 153332
rect 120776 153320 120782 153332
rect 207198 153320 207204 153332
rect 120776 153292 207204 153320
rect 120776 153280 120782 153292
rect 207198 153280 207204 153292
rect 207256 153280 207262 153332
rect 272886 153280 272892 153332
rect 272944 153320 272950 153332
rect 327258 153320 327264 153332
rect 272944 153292 327264 153320
rect 272944 153280 272950 153292
rect 327258 153280 327264 153292
rect 327316 153280 327322 153332
rect 119430 153212 119436 153264
rect 119488 153252 119494 153264
rect 207842 153252 207848 153264
rect 119488 153224 207848 153252
rect 119488 153212 119494 153224
rect 207842 153212 207848 153224
rect 207900 153212 207906 153264
rect 269482 153212 269488 153264
rect 269540 153252 269546 153264
rect 324682 153252 324688 153264
rect 269540 153224 324688 153252
rect 269540 153212 269546 153224
rect 324682 153212 324688 153224
rect 324740 153212 324746 153264
rect 433058 153252 433064 153264
rect 432340 153224 433064 153252
rect 118510 153144 118516 153196
rect 118568 153184 118574 153196
rect 120718 153184 120724 153196
rect 118568 153156 120724 153184
rect 118568 153144 118574 153156
rect 120718 153144 120724 153156
rect 120776 153144 120782 153196
rect 123478 153144 123484 153196
rect 123536 153184 123542 153196
rect 205910 153184 205916 153196
rect 123536 153156 205916 153184
rect 123536 153144 123542 153156
rect 205910 153144 205916 153156
rect 205968 153144 205974 153196
rect 225046 153144 225052 153196
rect 225104 153184 225110 153196
rect 229002 153184 229008 153196
rect 225104 153156 229008 153184
rect 225104 153144 225110 153156
rect 229002 153144 229008 153156
rect 229060 153144 229066 153196
rect 234430 153144 234436 153196
rect 234488 153184 234494 153196
rect 297726 153184 297732 153196
rect 234488 153156 297732 153184
rect 234488 153144 234494 153156
rect 297726 153144 297732 153156
rect 297784 153144 297790 153196
rect 300302 153144 300308 153196
rect 300360 153184 300366 153196
rect 342254 153184 342260 153196
rect 300360 153156 342260 153184
rect 300360 153144 300366 153156
rect 342254 153144 342260 153156
rect 342312 153144 342318 153196
rect 342346 153144 342352 153196
rect 342404 153184 342410 153196
rect 343910 153184 343916 153196
rect 342404 153156 343916 153184
rect 342404 153144 342410 153156
rect 343910 153144 343916 153156
rect 343968 153144 343974 153196
rect 345290 153144 345296 153196
rect 345348 153184 345354 153196
rect 345750 153184 345756 153196
rect 345348 153156 345756 153184
rect 345348 153144 345354 153156
rect 345750 153144 345756 153156
rect 345808 153144 345814 153196
rect 349430 153144 349436 153196
rect 349488 153184 349494 153196
rect 385586 153184 385592 153196
rect 349488 153156 385592 153184
rect 349488 153144 349494 153156
rect 385586 153144 385592 153156
rect 385644 153144 385650 153196
rect 390370 153144 390376 153196
rect 390428 153184 390434 153196
rect 415210 153184 415216 153196
rect 390428 153156 415216 153184
rect 390428 153144 390434 153156
rect 415210 153144 415216 153156
rect 415268 153144 415274 153196
rect 415854 153144 415860 153196
rect 415912 153184 415918 153196
rect 432340 153184 432368 153224
rect 433058 153212 433064 153224
rect 433116 153212 433122 153264
rect 435726 153184 435732 153196
rect 415912 153156 432368 153184
rect 432432 153156 435732 153184
rect 415912 153144 415918 153156
rect 103790 153076 103796 153128
rect 103848 153116 103854 153128
rect 198182 153116 198188 153128
rect 103848 153088 198188 153116
rect 103848 153076 103854 153088
rect 198182 153076 198188 153088
rect 198240 153076 198246 153128
rect 215294 153076 215300 153128
rect 215352 153116 215358 153128
rect 279694 153116 279700 153128
rect 215352 153088 279700 153116
rect 215352 153076 215358 153088
rect 279694 153076 279700 153088
rect 279752 153076 279758 153128
rect 279878 153076 279884 153128
rect 279936 153116 279942 153128
rect 331766 153116 331772 153128
rect 279936 153088 331772 153116
rect 279936 153076 279942 153088
rect 331766 153076 331772 153088
rect 331824 153076 331830 153128
rect 332594 153076 332600 153128
rect 332652 153116 332658 153128
rect 372798 153116 372804 153128
rect 332652 153088 372804 153116
rect 332652 153076 332658 153088
rect 372798 153076 372804 153088
rect 372856 153076 372862 153128
rect 372982 153076 372988 153128
rect 373040 153116 373046 153128
rect 403618 153116 403624 153128
rect 373040 153088 403624 153116
rect 373040 153076 373046 153088
rect 403618 153076 403624 153088
rect 403676 153076 403682 153128
rect 408494 153076 408500 153128
rect 408552 153116 408558 153128
rect 415118 153116 415124 153128
rect 408552 153088 415124 153116
rect 408552 153076 408558 153088
rect 415118 153076 415124 153088
rect 415176 153076 415182 153128
rect 415302 153076 415308 153128
rect 415360 153116 415366 153128
rect 432432 153116 432460 153156
rect 435726 153144 435732 153156
rect 435784 153144 435790 153196
rect 435818 153144 435824 153196
rect 435876 153184 435882 153196
rect 435876 153156 436508 153184
rect 435876 153144 435882 153156
rect 433150 153116 433156 153128
rect 415360 153088 432460 153116
rect 432524 153088 433156 153116
rect 415360 153076 415366 153088
rect 86862 153008 86868 153060
rect 86920 153048 86926 153060
rect 180242 153048 180248 153060
rect 86920 153020 180248 153048
rect 86920 153008 86926 153020
rect 180242 153008 180248 153020
rect 180300 153008 180306 153060
rect 181162 153008 181168 153060
rect 181220 153048 181226 153060
rect 257246 153048 257252 153060
rect 181220 153020 257252 153048
rect 181220 153008 181226 153020
rect 257246 153008 257252 153020
rect 257304 153008 257310 153060
rect 257706 153008 257712 153060
rect 257764 153048 257770 153060
rect 315666 153048 315672 153060
rect 257764 153020 315672 153048
rect 257764 153008 257770 153020
rect 315666 153008 315672 153020
rect 315724 153008 315730 153060
rect 317138 153008 317144 153060
rect 317196 153048 317202 153060
rect 318242 153048 318248 153060
rect 317196 153020 318248 153048
rect 317196 153008 317202 153020
rect 318242 153008 318248 153020
rect 318300 153008 318306 153060
rect 318426 153008 318432 153060
rect 318484 153048 318490 153060
rect 361298 153048 361304 153060
rect 318484 153020 361304 153048
rect 318484 153008 318490 153020
rect 361298 153008 361304 153020
rect 361356 153008 361362 153060
rect 367186 153008 367192 153060
rect 367244 153048 367250 153060
rect 368934 153048 368940 153060
rect 367244 153020 368940 153048
rect 367244 153008 367250 153020
rect 368934 153008 368940 153020
rect 368992 153008 368998 153060
rect 369026 153008 369032 153060
rect 369084 153048 369090 153060
rect 397178 153048 397184 153060
rect 369084 153020 397184 153048
rect 369084 153008 369090 153020
rect 397178 153008 397184 153020
rect 397236 153008 397242 153060
rect 398098 153008 398104 153060
rect 398156 153048 398162 153060
rect 408126 153048 408132 153060
rect 398156 153020 408132 153048
rect 398156 153008 398162 153020
rect 408126 153008 408132 153020
rect 408184 153008 408190 153060
rect 411622 153008 411628 153060
rect 411680 153048 411686 153060
rect 432524 153048 432552 153088
rect 433150 153076 433156 153088
rect 433208 153076 433214 153128
rect 433242 153076 433248 153128
rect 433300 153116 433306 153128
rect 436370 153116 436376 153128
rect 433300 153088 436376 153116
rect 433300 153076 433306 153088
rect 436370 153076 436376 153088
rect 436428 153076 436434 153128
rect 436480 153116 436508 153156
rect 437290 153144 437296 153196
rect 437348 153184 437354 153196
rect 452470 153184 452476 153196
rect 437348 153156 452476 153184
rect 437348 153144 437354 153156
rect 452470 153144 452476 153156
rect 452528 153144 452534 153196
rect 453942 153144 453948 153196
rect 454000 153184 454006 153196
rect 459462 153184 459468 153196
rect 454000 153156 459468 153184
rect 454000 153144 454006 153156
rect 459462 153144 459468 153156
rect 459520 153144 459526 153196
rect 461854 153144 461860 153196
rect 461912 153184 461918 153196
rect 465902 153184 465908 153196
rect 461912 153156 465908 153184
rect 461912 153144 461918 153156
rect 465902 153144 465908 153156
rect 465960 153144 465966 153196
rect 466454 153144 466460 153196
rect 466512 153184 466518 153196
rect 469766 153184 469772 153196
rect 466512 153156 469772 153184
rect 466512 153144 466518 153156
rect 469766 153144 469772 153156
rect 469824 153144 469830 153196
rect 471238 153144 471244 153196
rect 471296 153184 471302 153196
rect 472986 153184 472992 153196
rect 471296 153156 472992 153184
rect 471296 153144 471302 153156
rect 472986 153144 472992 153156
rect 473044 153144 473050 153196
rect 474826 153144 474832 153196
rect 474884 153184 474890 153196
rect 476850 153184 476856 153196
rect 474884 153156 476856 153184
rect 474884 153144 474890 153156
rect 476850 153144 476856 153156
rect 476908 153144 476914 153196
rect 485682 153144 485688 153196
rect 485740 153184 485746 153196
rect 489638 153184 489644 153196
rect 485740 153156 489644 153184
rect 485740 153144 485746 153156
rect 489638 153144 489644 153156
rect 489696 153144 489702 153196
rect 490742 153144 490748 153196
rect 490800 153184 490806 153196
rect 493502 153184 493508 153196
rect 490800 153156 493508 153184
rect 490800 153144 490806 153156
rect 493502 153144 493508 153156
rect 493560 153144 493566 153196
rect 494054 153144 494060 153196
rect 494112 153184 494118 153196
rect 496078 153184 496084 153196
rect 494112 153156 496084 153184
rect 494112 153144 494118 153156
rect 496078 153144 496084 153156
rect 496136 153144 496142 153196
rect 496630 153144 496636 153196
rect 496688 153184 496694 153196
rect 498010 153184 498016 153196
rect 496688 153156 498016 153184
rect 496688 153144 496694 153156
rect 498010 153144 498016 153156
rect 498068 153144 498074 153196
rect 498286 153144 498292 153196
rect 498344 153184 498350 153196
rect 499298 153184 499304 153196
rect 498344 153156 499304 153184
rect 498344 153144 498350 153156
rect 499298 153144 499304 153156
rect 499356 153144 499362 153196
rect 500954 153144 500960 153196
rect 501012 153184 501018 153196
rect 501874 153184 501880 153196
rect 501012 153156 501880 153184
rect 501012 153144 501018 153156
rect 501874 153144 501880 153156
rect 501932 153144 501938 153196
rect 511626 153144 511632 153196
rect 511684 153184 511690 153196
rect 513742 153184 513748 153196
rect 511684 153156 513748 153184
rect 511684 153144 511690 153156
rect 513742 153144 513748 153156
rect 513800 153144 513806 153196
rect 514202 153144 514208 153196
rect 514260 153184 514266 153196
rect 517422 153184 517428 153196
rect 514260 153156 517428 153184
rect 514260 153144 514266 153156
rect 517422 153144 517428 153156
rect 517480 153144 517486 153196
rect 438486 153116 438492 153128
rect 436480 153088 438492 153116
rect 438486 153076 438492 153088
rect 438544 153076 438550 153128
rect 438578 153076 438584 153128
rect 438636 153116 438642 153128
rect 453758 153116 453764 153128
rect 438636 153088 453764 153116
rect 438636 153076 438642 153088
rect 453758 153076 453764 153088
rect 453816 153076 453822 153128
rect 456886 153076 456892 153128
rect 456944 153116 456950 153128
rect 460750 153116 460756 153128
rect 456944 153088 460756 153116
rect 456944 153076 456950 153088
rect 460750 153076 460756 153088
rect 460808 153076 460814 153128
rect 462958 153076 462964 153128
rect 463016 153116 463022 153128
rect 467190 153116 467196 153128
rect 463016 153088 467196 153116
rect 463016 153076 463022 153088
rect 467190 153076 467196 153088
rect 467248 153076 467254 153128
rect 471606 153076 471612 153128
rect 471664 153116 471670 153128
rect 473630 153116 473636 153128
rect 471664 153088 473636 153116
rect 471664 153076 471670 153088
rect 473630 153076 473636 153088
rect 473688 153076 473694 153128
rect 476114 153076 476120 153128
rect 476172 153116 476178 153128
rect 478138 153116 478144 153128
rect 476172 153088 478144 153116
rect 476172 153076 476178 153088
rect 478138 153076 478144 153088
rect 478196 153076 478202 153128
rect 484854 153076 484860 153128
rect 484912 153116 484918 153128
rect 488994 153116 489000 153128
rect 484912 153088 489000 153116
rect 484912 153076 484918 153088
rect 488994 153076 489000 153088
rect 489052 153076 489058 153128
rect 489914 153076 489920 153128
rect 489972 153116 489978 153128
rect 492858 153116 492864 153128
rect 489972 153088 492864 153116
rect 489972 153076 489978 153088
rect 492858 153076 492864 153088
rect 492916 153076 492922 153128
rect 493226 153076 493232 153128
rect 493284 153116 493290 153128
rect 495434 153116 495440 153128
rect 493284 153088 495440 153116
rect 493284 153076 493290 153088
rect 495434 153076 495440 153088
rect 495492 153076 495498 153128
rect 495802 153076 495808 153128
rect 495860 153116 495866 153128
rect 497366 153116 497372 153128
rect 495860 153088 497372 153116
rect 495860 153076 495866 153088
rect 497366 153076 497372 153088
rect 497424 153076 497430 153128
rect 497458 153076 497464 153128
rect 497516 153116 497522 153128
rect 498654 153116 498660 153128
rect 497516 153088 498660 153116
rect 497516 153076 497522 153088
rect 498654 153076 498660 153088
rect 498712 153076 498718 153128
rect 510982 153076 510988 153128
rect 511040 153116 511046 153128
rect 513466 153116 513472 153128
rect 511040 153088 513472 153116
rect 511040 153076 511046 153088
rect 513466 153076 513472 153088
rect 513524 153076 513530 153128
rect 513558 153076 513564 153128
rect 513616 153116 513622 153128
rect 516134 153116 516140 153128
rect 513616 153088 516140 153116
rect 513616 153076 513622 153088
rect 516134 153076 516140 153088
rect 516192 153076 516198 153128
rect 411680 153020 432552 153048
rect 411680 153008 411686 153020
rect 432690 153008 432696 153060
rect 432748 153048 432754 153060
rect 449250 153048 449256 153060
rect 432748 153020 449256 153048
rect 432748 153008 432754 153020
rect 449250 153008 449256 153020
rect 449308 153008 449314 153060
rect 463326 153008 463332 153060
rect 463384 153048 463390 153060
rect 466546 153048 466552 153060
rect 463384 153020 466552 153048
rect 463384 153008 463390 153020
rect 466546 153008 466552 153020
rect 466604 153008 466610 153060
rect 466638 153008 466644 153060
rect 466696 153048 466702 153060
rect 470410 153048 470416 153060
rect 466696 153020 470416 153048
rect 466696 153008 466702 153020
rect 470410 153008 470416 153020
rect 470468 153008 470474 153060
rect 472434 153008 472440 153060
rect 472492 153048 472498 153060
rect 474274 153048 474280 153060
rect 472492 153020 474280 153048
rect 472492 153008 472498 153020
rect 474274 153008 474280 153020
rect 474332 153008 474338 153060
rect 484026 153008 484032 153060
rect 484084 153048 484090 153060
rect 488350 153048 488356 153060
rect 484084 153020 488356 153048
rect 484084 153008 484090 153020
rect 488350 153008 488356 153020
rect 488408 153008 488414 153060
rect 492398 153008 492404 153060
rect 492456 153048 492462 153060
rect 494790 153048 494796 153060
rect 492456 153020 494796 153048
rect 492456 153008 492462 153020
rect 494790 153008 494796 153020
rect 494848 153008 494854 153060
rect 495250 153008 495256 153060
rect 495308 153048 495314 153060
rect 496630 153048 496636 153060
rect 495308 153020 496636 153048
rect 495308 153008 495314 153020
rect 496630 153008 496636 153020
rect 496688 153008 496694 153060
rect 512270 153008 512276 153060
rect 512328 153048 512334 153060
rect 514846 153048 514852 153060
rect 512328 153020 514852 153048
rect 512328 153008 512334 153020
rect 514846 153008 514852 153020
rect 514904 153008 514910 153060
rect 97074 152940 97080 152992
rect 97132 152980 97138 152992
rect 193030 152980 193036 152992
rect 97132 152952 193036 152980
rect 97132 152940 97138 152952
rect 193030 152940 193036 152952
rect 193088 152940 193094 152992
rect 203702 152940 203708 152992
rect 203760 152980 203766 152992
rect 267550 152980 267556 152992
rect 203760 152952 267556 152980
rect 203760 152940 203766 152952
rect 267550 152940 267556 152952
rect 267608 152940 267614 152992
rect 267642 152940 267648 152992
rect 267700 152980 267706 152992
rect 320910 152980 320916 152992
rect 267700 152952 320916 152980
rect 267700 152940 267706 152952
rect 320910 152940 320916 152952
rect 320968 152940 320974 152992
rect 325878 152940 325884 152992
rect 325936 152980 325942 152992
rect 367646 152980 367652 152992
rect 325936 152952 367652 152980
rect 325936 152940 325942 152952
rect 367646 152940 367652 152952
rect 367704 152940 367710 152992
rect 368750 152940 368756 152992
rect 368808 152980 368814 152992
rect 400398 152980 400404 152992
rect 368808 152952 400404 152980
rect 368808 152940 368814 152952
rect 400398 152940 400404 152952
rect 400456 152940 400462 152992
rect 407022 152940 407028 152992
rect 407080 152980 407086 152992
rect 429194 152980 429200 152992
rect 407080 152952 429200 152980
rect 407080 152940 407086 152952
rect 429194 152940 429200 152952
rect 429252 152940 429258 152992
rect 429286 152940 429292 152992
rect 429344 152980 429350 152992
rect 446674 152980 446680 152992
rect 429344 152952 446680 152980
rect 429344 152940 429350 152952
rect 446674 152940 446680 152952
rect 446732 152940 446738 152992
rect 459554 152940 459560 152992
rect 459612 152980 459618 152992
rect 464614 152980 464620 152992
rect 459612 152952 464620 152980
rect 459612 152940 459618 152952
rect 464614 152940 464620 152952
rect 464672 152940 464678 152992
rect 465074 152940 465080 152992
rect 465132 152980 465138 152992
rect 469122 152980 469128 152992
rect 465132 152952 469128 152980
rect 465132 152940 465138 152952
rect 469122 152940 469128 152952
rect 469180 152940 469186 152992
rect 472526 152940 472532 152992
rect 472584 152980 472590 152992
rect 474918 152980 474924 152992
rect 472584 152952 474924 152980
rect 472584 152940 472590 152952
rect 474918 152940 474924 152952
rect 474976 152940 474982 152992
rect 483198 152940 483204 152992
rect 483256 152980 483262 152992
rect 487798 152980 487804 152992
rect 483256 152952 487804 152980
rect 483256 152940 483262 152952
rect 487798 152940 487804 152952
rect 487856 152940 487862 152992
rect 491570 152940 491576 152992
rect 491628 152980 491634 152992
rect 494146 152980 494152 152992
rect 491628 152952 494152 152980
rect 491628 152940 491634 152952
rect 494146 152940 494152 152952
rect 494204 152940 494210 152992
rect 512914 152940 512920 152992
rect 512972 152980 512978 152992
rect 515950 152980 515956 152992
rect 512972 152952 515956 152980
rect 512972 152940 512978 152952
rect 515950 152940 515956 152952
rect 516008 152940 516014 152992
rect 90358 152872 90364 152924
rect 90416 152912 90422 152924
rect 187878 152912 187884 152924
rect 90416 152884 187884 152912
rect 90416 152872 90422 152884
rect 187878 152872 187884 152884
rect 187936 152872 187942 152924
rect 187970 152872 187976 152924
rect 188028 152912 188034 152924
rect 262398 152912 262404 152924
rect 188028 152884 262404 152912
rect 188028 152872 188034 152884
rect 262398 152872 262404 152884
rect 262456 152872 262462 152924
rect 270862 152872 270868 152924
rect 270920 152912 270926 152924
rect 321462 152912 321468 152924
rect 270920 152884 321468 152912
rect 270920 152872 270926 152884
rect 321462 152872 321468 152884
rect 321520 152872 321526 152924
rect 321554 152872 321560 152924
rect 321612 152912 321618 152924
rect 323486 152912 323492 152924
rect 321612 152884 323492 152912
rect 321612 152872 321618 152884
rect 323486 152872 323492 152884
rect 323544 152872 323550 152924
rect 324222 152872 324228 152924
rect 324280 152912 324286 152924
rect 366358 152912 366364 152924
rect 324280 152884 366364 152912
rect 324280 152872 324286 152884
rect 366358 152872 366364 152884
rect 366416 152872 366422 152924
rect 366450 152872 366456 152924
rect 366508 152912 366514 152924
rect 398466 152912 398472 152924
rect 366508 152884 398472 152912
rect 366508 152872 366514 152884
rect 398466 152872 398472 152884
rect 398524 152872 398530 152924
rect 402422 152872 402428 152924
rect 402480 152912 402486 152924
rect 426158 152912 426164 152924
rect 402480 152884 426164 152912
rect 402480 152872 402486 152884
rect 426158 152872 426164 152884
rect 426216 152872 426222 152924
rect 426250 152872 426256 152924
rect 426308 152912 426314 152924
rect 427170 152912 427176 152924
rect 426308 152884 427176 152912
rect 426308 152872 426314 152884
rect 427170 152872 427176 152884
rect 427228 152872 427234 152924
rect 430482 152872 430488 152924
rect 430540 152912 430546 152924
rect 447318 152912 447324 152924
rect 430540 152884 447324 152912
rect 430540 152872 430546 152884
rect 447318 152872 447324 152884
rect 447376 152872 447382 152924
rect 464154 152872 464160 152924
rect 464212 152912 464218 152924
rect 467834 152912 467840 152924
rect 464212 152884 467840 152912
rect 464212 152872 464218 152884
rect 467834 152872 467840 152884
rect 467892 152872 467898 152924
rect 473354 152872 473360 152924
rect 473412 152912 473418 152924
rect 475562 152912 475568 152924
rect 473412 152884 475568 152912
rect 473412 152872 473418 152884
rect 475562 152872 475568 152884
rect 475620 152872 475626 152924
rect 66806 152804 66812 152856
rect 66864 152844 66870 152856
rect 169938 152844 169944 152856
rect 66864 152816 169944 152844
rect 66864 152804 66870 152816
rect 169938 152804 169944 152816
rect 169996 152804 170002 152856
rect 174538 152804 174544 152856
rect 174596 152844 174602 152856
rect 252094 152844 252100 152856
rect 174596 152816 252100 152844
rect 174596 152804 174602 152816
rect 252094 152804 252100 152816
rect 252152 152804 252158 152856
rect 252186 152804 252192 152856
rect 252244 152844 252250 152856
rect 311158 152844 311164 152856
rect 252244 152816 311164 152844
rect 252244 152804 252250 152816
rect 311158 152804 311164 152816
rect 311216 152804 311222 152856
rect 318702 152804 318708 152856
rect 318760 152844 318766 152856
rect 361942 152844 361948 152856
rect 318760 152816 361948 152844
rect 318760 152804 318766 152816
rect 361942 152804 361948 152816
rect 362000 152804 362006 152856
rect 362034 152804 362040 152856
rect 362092 152844 362098 152856
rect 395430 152844 395436 152856
rect 362092 152816 395436 152844
rect 362092 152804 362098 152816
rect 395430 152804 395436 152816
rect 395488 152804 395494 152856
rect 395522 152804 395528 152856
rect 395580 152844 395586 152856
rect 397822 152844 397828 152856
rect 395580 152816 397828 152844
rect 395580 152804 395586 152816
rect 397822 152804 397828 152816
rect 397880 152804 397886 152856
rect 400122 152804 400128 152856
rect 400180 152844 400186 152856
rect 424226 152844 424232 152856
rect 400180 152816 424232 152844
rect 400180 152804 400186 152816
rect 424226 152804 424232 152816
rect 424284 152804 424290 152856
rect 425146 152804 425152 152856
rect 425204 152844 425210 152856
rect 443454 152844 443460 152856
rect 425204 152816 443460 152844
rect 425204 152804 425210 152816
rect 443454 152804 443460 152816
rect 443512 152804 443518 152856
rect 444466 152804 444472 152856
rect 444524 152844 444530 152856
rect 458266 152844 458272 152856
rect 444524 152816 458272 152844
rect 444524 152804 444530 152816
rect 458266 152804 458272 152816
rect 458324 152804 458330 152856
rect 464522 152804 464528 152856
rect 464580 152844 464586 152856
rect 468386 152844 468392 152856
rect 464580 152816 468392 152844
rect 464580 152804 464586 152816
rect 468386 152804 468392 152816
rect 468444 152804 468450 152856
rect 510338 152804 510344 152856
rect 510396 152844 510402 152856
rect 511994 152844 512000 152856
rect 510396 152816 512000 152844
rect 510396 152804 510402 152816
rect 511994 152804 512000 152816
rect 512052 152804 512058 152856
rect 26418 152736 26424 152788
rect 26476 152776 26482 152788
rect 139118 152776 139124 152788
rect 26476 152748 139124 152776
rect 26476 152736 26482 152748
rect 139118 152736 139124 152748
rect 139176 152736 139182 152788
rect 143534 152776 143540 152788
rect 139228 152748 143540 152776
rect 22186 152668 22192 152720
rect 22244 152708 22250 152720
rect 135898 152708 135904 152720
rect 22244 152680 135904 152708
rect 22244 152668 22250 152680
rect 135898 152668 135904 152680
rect 135956 152668 135962 152720
rect 137462 152668 137468 152720
rect 137520 152708 137526 152720
rect 139228 152708 139256 152748
rect 143534 152736 143540 152748
rect 143592 152736 143598 152788
rect 151906 152776 151912 152788
rect 143736 152748 151912 152776
rect 137520 152680 139256 152708
rect 137520 152668 137526 152680
rect 139394 152668 139400 152720
rect 139452 152708 139458 152720
rect 141694 152708 141700 152720
rect 139452 152680 141700 152708
rect 139452 152668 139458 152680
rect 141694 152668 141700 152680
rect 141752 152668 141758 152720
rect 141786 152668 141792 152720
rect 141844 152708 141850 152720
rect 143736 152708 143764 152748
rect 151906 152736 151912 152748
rect 151964 152736 151970 152788
rect 154298 152736 154304 152788
rect 154356 152776 154362 152788
rect 236730 152776 236736 152788
rect 154356 152748 236736 152776
rect 154356 152736 154362 152748
rect 236730 152736 236736 152748
rect 236788 152736 236794 152788
rect 240318 152736 240324 152788
rect 240376 152776 240382 152788
rect 241882 152776 241888 152788
rect 240376 152748 241888 152776
rect 240376 152736 240382 152748
rect 241882 152736 241888 152748
rect 241940 152736 241946 152788
rect 247678 152736 247684 152788
rect 247736 152776 247742 152788
rect 307938 152776 307944 152788
rect 247736 152748 307944 152776
rect 247736 152736 247742 152748
rect 307938 152736 307944 152748
rect 307996 152736 308002 152788
rect 311802 152736 311808 152788
rect 311860 152776 311866 152788
rect 356790 152776 356796 152788
rect 311860 152748 356796 152776
rect 311860 152736 311866 152748
rect 356790 152736 356796 152748
rect 356848 152736 356854 152788
rect 357434 152736 357440 152788
rect 357492 152776 357498 152788
rect 359366 152776 359372 152788
rect 357492 152748 359372 152776
rect 357492 152736 357498 152748
rect 359366 152736 359372 152748
rect 359424 152736 359430 152788
rect 359550 152736 359556 152788
rect 359608 152776 359614 152788
rect 393406 152776 393412 152788
rect 359608 152748 393412 152776
rect 359608 152736 359614 152748
rect 393406 152736 393412 152748
rect 393464 152736 393470 152788
rect 394878 152736 394884 152788
rect 394936 152776 394942 152788
rect 420362 152776 420368 152788
rect 394936 152748 420368 152776
rect 394936 152736 394942 152748
rect 420362 152736 420368 152748
rect 420420 152736 420426 152788
rect 421742 152736 421748 152788
rect 421800 152776 421806 152788
rect 433334 152776 433340 152788
rect 421800 152748 433340 152776
rect 421800 152736 421806 152748
rect 433334 152736 433340 152748
rect 433392 152736 433398 152788
rect 433426 152736 433432 152788
rect 433484 152776 433490 152788
rect 438946 152776 438952 152788
rect 433484 152748 438952 152776
rect 433484 152736 433490 152748
rect 438946 152736 438952 152748
rect 439004 152736 439010 152788
rect 442810 152736 442816 152788
rect 442868 152776 442874 152788
rect 456978 152776 456984 152788
rect 442868 152748 456984 152776
rect 442868 152736 442874 152748
rect 456978 152736 456984 152748
rect 457036 152736 457042 152788
rect 141844 152680 143764 152708
rect 141844 152668 141850 152680
rect 143810 152668 143816 152720
rect 143868 152708 143874 152720
rect 221274 152708 221280 152720
rect 143868 152680 221280 152708
rect 143868 152668 143874 152680
rect 221274 152668 221280 152680
rect 221332 152668 221338 152720
rect 224770 152668 224776 152720
rect 224828 152708 224834 152720
rect 288066 152708 288072 152720
rect 224828 152680 288072 152708
rect 224828 152668 224834 152680
rect 288066 152668 288072 152680
rect 288124 152668 288130 152720
rect 288342 152668 288348 152720
rect 288400 152708 288406 152720
rect 289998 152708 290004 152720
rect 288400 152680 290004 152708
rect 288400 152668 288406 152680
rect 289998 152668 290004 152680
rect 290056 152668 290062 152720
rect 291378 152668 291384 152720
rect 291436 152708 291442 152720
rect 341334 152708 341340 152720
rect 291436 152680 341340 152708
rect 291436 152668 291442 152680
rect 341334 152668 341340 152680
rect 341392 152668 341398 152720
rect 342438 152668 342444 152720
rect 342496 152708 342502 152720
rect 344554 152708 344560 152720
rect 342496 152680 344560 152708
rect 342496 152668 342502 152680
rect 344554 152668 344560 152680
rect 344612 152668 344618 152720
rect 347130 152708 347136 152720
rect 345492 152680 347136 152708
rect 15470 152600 15476 152652
rect 15528 152640 15534 152652
rect 130746 152640 130752 152652
rect 15528 152612 130752 152640
rect 15528 152600 15534 152612
rect 130746 152600 130752 152612
rect 130804 152600 130810 152652
rect 130838 152600 130844 152652
rect 130896 152640 130902 152652
rect 216122 152640 216128 152652
rect 130896 152612 216128 152640
rect 130896 152600 130902 152612
rect 216122 152600 216128 152612
rect 216180 152600 216186 152652
rect 220446 152600 220452 152652
rect 220504 152640 220510 152652
rect 284846 152640 284852 152652
rect 220504 152612 284852 152640
rect 220504 152600 220510 152612
rect 284846 152600 284852 152612
rect 284904 152600 284910 152652
rect 293218 152640 293224 152652
rect 287026 152612 293224 152640
rect 19702 152532 19708 152584
rect 19760 152572 19766 152584
rect 133966 152572 133972 152584
rect 19760 152544 133972 152572
rect 19760 152532 19766 152544
rect 133966 152532 133972 152544
rect 134024 152532 134030 152584
rect 135162 152532 135168 152584
rect 135220 152572 135226 152584
rect 138566 152572 138572 152584
rect 135220 152544 138572 152572
rect 135220 152532 135226 152544
rect 138566 152532 138572 152544
rect 138624 152532 138630 152584
rect 140774 152532 140780 152584
rect 140832 152572 140838 152584
rect 226426 152572 226432 152584
rect 140832 152544 226432 152572
rect 140832 152532 140838 152544
rect 226426 152532 226432 152544
rect 226484 152532 226490 152584
rect 228266 152532 228272 152584
rect 228324 152572 228330 152584
rect 287026 152572 287054 152612
rect 293218 152600 293224 152612
rect 293276 152600 293282 152652
rect 336182 152640 336188 152652
rect 296686 152612 336188 152640
rect 296686 152572 296714 152612
rect 336182 152600 336188 152612
rect 336240 152600 336246 152652
rect 336274 152600 336280 152652
rect 336332 152640 336338 152652
rect 345382 152640 345388 152652
rect 336332 152612 345388 152640
rect 336332 152600 336338 152612
rect 345382 152600 345388 152612
rect 345440 152600 345446 152652
rect 228324 152544 287054 152572
rect 290200 152544 296714 152572
rect 228324 152532 228330 152544
rect 2866 152464 2872 152516
rect 2924 152504 2930 152516
rect 121086 152504 121092 152516
rect 2924 152476 121092 152504
rect 2924 152464 2930 152476
rect 121086 152464 121092 152476
rect 121144 152464 121150 152516
rect 121178 152464 121184 152516
rect 121236 152504 121242 152516
rect 211062 152504 211068 152516
rect 121236 152476 211068 152504
rect 121236 152464 121242 152476
rect 211062 152464 211068 152476
rect 211120 152464 211126 152516
rect 211982 152464 211988 152516
rect 212040 152504 212046 152516
rect 277762 152504 277768 152516
rect 212040 152476 277768 152504
rect 212040 152464 212046 152476
rect 277762 152464 277768 152476
rect 277820 152464 277826 152516
rect 285858 152464 285864 152516
rect 285916 152504 285922 152516
rect 290200 152504 290228 152544
rect 299382 152532 299388 152584
rect 299440 152572 299446 152584
rect 345492 152572 345520 152680
rect 347130 152668 347136 152680
rect 347188 152668 347194 152720
rect 349062 152668 349068 152720
rect 349120 152708 349126 152720
rect 352374 152708 352380 152720
rect 349120 152680 352380 152708
rect 349120 152668 349126 152680
rect 352374 152668 352380 152680
rect 352432 152668 352438 152720
rect 352466 152668 352472 152720
rect 352524 152708 352530 152720
rect 382458 152708 382464 152720
rect 352524 152680 382464 152708
rect 352524 152668 352530 152680
rect 382458 152668 382464 152680
rect 382516 152668 382522 152720
rect 382550 152668 382556 152720
rect 382608 152708 382614 152720
rect 386966 152708 386972 152720
rect 382608 152680 386972 152708
rect 382608 152668 382614 152680
rect 386966 152668 386972 152680
rect 387024 152668 387030 152720
rect 387702 152668 387708 152720
rect 387760 152708 387766 152720
rect 413922 152708 413928 152720
rect 387760 152680 413928 152708
rect 387760 152668 387766 152680
rect 413922 152668 413928 152680
rect 413980 152668 413986 152720
rect 414014 152668 414020 152720
rect 414072 152708 414078 152720
rect 427078 152708 427084 152720
rect 414072 152680 427084 152708
rect 414072 152668 414078 152680
rect 427078 152668 427084 152680
rect 427136 152668 427142 152720
rect 427170 152668 427176 152720
rect 427228 152708 427234 152720
rect 431586 152708 431592 152720
rect 427228 152680 431592 152708
rect 427228 152668 427234 152680
rect 431586 152668 431592 152680
rect 431644 152668 431650 152720
rect 434622 152668 434628 152720
rect 434680 152708 434686 152720
rect 450538 152708 450544 152720
rect 434680 152680 450544 152708
rect 434680 152668 434686 152680
rect 450538 152668 450544 152680
rect 450596 152668 450602 152720
rect 458174 152668 458180 152720
rect 458232 152708 458238 152720
rect 463970 152708 463976 152720
rect 458232 152680 463976 152708
rect 458232 152668 458238 152680
rect 463970 152668 463976 152680
rect 464028 152668 464034 152720
rect 345566 152600 345572 152652
rect 345624 152640 345630 152652
rect 375374 152640 375380 152652
rect 345624 152612 375380 152640
rect 345624 152600 345630 152612
rect 375374 152600 375380 152612
rect 375432 152600 375438 152652
rect 375466 152600 375472 152652
rect 375524 152640 375530 152652
rect 405550 152640 405556 152652
rect 375524 152612 405556 152640
rect 375524 152600 375530 152612
rect 405550 152600 405556 152612
rect 405608 152600 405614 152652
rect 405642 152600 405648 152652
rect 405700 152640 405706 152652
rect 427998 152640 428004 152652
rect 405700 152612 428004 152640
rect 405700 152600 405706 152612
rect 427998 152600 428004 152612
rect 428056 152600 428062 152652
rect 428458 152600 428464 152652
rect 428516 152640 428522 152652
rect 446030 152640 446036 152652
rect 428516 152612 446036 152640
rect 428516 152600 428522 152612
rect 446030 152600 446036 152612
rect 446088 152600 446094 152652
rect 446950 152600 446956 152652
rect 447008 152640 447014 152652
rect 447008 152612 455828 152640
rect 447008 152600 447014 152612
rect 299440 152544 345520 152572
rect 299440 152532 299446 152544
rect 345658 152532 345664 152584
rect 345716 152572 345722 152584
rect 352282 152572 352288 152584
rect 345716 152544 352288 152572
rect 345716 152532 345722 152544
rect 352282 152532 352288 152544
rect 352340 152532 352346 152584
rect 352374 152532 352380 152584
rect 352432 152572 352438 152584
rect 385034 152572 385040 152584
rect 352432 152544 385040 152572
rect 352432 152532 352438 152544
rect 385034 152532 385040 152544
rect 385092 152532 385098 152584
rect 385494 152532 385500 152584
rect 385552 152572 385558 152584
rect 387610 152572 387616 152584
rect 385552 152544 387616 152572
rect 385552 152532 385558 152544
rect 387610 152532 387616 152544
rect 387668 152532 387674 152584
rect 393130 152532 393136 152584
rect 393188 152572 393194 152584
rect 419074 152572 419080 152584
rect 393188 152544 419080 152572
rect 393188 152532 393194 152544
rect 419074 152532 419080 152544
rect 419132 152532 419138 152584
rect 419258 152532 419264 152584
rect 419316 152572 419322 152584
rect 433426 152572 433432 152584
rect 419316 152544 433432 152572
rect 419316 152532 419322 152544
rect 433426 152532 433432 152544
rect 433484 152532 433490 152584
rect 433518 152532 433524 152584
rect 433576 152572 433582 152584
rect 433576 152544 438440 152572
rect 433576 152532 433582 152544
rect 285916 152476 290228 152504
rect 285916 152464 285922 152476
rect 291838 152464 291844 152516
rect 291896 152504 291902 152516
rect 336826 152504 336832 152516
rect 291896 152476 336832 152504
rect 291896 152464 291902 152476
rect 336826 152464 336832 152476
rect 336884 152464 336890 152516
rect 339494 152464 339500 152516
rect 339552 152504 339558 152516
rect 377306 152504 377312 152516
rect 339552 152476 377312 152504
rect 339552 152464 339558 152476
rect 377306 152464 377312 152476
rect 377364 152464 377370 152516
rect 378226 152464 378232 152516
rect 378284 152504 378290 152516
rect 379882 152504 379888 152516
rect 378284 152476 379888 152504
rect 378284 152464 378290 152476
rect 379882 152464 379888 152476
rect 379940 152464 379946 152516
rect 382182 152464 382188 152516
rect 382240 152504 382246 152516
rect 410702 152504 410708 152516
rect 382240 152476 410708 152504
rect 382240 152464 382246 152476
rect 410702 152464 410708 152476
rect 410760 152464 410766 152516
rect 431218 152504 431224 152516
rect 416516 152476 431224 152504
rect 56226 152396 56232 152448
rect 56284 152436 56290 152448
rect 141050 152436 141056 152448
rect 56284 152408 141056 152436
rect 56284 152396 56290 152408
rect 141050 152396 141056 152408
rect 141108 152396 141114 152448
rect 144086 152396 144092 152448
rect 144144 152436 144150 152448
rect 144144 152408 144408 152436
rect 144144 152396 144150 152408
rect 59998 152328 60004 152380
rect 60056 152368 60062 152380
rect 144270 152368 144276 152380
rect 60056 152340 144276 152368
rect 60056 152328 60062 152340
rect 144270 152328 144276 152340
rect 144328 152328 144334 152380
rect 144380 152368 144408 152408
rect 149054 152396 149060 152448
rect 149112 152436 149118 152448
rect 231578 152436 231584 152448
rect 149112 152408 231584 152436
rect 149112 152396 149118 152408
rect 231578 152396 231584 152408
rect 231636 152396 231642 152448
rect 245102 152396 245108 152448
rect 245160 152436 245166 152448
rect 306006 152436 306012 152448
rect 245160 152408 306012 152436
rect 245160 152396 245166 152408
rect 306006 152396 306012 152408
rect 306064 152396 306070 152448
rect 307294 152396 307300 152448
rect 307352 152436 307358 152448
rect 345658 152436 345664 152448
rect 307352 152408 345664 152436
rect 307352 152396 307358 152408
rect 345658 152396 345664 152408
rect 345716 152396 345722 152448
rect 345750 152396 345756 152448
rect 345808 152436 345814 152448
rect 346670 152436 346676 152448
rect 345808 152408 346676 152436
rect 345808 152396 345814 152408
rect 346670 152396 346676 152408
rect 346728 152396 346734 152448
rect 356146 152436 356152 152448
rect 350506 152408 356152 152436
rect 162210 152368 162216 152380
rect 144380 152340 162216 152368
rect 162210 152328 162216 152340
rect 162268 152328 162274 152380
rect 164418 152328 164424 152380
rect 164476 152368 164482 152380
rect 244366 152368 244372 152380
rect 164476 152340 244372 152368
rect 164476 152328 164482 152340
rect 244366 152328 244372 152340
rect 244424 152328 244430 152380
rect 255406 152328 255412 152380
rect 255464 152368 255470 152380
rect 313090 152368 313096 152380
rect 255464 152340 313096 152368
rect 255464 152328 255470 152340
rect 313090 152328 313096 152340
rect 313148 152328 313154 152380
rect 313182 152328 313188 152380
rect 313240 152368 313246 152380
rect 350506 152368 350534 152408
rect 356146 152396 356152 152408
rect 356204 152396 356210 152448
rect 389542 152436 389548 152448
rect 364306 152408 389548 152436
rect 313240 152340 350534 152368
rect 313240 152328 313246 152340
rect 354490 152328 354496 152380
rect 354548 152368 354554 152380
rect 364306 152368 364334 152408
rect 389542 152396 389548 152408
rect 389600 152396 389606 152448
rect 389634 152396 389640 152448
rect 389692 152436 389698 152448
rect 412634 152436 412640 152448
rect 389692 152408 412640 152436
rect 389692 152396 389698 152408
rect 412634 152396 412640 152408
rect 412692 152396 412698 152448
rect 354548 152340 364334 152368
rect 354548 152328 354554 152340
rect 364518 152328 364524 152380
rect 364576 152368 364582 152380
rect 369026 152368 369032 152380
rect 364576 152340 369032 152368
rect 364576 152328 364582 152340
rect 369026 152328 369032 152340
rect 369084 152328 369090 152380
rect 371326 152328 371332 152380
rect 371384 152368 371390 152380
rect 402330 152368 402336 152380
rect 371384 152340 402336 152368
rect 371384 152328 371390 152340
rect 402330 152328 402336 152340
rect 402388 152328 402394 152380
rect 405826 152328 405832 152380
rect 405884 152368 405890 152380
rect 408770 152368 408776 152380
rect 405884 152340 408776 152368
rect 405884 152328 405890 152340
rect 408770 152328 408776 152340
rect 408828 152328 408834 152380
rect 409138 152328 409144 152380
rect 409196 152368 409202 152380
rect 409196 152340 410196 152368
rect 409196 152328 409202 152340
rect 76742 152260 76748 152312
rect 76800 152300 76806 152312
rect 159634 152300 159640 152312
rect 76800 152272 159640 152300
rect 76800 152260 76806 152272
rect 159634 152260 159640 152272
rect 159692 152260 159698 152312
rect 172606 152260 172612 152312
rect 172664 152300 172670 152312
rect 249518 152300 249524 152312
rect 172664 152272 249524 152300
rect 172664 152260 172670 152272
rect 249518 152260 249524 152272
rect 249576 152260 249582 152312
rect 265342 152260 265348 152312
rect 265400 152300 265406 152312
rect 270862 152300 270868 152312
rect 265400 152272 270868 152300
rect 265400 152260 265406 152272
rect 270862 152260 270868 152272
rect 270920 152260 270926 152312
rect 272518 152260 272524 152312
rect 272576 152300 272582 152312
rect 316310 152300 316316 152312
rect 272576 152272 316316 152300
rect 272576 152260 272582 152272
rect 316310 152260 316316 152272
rect 316368 152260 316374 152312
rect 320266 152260 320272 152312
rect 320324 152300 320330 152312
rect 323394 152300 323400 152312
rect 320324 152272 323400 152300
rect 320324 152260 320330 152272
rect 323394 152260 323400 152272
rect 323452 152260 323458 152312
rect 323486 152260 323492 152312
rect 323544 152300 323550 152312
rect 330386 152300 330392 152312
rect 323544 152272 330392 152300
rect 323544 152260 323550 152272
rect 330386 152260 330392 152272
rect 330444 152260 330450 152312
rect 330938 152260 330944 152312
rect 330996 152300 331002 152312
rect 371510 152300 371516 152312
rect 330996 152272 371516 152300
rect 330996 152260 331002 152272
rect 371510 152260 371516 152272
rect 371568 152260 371574 152312
rect 381354 152260 381360 152312
rect 381412 152300 381418 152312
rect 410058 152300 410064 152312
rect 381412 152272 410064 152300
rect 381412 152260 381418 152272
rect 410058 152260 410064 152272
rect 410116 152260 410122 152312
rect 410168 152300 410196 152340
rect 410886 152328 410892 152380
rect 410944 152368 410950 152380
rect 416516 152368 416544 152476
rect 431218 152464 431224 152476
rect 431276 152464 431282 152516
rect 431310 152464 431316 152516
rect 431368 152504 431374 152516
rect 436738 152504 436744 152516
rect 431368 152476 436744 152504
rect 431368 152464 431374 152476
rect 436738 152464 436744 152476
rect 436796 152464 436802 152516
rect 438302 152504 438308 152516
rect 436848 152476 438308 152504
rect 418430 152396 418436 152448
rect 418488 152436 418494 152448
rect 436848 152436 436876 152476
rect 438302 152464 438308 152476
rect 438360 152464 438366 152516
rect 438412 152504 438440 152544
rect 438486 152532 438492 152584
rect 438544 152572 438550 152584
rect 440970 152572 440976 152584
rect 438544 152544 440976 152572
rect 438544 152532 438550 152544
rect 440970 152532 440976 152544
rect 441028 152532 441034 152584
rect 441430 152532 441436 152584
rect 441488 152572 441494 152584
rect 455690 152572 455696 152584
rect 441488 152544 455696 152572
rect 441488 152532 441494 152544
rect 455690 152532 455696 152544
rect 455748 152532 455754 152584
rect 455800 152572 455828 152612
rect 459646 152600 459652 152652
rect 459704 152640 459710 152652
rect 465258 152640 465264 152652
rect 459704 152612 465264 152640
rect 459704 152600 459710 152612
rect 465258 152600 465264 152612
rect 465316 152600 465322 152652
rect 460106 152572 460112 152584
rect 455800 152544 460112 152572
rect 460106 152532 460112 152544
rect 460164 152532 460170 152584
rect 449894 152504 449900 152516
rect 438412 152476 449900 152504
rect 449894 152464 449900 152476
rect 449952 152464 449958 152516
rect 418488 152408 436876 152436
rect 418488 152396 418494 152408
rect 437750 152396 437756 152448
rect 437808 152436 437814 152448
rect 453114 152436 453120 152448
rect 437808 152408 453120 152436
rect 437808 152396 437814 152408
rect 453114 152396 453120 152408
rect 453172 152396 453178 152448
rect 428642 152368 428648 152380
rect 410944 152340 416544 152368
rect 422266 152340 428648 152368
rect 410944 152328 410950 152340
rect 422266 152300 422294 152340
rect 428642 152328 428648 152340
rect 428700 152328 428706 152380
rect 431034 152328 431040 152380
rect 431092 152368 431098 152380
rect 447962 152368 447968 152380
rect 431092 152340 447968 152368
rect 431092 152328 431098 152340
rect 447962 152328 447968 152340
rect 448020 152328 448026 152380
rect 410168 152272 422294 152300
rect 423582 152260 423588 152312
rect 423640 152300 423646 152312
rect 426250 152300 426256 152312
rect 423640 152272 426256 152300
rect 423640 152260 423646 152272
rect 426250 152260 426256 152272
rect 426308 152260 426314 152312
rect 426342 152260 426348 152312
rect 426400 152300 426406 152312
rect 431310 152300 431316 152312
rect 426400 152272 431316 152300
rect 426400 152260 426406 152272
rect 431310 152260 431316 152272
rect 431368 152260 431374 152312
rect 442166 152300 442172 152312
rect 431420 152272 442172 152300
rect 85482 152192 85488 152244
rect 85540 152232 85546 152244
rect 164786 152232 164792 152244
rect 85540 152204 164792 152232
rect 85540 152192 85546 152204
rect 164786 152192 164792 152204
rect 164844 152192 164850 152244
rect 166994 152192 167000 152244
rect 167052 152232 167058 152244
rect 182726 152232 182732 152244
rect 167052 152204 182732 152232
rect 167052 152192 167058 152204
rect 182726 152192 182732 152204
rect 182784 152192 182790 152244
rect 183094 152192 183100 152244
rect 183152 152232 183158 152244
rect 195606 152232 195612 152244
rect 183152 152204 195612 152232
rect 183152 152192 183158 152204
rect 195606 152192 195612 152204
rect 195664 152192 195670 152244
rect 218698 152232 218704 152244
rect 195716 152204 218704 152232
rect 75086 152124 75092 152176
rect 75144 152164 75150 152176
rect 154482 152164 154488 152176
rect 75144 152136 154488 152164
rect 75144 152124 75150 152136
rect 154482 152124 154488 152136
rect 154540 152124 154546 152176
rect 156046 152124 156052 152176
rect 156104 152164 156110 152176
rect 172514 152164 172520 152176
rect 156104 152136 172520 152164
rect 156104 152124 156110 152136
rect 172514 152124 172520 152136
rect 172572 152124 172578 152176
rect 176654 152124 176660 152176
rect 176712 152164 176718 152176
rect 190454 152164 190460 152176
rect 176712 152136 190460 152164
rect 176712 152124 176718 152136
rect 190454 152124 190460 152136
rect 190512 152124 190518 152176
rect 195146 152124 195152 152176
rect 195204 152164 195210 152176
rect 195716 152164 195744 152204
rect 218698 152192 218704 152204
rect 218756 152192 218762 152244
rect 221458 152192 221464 152244
rect 221516 152232 221522 152244
rect 282914 152232 282920 152244
rect 221516 152204 282920 152232
rect 221516 152192 221522 152204
rect 282914 152192 282920 152204
rect 282972 152192 282978 152244
rect 285490 152192 285496 152244
rect 285548 152232 285554 152244
rect 291838 152232 291844 152244
rect 285548 152204 291844 152232
rect 285548 152192 285554 152204
rect 291838 152192 291844 152204
rect 291896 152192 291902 152244
rect 292482 152192 292488 152244
rect 292540 152232 292546 152244
rect 341978 152232 341984 152244
rect 292540 152204 341984 152232
rect 292540 152192 292546 152204
rect 341978 152192 341984 152204
rect 342036 152192 342042 152244
rect 342254 152192 342260 152244
rect 342312 152232 342318 152244
rect 346486 152232 346492 152244
rect 342312 152204 346492 152232
rect 342312 152192 342318 152204
rect 346486 152192 346492 152204
rect 346544 152192 346550 152244
rect 346578 152192 346584 152244
rect 346636 152232 346642 152244
rect 380526 152232 380532 152244
rect 346636 152204 380532 152232
rect 346636 152192 346642 152204
rect 380526 152192 380532 152204
rect 380584 152192 380590 152244
rect 384942 152192 384948 152244
rect 385000 152232 385006 152244
rect 392118 152232 392124 152244
rect 385000 152204 392124 152232
rect 385000 152192 385006 152204
rect 392118 152192 392124 152204
rect 392176 152192 392182 152244
rect 394326 152192 394332 152244
rect 394384 152232 394390 152244
rect 417786 152232 417792 152244
rect 394384 152204 417792 152232
rect 394384 152192 394390 152204
rect 417786 152192 417792 152204
rect 417844 152192 417850 152244
rect 417878 152192 417884 152244
rect 417936 152232 417942 152244
rect 421742 152232 421748 152244
rect 417936 152204 421748 152232
rect 417936 152192 417942 152204
rect 421742 152192 421748 152204
rect 421800 152192 421806 152244
rect 423398 152192 423404 152244
rect 423456 152232 423462 152244
rect 431420 152232 431448 152272
rect 442166 152260 442172 152272
rect 442224 152260 442230 152312
rect 456334 152300 456340 152312
rect 442276 152272 456340 152300
rect 423456 152204 431448 152232
rect 423456 152192 423462 152204
rect 431494 152192 431500 152244
rect 431552 152232 431558 152244
rect 441522 152232 441528 152244
rect 431552 152204 441528 152232
rect 431552 152192 431558 152204
rect 441522 152192 441528 152204
rect 441580 152192 441586 152244
rect 441982 152192 441988 152244
rect 442040 152232 442046 152244
rect 442276 152232 442304 152272
rect 456334 152260 456340 152272
rect 456392 152260 456398 152312
rect 442040 152204 442304 152232
rect 442040 152192 442046 152204
rect 443638 152192 443644 152244
rect 443696 152232 443702 152244
rect 457622 152232 457628 152244
rect 443696 152204 457628 152232
rect 443696 152192 443702 152204
rect 457622 152192 457628 152204
rect 457680 152192 457686 152244
rect 213546 152164 213552 152176
rect 195204 152136 195744 152164
rect 195808 152136 213552 152164
rect 195204 152124 195210 152136
rect 71774 152056 71780 152108
rect 71832 152096 71838 152108
rect 149422 152096 149428 152108
rect 71832 152068 149428 152096
rect 71832 152056 71838 152068
rect 149422 152056 149428 152068
rect 149480 152056 149486 152108
rect 150434 152056 150440 152108
rect 150492 152096 150498 152108
rect 167362 152096 167368 152108
rect 150492 152068 167368 152096
rect 150492 152056 150498 152068
rect 167362 152056 167368 152068
rect 167420 152056 167426 152108
rect 169754 152056 169760 152108
rect 169812 152096 169818 152108
rect 185302 152096 185308 152108
rect 169812 152068 185308 152096
rect 169812 152056 169818 152068
rect 185302 152056 185308 152068
rect 185360 152056 185366 152108
rect 193122 152056 193128 152108
rect 193180 152096 193186 152108
rect 195808 152096 195836 152136
rect 213546 152124 213552 152136
rect 213604 152124 213610 152176
rect 213730 152124 213736 152176
rect 213788 152164 213794 152176
rect 274542 152164 274548 152176
rect 213788 152136 274548 152164
rect 213788 152124 213794 152136
rect 274542 152124 274548 152136
rect 274600 152124 274606 152176
rect 277946 152124 277952 152176
rect 278004 152164 278010 152176
rect 331122 152164 331128 152176
rect 278004 152136 331128 152164
rect 278004 152124 278010 152136
rect 331122 152124 331128 152136
rect 331180 152124 331186 152176
rect 331858 152124 331864 152176
rect 331916 152164 331922 152176
rect 372154 152164 372160 152176
rect 331916 152136 372160 152164
rect 331916 152124 331922 152136
rect 372154 152124 372160 152136
rect 372212 152124 372218 152176
rect 388346 152124 388352 152176
rect 388404 152164 388410 152176
rect 407482 152164 407488 152176
rect 388404 152136 407488 152164
rect 388404 152124 388410 152136
rect 407482 152124 407488 152136
rect 407540 152124 407546 152176
rect 415118 152124 415124 152176
rect 415176 152164 415182 152176
rect 423582 152164 423588 152176
rect 415176 152136 423588 152164
rect 415176 152124 415182 152136
rect 423582 152124 423588 152136
rect 423640 152124 423646 152176
rect 427078 152124 427084 152176
rect 427136 152164 427142 152176
rect 433794 152164 433800 152176
rect 427136 152136 433800 152164
rect 427136 152124 427142 152136
rect 433794 152124 433800 152136
rect 433852 152124 433858 152176
rect 436738 152124 436744 152176
rect 436796 152164 436802 152176
rect 444098 152164 444104 152176
rect 436796 152136 444104 152164
rect 436796 152124 436802 152136
rect 444098 152124 444104 152136
rect 444156 152124 444162 152176
rect 445662 152124 445668 152176
rect 445720 152164 445726 152176
rect 458818 152164 458824 152176
rect 445720 152136 458824 152164
rect 445720 152124 445726 152136
rect 458818 152124 458824 152136
rect 458876 152124 458882 152176
rect 516686 152124 516692 152176
rect 516744 152164 516750 152176
rect 520274 152164 520280 152176
rect 516744 152136 520280 152164
rect 516744 152124 516750 152136
rect 520274 152124 520280 152136
rect 520332 152124 520338 152176
rect 193180 152068 195836 152096
rect 193180 152056 193186 152068
rect 195882 152056 195888 152108
rect 195940 152096 195946 152108
rect 208486 152096 208492 152108
rect 195940 152068 208492 152096
rect 195940 152056 195946 152068
rect 208486 152056 208492 152068
rect 208544 152056 208550 152108
rect 272702 152096 272708 152108
rect 215266 152068 272708 152096
rect 109678 151988 109684 152040
rect 109736 152028 109742 152040
rect 128170 152028 128176 152040
rect 109736 152000 128176 152028
rect 109736 151988 109742 152000
rect 128170 151988 128176 152000
rect 128228 151988 128234 152040
rect 128354 151988 128360 152040
rect 128412 152028 128418 152040
rect 203334 152028 203340 152040
rect 128412 152000 203340 152028
rect 128412 151988 128418 152000
rect 203334 151988 203340 152000
rect 203392 151988 203398 152040
rect 212626 151988 212632 152040
rect 212684 152028 212690 152040
rect 215266 152028 215294 152068
rect 272702 152056 272708 152068
rect 272760 152056 272766 152108
rect 272794 152056 272800 152108
rect 272852 152096 272858 152108
rect 325970 152096 325976 152108
rect 272852 152068 325976 152096
rect 272852 152056 272858 152068
rect 325970 152056 325976 152068
rect 326028 152056 326034 152108
rect 330386 152056 330392 152108
rect 330444 152096 330450 152108
rect 362586 152096 362592 152108
rect 330444 152068 362592 152096
rect 330444 152056 330450 152068
rect 362586 152056 362592 152068
rect 362644 152056 362650 152108
rect 388438 152056 388444 152108
rect 388496 152096 388502 152108
rect 404906 152096 404912 152108
rect 388496 152068 404912 152096
rect 388496 152056 388502 152068
rect 404906 152056 404912 152068
rect 404964 152056 404970 152108
rect 405366 152056 405372 152108
rect 405424 152096 405430 152108
rect 421006 152096 421012 152108
rect 405424 152068 421012 152096
rect 405424 152056 405430 152068
rect 421006 152056 421012 152068
rect 421064 152056 421070 152108
rect 426802 152096 426808 152108
rect 422266 152068 426808 152096
rect 212684 152000 215294 152028
rect 212684 151988 212690 152000
rect 242434 151988 242440 152040
rect 242492 152028 242498 152040
rect 300946 152028 300952 152040
rect 242492 152000 300952 152028
rect 242492 151988 242498 152000
rect 300946 151988 300952 152000
rect 301004 151988 301010 152040
rect 304810 151988 304816 152040
rect 304868 152028 304874 152040
rect 351638 152028 351644 152040
rect 304868 152000 351644 152028
rect 304868 151988 304874 152000
rect 351638 151988 351644 152000
rect 351696 151988 351702 152040
rect 352742 151988 352748 152040
rect 352800 152028 352806 152040
rect 388254 152028 388260 152040
rect 352800 152000 388260 152028
rect 352800 151988 352806 152000
rect 388254 151988 388260 152000
rect 388312 151988 388318 152040
rect 403434 151988 403440 152040
rect 403492 152028 403498 152040
rect 418430 152028 418436 152040
rect 403492 152000 418436 152028
rect 403492 151988 403498 152000
rect 418430 151988 418436 152000
rect 418488 151988 418494 152040
rect 422266 152028 422294 152068
rect 426802 152056 426808 152068
rect 426860 152056 426866 152108
rect 426894 152056 426900 152108
rect 426952 152096 426958 152108
rect 444742 152096 444748 152108
rect 426952 152068 444748 152096
rect 426952 152056 426958 152068
rect 444742 152056 444748 152068
rect 444800 152056 444806 152108
rect 515490 152056 515496 152108
rect 515548 152096 515554 152108
rect 518986 152096 518992 152108
rect 515548 152068 518992 152096
rect 515548 152056 515554 152068
rect 518986 152056 518992 152068
rect 519044 152056 519050 152108
rect 418540 152000 422294 152028
rect 107562 151920 107568 151972
rect 107620 151960 107626 151972
rect 175090 151960 175096 151972
rect 107620 151932 175096 151960
rect 107620 151920 107626 151932
rect 175090 151920 175096 151932
rect 175148 151920 175154 151972
rect 185578 151920 185584 151972
rect 185636 151960 185642 151972
rect 200758 151960 200764 151972
rect 185636 151932 200764 151960
rect 185636 151920 185642 151932
rect 200758 151920 200764 151932
rect 200816 151920 200822 151972
rect 243354 151920 243360 151972
rect 243412 151960 243418 151972
rect 302878 151960 302884 151972
rect 243412 151932 302884 151960
rect 243412 151920 243418 151932
rect 302878 151920 302884 151932
rect 302936 151920 302942 151972
rect 326614 151960 326620 151972
rect 316006 151932 326620 151960
rect 30190 151852 30196 151904
rect 30248 151892 30254 151904
rect 74534 151892 74540 151904
rect 30248 151864 74540 151892
rect 30248 151852 30254 151864
rect 74534 151852 74540 151864
rect 74592 151852 74598 151904
rect 109126 151852 109132 151904
rect 109184 151892 109190 151904
rect 138474 151892 138480 151904
rect 109184 151864 138480 151892
rect 109184 151852 109190 151864
rect 138474 151852 138480 151864
rect 138532 151852 138538 151904
rect 138566 151852 138572 151904
rect 138624 151892 138630 151904
rect 146846 151892 146852 151904
rect 138624 151864 146852 151892
rect 138624 151852 138630 151864
rect 146846 151852 146852 151864
rect 146904 151852 146910 151904
rect 157058 151892 157064 151904
rect 151786 151864 157064 151892
rect 33594 151784 33600 151836
rect 33652 151824 33658 151836
rect 84194 151824 84200 151836
rect 33652 151796 84200 151824
rect 33652 151784 33658 151796
rect 84194 151784 84200 151796
rect 84252 151784 84258 151836
rect 105814 151784 105820 151836
rect 105872 151824 105878 151836
rect 110322 151824 110328 151836
rect 105872 151796 110328 151824
rect 105872 151784 105878 151796
rect 110322 151784 110328 151796
rect 110380 151784 110386 151836
rect 113910 151784 113916 151836
rect 113968 151824 113974 151836
rect 123478 151824 123484 151836
rect 113968 151796 123484 151824
rect 113968 151784 113974 151796
rect 123478 151784 123484 151796
rect 123536 151784 123542 151836
rect 138014 151784 138020 151836
rect 138072 151824 138078 151836
rect 141786 151824 141792 151836
rect 138072 151796 141792 151824
rect 138072 151784 138078 151796
rect 141786 151784 141792 151796
rect 141844 151784 141850 151836
rect 143258 151784 143264 151836
rect 143316 151824 143322 151836
rect 151786 151824 151814 151864
rect 157058 151852 157064 151864
rect 157116 151852 157122 151904
rect 160186 151852 160192 151904
rect 160244 151892 160250 151904
rect 177666 151892 177672 151904
rect 160244 151864 177672 151892
rect 160244 151852 160250 151864
rect 177666 151852 177672 151864
rect 177724 151852 177730 151904
rect 191650 151852 191656 151904
rect 191708 151892 191714 151904
rect 195882 151892 195888 151904
rect 191708 151864 195888 151892
rect 191708 151852 191714 151864
rect 195882 151852 195888 151864
rect 195940 151852 195946 151904
rect 272610 151852 272616 151904
rect 272668 151892 272674 151904
rect 316006 151892 316034 151932
rect 326614 151920 326620 151932
rect 326672 151920 326678 151972
rect 335326 151932 354674 151960
rect 272668 151864 316034 151892
rect 272668 151852 272674 151864
rect 325050 151852 325056 151904
rect 325108 151892 325114 151904
rect 335326 151892 335354 151932
rect 325108 151864 335354 151892
rect 325108 151852 325114 151864
rect 343818 151852 343824 151904
rect 343876 151892 343882 151904
rect 346578 151892 346584 151904
rect 343876 151864 346584 151892
rect 343876 151852 343882 151864
rect 346578 151852 346584 151864
rect 346636 151852 346642 151904
rect 346670 151852 346676 151904
rect 346728 151892 346734 151904
rect 352466 151892 352472 151904
rect 346728 151864 352472 151892
rect 346728 151852 346734 151864
rect 352466 151852 352472 151864
rect 352524 151852 352530 151904
rect 143316 151796 151814 151824
rect 143316 151784 143322 151796
rect 261018 151784 261024 151836
rect 261076 151824 261082 151836
rect 272518 151824 272524 151836
rect 261076 151796 272524 151824
rect 261076 151784 261082 151796
rect 272518 151784 272524 151796
rect 272576 151784 272582 151836
rect 283006 151784 283012 151836
rect 283064 151824 283070 151836
rect 287422 151824 287428 151836
rect 283064 151796 287428 151824
rect 283064 151784 283070 151796
rect 287422 151784 287428 151796
rect 287480 151784 287486 151836
rect 303982 151784 303988 151836
rect 304040 151824 304046 151836
rect 350994 151824 351000 151836
rect 304040 151796 351000 151824
rect 304040 151784 304046 151796
rect 350994 151784 351000 151796
rect 351052 151784 351058 151836
rect 354646 151824 354674 151932
rect 362954 151920 362960 151972
rect 363012 151960 363018 151972
rect 364518 151960 364524 151972
rect 363012 151932 364524 151960
rect 363012 151920 363018 151932
rect 364518 151920 364524 151932
rect 364576 151920 364582 151972
rect 386230 151920 386236 151972
rect 386288 151960 386294 151972
rect 399754 151960 399760 151972
rect 386288 151932 399760 151960
rect 386288 151920 386294 151932
rect 399754 151920 399760 151932
rect 399812 151920 399818 151972
rect 399846 151920 399852 151972
rect 399904 151960 399910 151972
rect 399904 151932 403848 151960
rect 399904 151920 399910 151932
rect 355318 151852 355324 151904
rect 355376 151892 355382 151904
rect 390186 151892 390192 151904
rect 355376 151864 390192 151892
rect 355376 151852 355382 151864
rect 390186 151852 390192 151864
rect 390244 151852 390250 151904
rect 367002 151824 367008 151836
rect 354646 151796 367008 151824
rect 367002 151784 367008 151796
rect 367060 151784 367066 151836
rect 378778 151784 378784 151836
rect 378836 151824 378842 151836
rect 384390 151824 384396 151836
rect 378836 151796 384396 151824
rect 378836 151784 378842 151796
rect 384390 151784 384396 151796
rect 384448 151784 384454 151836
rect 385310 151784 385316 151836
rect 385368 151824 385374 151836
rect 394694 151824 394700 151836
rect 385368 151796 394700 151824
rect 385368 151784 385374 151796
rect 394694 151784 394700 151796
rect 394752 151784 394758 151836
rect 396166 151784 396172 151836
rect 396224 151824 396230 151836
rect 402974 151824 402980 151836
rect 396224 151796 402980 151824
rect 396224 151784 396230 151796
rect 402974 151784 402980 151796
rect 403032 151784 403038 151836
rect 403820 151824 403848 151932
rect 413830 151920 413836 151972
rect 413888 151960 413894 151972
rect 416498 151960 416504 151972
rect 413888 151932 416504 151960
rect 413888 151920 413894 151932
rect 416498 151920 416504 151932
rect 416556 151920 416562 151972
rect 416590 151920 416596 151972
rect 416648 151960 416654 151972
rect 418540 151960 418568 152000
rect 422570 151988 422576 152040
rect 422628 152028 422634 152040
rect 431494 152028 431500 152040
rect 422628 152000 431500 152028
rect 422628 151988 422634 152000
rect 431494 151988 431500 152000
rect 431552 151988 431558 152040
rect 431586 151988 431592 152040
rect 431644 152028 431650 152040
rect 439590 152028 439596 152040
rect 431644 152000 439596 152028
rect 431644 151988 431650 152000
rect 439590 151988 439596 152000
rect 439648 151988 439654 152040
rect 454402 152028 454408 152040
rect 439700 152000 454408 152028
rect 416648 151932 418568 151960
rect 416648 151920 416654 151932
rect 419534 151920 419540 151972
rect 419592 151960 419598 151972
rect 437014 151960 437020 151972
rect 419592 151932 437020 151960
rect 419592 151920 419598 151932
rect 437014 151920 437020 151932
rect 437072 151920 437078 151972
rect 439406 151920 439412 151972
rect 439464 151960 439470 151972
rect 439700 151960 439728 152000
rect 454402 151988 454408 152000
rect 454460 151988 454466 152040
rect 456794 151988 456800 152040
rect 456852 152028 456858 152040
rect 463326 152028 463332 152040
rect 456852 152000 463332 152028
rect 456852 151988 456858 152000
rect 463326 151988 463332 152000
rect 463384 151988 463390 152040
rect 486510 151988 486516 152040
rect 486568 152028 486574 152040
rect 490282 152028 490288 152040
rect 486568 152000 490288 152028
rect 486568 151988 486574 152000
rect 490282 151988 490288 152000
rect 490340 151988 490346 152040
rect 515950 151988 515956 152040
rect 516008 152028 516014 152040
rect 519906 152028 519912 152040
rect 516008 152000 519912 152028
rect 516008 151988 516014 152000
rect 519906 151988 519912 152000
rect 519964 151988 519970 152040
rect 451826 151960 451832 151972
rect 439464 151932 439728 151960
rect 439792 151932 451832 151960
rect 439464 151920 439470 151932
rect 403894 151852 403900 151904
rect 403952 151892 403958 151904
rect 415854 151892 415860 151904
rect 403952 151864 415860 151892
rect 403952 151852 403958 151864
rect 415854 151852 415860 151864
rect 415912 151852 415918 151904
rect 421650 151892 421656 151904
rect 415964 151864 421656 151892
rect 413278 151824 413284 151836
rect 403820 151796 413284 151824
rect 413278 151784 413284 151796
rect 413336 151784 413342 151836
rect 413646 151784 413652 151836
rect 413704 151824 413710 151836
rect 415964 151824 415992 151864
rect 421650 151852 421656 151864
rect 421708 151852 421714 151904
rect 421742 151852 421748 151904
rect 421800 151892 421806 151904
rect 431862 151892 431868 151904
rect 421800 151864 431868 151892
rect 421800 151852 421806 151864
rect 431862 151852 431868 151864
rect 431920 151852 431926 151904
rect 433334 151852 433340 151904
rect 433392 151892 433398 151904
rect 433392 151864 434576 151892
rect 433392 151852 433398 151864
rect 413704 151796 415992 151824
rect 413704 151784 413710 151796
rect 419626 151784 419632 151836
rect 419684 151824 419690 151836
rect 434438 151824 434444 151836
rect 419684 151796 434444 151824
rect 419684 151784 419690 151796
rect 434438 151784 434444 151796
rect 434496 151784 434502 151836
rect 434548 151824 434576 151864
rect 436094 151852 436100 151904
rect 436152 151892 436158 151904
rect 439792 151892 439820 151932
rect 451826 151920 451832 151932
rect 451884 151920 451890 151972
rect 456058 151920 456064 151972
rect 456116 151960 456122 151972
rect 461394 151960 461400 151972
rect 456116 151932 461400 151960
rect 456116 151920 456122 151932
rect 461394 151920 461400 151932
rect 461452 151920 461458 151972
rect 469214 151920 469220 151972
rect 469272 151960 469278 151972
rect 472342 151960 472348 151972
rect 469272 151932 472348 151960
rect 469272 151920 469278 151932
rect 472342 151920 472348 151932
rect 472400 151920 472406 151972
rect 487338 151920 487344 151972
rect 487396 151960 487402 151972
rect 490926 151960 490932 151972
rect 487396 151932 490932 151960
rect 487396 151920 487402 151932
rect 490926 151920 490932 151932
rect 490984 151920 490990 151972
rect 507670 151920 507676 151972
rect 507728 151960 507734 151972
rect 509234 151960 509240 151972
rect 507728 151932 509240 151960
rect 507728 151920 507734 151932
rect 509234 151920 509240 151932
rect 509292 151920 509298 151972
rect 517422 151920 517428 151972
rect 517480 151960 517486 151972
rect 521562 151960 521568 151972
rect 517480 151932 521568 151960
rect 517480 151920 517486 151932
rect 521562 151920 521568 151932
rect 521620 151920 521626 151972
rect 440878 151892 440884 151904
rect 436152 151864 439820 151892
rect 439884 151864 440884 151892
rect 436152 151852 436158 151864
rect 439884 151824 439912 151864
rect 440878 151852 440884 151864
rect 440936 151852 440942 151904
rect 440970 151852 440976 151904
rect 441028 151892 441034 151904
rect 451182 151892 451188 151904
rect 441028 151864 451188 151892
rect 441028 151852 441034 151864
rect 451182 151852 451188 151864
rect 451240 151852 451246 151904
rect 457162 151852 457168 151904
rect 457220 151892 457226 151904
rect 462682 151892 462688 151904
rect 457220 151864 462688 151892
rect 457220 151852 457226 151864
rect 462682 151852 462688 151864
rect 462740 151852 462746 151904
rect 468018 151852 468024 151904
rect 468076 151892 468082 151904
rect 471054 151892 471060 151904
rect 468076 151864 471060 151892
rect 468076 151852 468082 151864
rect 471054 151852 471060 151864
rect 471112 151852 471118 151904
rect 489086 151852 489092 151904
rect 489144 151892 489150 151904
rect 492214 151892 492220 151904
rect 489144 151864 492220 151892
rect 489144 151852 489150 151864
rect 492214 151852 492220 151864
rect 492272 151852 492278 151904
rect 499482 151852 499488 151904
rect 499540 151892 499546 151904
rect 499942 151892 499948 151904
rect 499540 151864 499948 151892
rect 499540 151852 499546 151864
rect 499942 151852 499948 151864
rect 500000 151852 500006 151904
rect 434548 151796 439912 151824
rect 440234 151784 440240 151836
rect 440292 151824 440298 151836
rect 455046 151824 455052 151836
rect 440292 151796 455052 151824
rect 440292 151784 440298 151796
rect 455046 151784 455052 151796
rect 455104 151784 455110 151836
rect 455782 151784 455788 151836
rect 455840 151824 455846 151836
rect 462038 151824 462044 151836
rect 455840 151796 462044 151824
rect 455840 151784 455846 151796
rect 462038 151784 462044 151796
rect 462096 151784 462102 151836
rect 467926 151784 467932 151836
rect 467984 151824 467990 151836
rect 471698 151824 471704 151836
rect 467984 151796 471704 151824
rect 467984 151784 467990 151796
rect 471698 151784 471704 151796
rect 471756 151784 471762 151836
rect 488442 151784 488448 151836
rect 488500 151824 488506 151836
rect 491570 151824 491576 151836
rect 488500 151796 491576 151824
rect 488500 151784 488506 151796
rect 491570 151784 491576 151796
rect 491628 151784 491634 151836
rect 509050 151784 509056 151836
rect 509108 151824 509114 151836
rect 510890 151824 510896 151836
rect 509108 151796 510896 151824
rect 509108 151784 509114 151796
rect 510890 151784 510896 151796
rect 510948 151784 510954 151836
rect 84194 151376 84200 151428
rect 84252 151416 84258 151428
rect 117222 151416 117228 151428
rect 84252 151388 117228 151416
rect 84252 151376 84258 151388
rect 117222 151376 117228 151388
rect 117280 151376 117286 151428
rect 74534 151308 74540 151360
rect 74592 151348 74598 151360
rect 117130 151348 117136 151360
rect 74592 151320 117136 151348
rect 74592 151308 74598 151320
rect 117130 151308 117136 151320
rect 117188 151308 117194 151360
rect 68002 151240 68008 151292
rect 68060 151280 68066 151292
rect 112806 151280 112812 151292
rect 68060 151252 112812 151280
rect 68060 151240 68066 151252
rect 112806 151240 112812 151252
rect 112864 151240 112870 151292
rect 64506 151172 64512 151224
rect 64564 151212 64570 151224
rect 112714 151212 112720 151224
rect 64564 151184 112720 151212
rect 64564 151172 64570 151184
rect 112714 151172 112720 151184
rect 112772 151172 112778 151224
rect 61102 151104 61108 151156
rect 61160 151144 61166 151156
rect 112622 151144 112628 151156
rect 61160 151116 112628 151144
rect 61160 151104 61166 151116
rect 112622 151104 112628 151116
rect 112680 151104 112686 151156
rect 57698 151036 57704 151088
rect 57756 151076 57762 151088
rect 112530 151076 112536 151088
rect 57756 151048 112536 151076
rect 57756 151036 57762 151048
rect 112530 151036 112536 151048
rect 112588 151036 112594 151088
rect 54202 150968 54208 151020
rect 54260 151008 54266 151020
rect 111610 151008 111616 151020
rect 54260 150980 111616 151008
rect 54260 150968 54266 150980
rect 111610 150968 111616 150980
rect 111668 150968 111674 151020
rect 50798 150900 50804 150952
rect 50856 150940 50862 150952
rect 112438 150940 112444 150952
rect 50856 150912 112444 150940
rect 50856 150900 50862 150912
rect 112438 150900 112444 150912
rect 112496 150900 112502 150952
rect 47302 150832 47308 150884
rect 47360 150872 47366 150884
rect 111518 150872 111524 150884
rect 47360 150844 111524 150872
rect 47360 150832 47366 150844
rect 111518 150832 111524 150844
rect 111576 150832 111582 150884
rect 43898 150764 43904 150816
rect 43956 150804 43962 150816
rect 111426 150804 111432 150816
rect 43956 150776 111432 150804
rect 43956 150764 43962 150776
rect 111426 150764 111432 150776
rect 111484 150764 111490 150816
rect 40494 150696 40500 150748
rect 40552 150736 40558 150748
rect 111334 150736 111340 150748
rect 40552 150708 111340 150736
rect 40552 150696 40558 150708
rect 111334 150696 111340 150708
rect 111392 150696 111398 150748
rect 36998 150628 37004 150680
rect 37056 150668 37062 150680
rect 111242 150668 111248 150680
rect 37056 150640 111248 150668
rect 37056 150628 37062 150640
rect 111242 150628 111248 150640
rect 111300 150628 111306 150680
rect 19794 150560 19800 150612
rect 19852 150600 19858 150612
rect 116854 150600 116860 150612
rect 19852 150572 116860 150600
rect 19852 150560 19858 150572
rect 116854 150560 116860 150572
rect 116912 150560 116918 150612
rect 16390 150492 16396 150544
rect 16448 150532 16454 150544
rect 116762 150532 116768 150544
rect 16448 150504 116768 150532
rect 16448 150492 16454 150504
rect 116762 150492 116768 150504
rect 116820 150492 116826 150544
rect 2682 150424 2688 150476
rect 2740 150464 2746 150476
rect 111058 150464 111064 150476
rect 2740 150436 111064 150464
rect 2740 150424 2746 150436
rect 111058 150424 111064 150436
rect 111116 150424 111122 150476
rect 118418 150152 118424 150204
rect 118476 150192 118482 150204
rect 121776 150192 121782 150204
rect 118476 150164 121782 150192
rect 118476 150152 118482 150164
rect 121776 150152 121782 150164
rect 121834 150152 121840 150204
rect 135438 150152 135444 150204
rect 135496 150192 135502 150204
rect 136588 150192 136594 150204
rect 135496 150164 136594 150192
rect 135496 150152 135502 150164
rect 136588 150152 136594 150164
rect 136646 150152 136652 150204
rect 146386 150152 146392 150204
rect 146444 150192 146450 150204
rect 147536 150192 147542 150204
rect 146444 150164 147542 150192
rect 146444 150152 146450 150164
rect 147536 150152 147542 150164
rect 147594 150152 147600 150204
rect 147674 150152 147680 150204
rect 147732 150192 147738 150204
rect 148824 150192 148830 150204
rect 147732 150164 148830 150192
rect 147732 150152 147738 150164
rect 148824 150152 148830 150164
rect 148882 150152 148888 150204
rect 164326 150152 164332 150204
rect 164384 150192 164390 150204
rect 165476 150192 165482 150204
rect 164384 150164 165482 150192
rect 164384 150152 164390 150164
rect 165476 150152 165482 150164
rect 165534 150152 165540 150204
rect 165614 150152 165620 150204
rect 165672 150192 165678 150204
rect 166764 150192 166770 150204
rect 165672 150164 166770 150192
rect 165672 150152 165678 150164
rect 166764 150152 166770 150164
rect 166822 150152 166828 150204
rect 171134 150152 171140 150204
rect 171192 150192 171198 150204
rect 171916 150192 171922 150204
rect 171192 150164 171922 150192
rect 171192 150152 171198 150164
rect 171916 150152 171922 150164
rect 171974 150152 171980 150204
rect 182266 150152 182272 150204
rect 182324 150192 182330 150204
rect 183416 150192 183422 150204
rect 182324 150164 183422 150192
rect 182324 150152 182330 150164
rect 183416 150152 183422 150164
rect 183474 150152 183480 150204
rect 183554 150152 183560 150204
rect 183612 150192 183618 150204
rect 184704 150192 184710 150204
rect 183612 150164 184710 150192
rect 183612 150152 183618 150164
rect 184704 150152 184710 150164
rect 184762 150152 184768 150204
rect 200298 150152 200304 150204
rect 200356 150192 200362 150204
rect 201448 150192 201454 150204
rect 200356 150164 201454 150192
rect 200356 150152 200362 150164
rect 201448 150152 201454 150164
rect 201506 150152 201512 150204
rect 204254 150152 204260 150204
rect 204312 150192 204318 150204
rect 205312 150192 205318 150204
rect 204312 150164 205318 150192
rect 204312 150152 204318 150164
rect 205312 150152 205318 150164
rect 205370 150152 205376 150204
rect 211246 150152 211252 150204
rect 211304 150192 211310 150204
rect 212304 150192 212310 150204
rect 211304 150164 212310 150192
rect 211304 150152 211310 150164
rect 212304 150152 212310 150164
rect 212362 150152 212368 150204
rect 218238 150152 218244 150204
rect 218296 150192 218302 150204
rect 219388 150192 219394 150204
rect 218296 150164 219394 150192
rect 218296 150152 218302 150164
rect 219388 150152 219394 150164
rect 219446 150152 219452 150204
rect 229186 150152 229192 150204
rect 229244 150192 229250 150204
rect 230336 150192 230342 150204
rect 229244 150164 230342 150192
rect 229244 150152 229250 150164
rect 230336 150152 230342 150164
rect 230394 150152 230400 150204
rect 238846 150152 238852 150204
rect 238904 150192 238910 150204
rect 239996 150192 240002 150204
rect 238904 150164 240002 150192
rect 238904 150152 238910 150164
rect 239996 150152 240002 150164
rect 240054 150152 240060 150204
rect 245838 150152 245844 150204
rect 245896 150192 245902 150204
rect 246988 150192 246994 150204
rect 245896 150164 246994 150192
rect 245896 150152 245902 150164
rect 246988 150152 246994 150164
rect 247046 150152 247052 150204
rect 247126 150152 247132 150204
rect 247184 150192 247190 150204
rect 248276 150192 248282 150204
rect 247184 150164 248282 150192
rect 247184 150152 247190 150164
rect 248276 150152 248282 150164
rect 248334 150152 248340 150204
rect 253934 150152 253940 150204
rect 253992 150192 253998 150204
rect 254716 150192 254722 150204
rect 253992 150164 254722 150192
rect 253992 150152 253998 150164
rect 254716 150152 254722 150164
rect 254774 150152 254780 150204
rect 256786 150152 256792 150204
rect 256844 150192 256850 150204
rect 257936 150192 257942 150204
rect 256844 150164 257942 150192
rect 256844 150152 256850 150164
rect 257936 150152 257942 150164
rect 257994 150152 258000 150204
rect 258074 150152 258080 150204
rect 258132 150192 258138 150204
rect 259224 150192 259230 150204
rect 258132 150164 259230 150192
rect 258132 150152 258138 150164
rect 259224 150152 259230 150164
rect 259282 150152 259288 150204
rect 259454 150152 259460 150204
rect 259512 150192 259518 150204
rect 260512 150192 260518 150204
rect 259512 150164 260518 150192
rect 259512 150152 259518 150164
rect 260512 150152 260518 150164
rect 260570 150152 260576 150204
rect 263594 150152 263600 150204
rect 263652 150192 263658 150204
rect 264376 150192 264382 150204
rect 263652 150164 264382 150192
rect 263652 150152 263658 150164
rect 264376 150152 264382 150164
rect 264434 150152 264440 150204
rect 281534 150152 281540 150204
rect 281592 150192 281598 150204
rect 282316 150192 282322 150204
rect 281592 150164 282322 150192
rect 281592 150152 281598 150164
rect 282316 150152 282322 150164
rect 282374 150152 282380 150204
rect 283098 150152 283104 150204
rect 283156 150192 283162 150204
rect 284248 150192 284254 150204
rect 283156 150164 284254 150192
rect 283156 150152 283162 150164
rect 284248 150152 284254 150164
rect 284306 150152 284312 150204
rect 285674 150152 285680 150204
rect 285732 150192 285738 150204
rect 286824 150192 286830 150204
rect 285732 150164 286830 150192
rect 285732 150152 285738 150164
rect 286824 150152 286830 150164
rect 286882 150152 286888 150204
rect 299474 150152 299480 150204
rect 299532 150192 299538 150204
rect 300348 150192 300354 150204
rect 299532 150164 300354 150192
rect 299532 150152 299538 150164
rect 300348 150152 300354 150164
rect 300406 150152 300412 150204
rect 302418 150152 302424 150204
rect 302476 150192 302482 150204
rect 303568 150192 303574 150204
rect 302476 150164 303574 150192
rect 302476 150152 302482 150164
rect 303568 150152 303574 150164
rect 303626 150152 303632 150204
rect 347958 150152 347964 150204
rect 348016 150192 348022 150204
rect 349108 150192 349114 150204
rect 348016 150164 349114 150192
rect 348016 150152 348022 150164
rect 349108 150152 349114 150164
rect 349166 150152 349172 150204
rect 354674 150152 354680 150204
rect 354732 150192 354738 150204
rect 355548 150192 355554 150204
rect 354732 150164 355554 150192
rect 354732 150152 354738 150164
rect 355548 150152 355554 150164
rect 355606 150152 355612 150204
rect 358906 150152 358912 150204
rect 358964 150192 358970 150204
rect 360056 150192 360062 150204
rect 358964 150164 360062 150192
rect 358964 150152 358970 150164
rect 360056 150152 360062 150164
rect 360114 150152 360120 150204
rect 369854 150152 369860 150204
rect 369912 150192 369918 150204
rect 370912 150192 370918 150204
rect 369912 150164 370918 150192
rect 369912 150152 369918 150164
rect 370912 150152 370918 150164
rect 370970 150152 370976 150204
rect 375558 150152 375564 150204
rect 375616 150192 375622 150204
rect 376708 150192 376714 150204
rect 375616 150164 376714 150192
rect 375616 150152 375622 150164
rect 376708 150152 376714 150164
rect 376766 150152 376772 150204
rect 378134 150152 378140 150204
rect 378192 150192 378198 150204
rect 379284 150192 379290 150204
rect 378192 150164 379290 150192
rect 378192 150152 378198 150164
rect 379284 150152 379290 150164
rect 379342 150152 379348 150204
rect 394878 150152 394884 150204
rect 394936 150192 394942 150204
rect 396028 150192 396034 150204
rect 394936 150164 396034 150192
rect 394936 150152 394942 150164
rect 396028 150152 396034 150164
rect 396086 150152 396092 150204
rect 403158 150152 403164 150204
rect 403216 150192 403222 150204
rect 404308 150192 404314 150204
rect 403216 150164 404314 150192
rect 403216 150152 403222 150164
rect 404308 150152 404314 150164
rect 404366 150152 404372 150204
rect 477678 150152 477684 150204
rect 477736 150192 477742 150204
rect 478828 150192 478834 150204
rect 477736 150164 478834 150192
rect 477736 150152 477742 150164
rect 478828 150152 478834 150164
rect 478886 150152 478892 150204
rect 478966 150152 478972 150204
rect 479024 150192 479030 150204
rect 480116 150192 480122 150204
rect 479024 150164 480122 150192
rect 479024 150152 479030 150164
rect 480116 150152 480122 150164
rect 480174 150152 480180 150204
rect 481634 150152 481640 150204
rect 481692 150192 481698 150204
rect 482692 150192 482698 150204
rect 481692 150164 482698 150192
rect 481692 150152 481698 150164
rect 482692 150152 482698 150164
rect 482750 150152 482756 150204
rect 6362 150016 6368 150068
rect 6420 150056 6426 150068
rect 111150 150056 111156 150068
rect 6420 150028 111156 150056
rect 6420 150016 6426 150028
rect 111150 150016 111156 150028
rect 111208 150016 111214 150068
rect 23382 149948 23388 150000
rect 23440 149988 23446 150000
rect 116946 149988 116952 150000
rect 23440 149960 116952 149988
rect 23440 149948 23446 149960
rect 116946 149948 116952 149960
rect 117004 149948 117010 150000
rect 13354 149880 13360 149932
rect 13412 149920 13418 149932
rect 116670 149920 116676 149932
rect 13412 149892 116676 149920
rect 13412 149880 13418 149892
rect 116670 149880 116676 149892
rect 116728 149880 116734 149932
rect 9582 149812 9588 149864
rect 9640 149852 9646 149864
rect 116578 149852 116584 149864
rect 9640 149824 116584 149852
rect 9640 149812 9646 149824
rect 116578 149812 116584 149824
rect 116636 149812 116642 149864
rect 88978 149744 88984 149796
rect 89036 149784 89042 149796
rect 114002 149784 114008 149796
rect 89036 149756 114008 149784
rect 89036 149744 89042 149756
rect 114002 149744 114008 149756
rect 114060 149744 114066 149796
rect 85482 149676 85488 149728
rect 85540 149716 85546 149728
rect 113910 149716 113916 149728
rect 85540 149688 113916 149716
rect 85540 149676 85546 149688
rect 113910 149676 113916 149688
rect 113968 149676 113974 149728
rect 81986 149608 81992 149660
rect 82044 149648 82050 149660
rect 112346 149648 112352 149660
rect 82044 149620 112352 149648
rect 82044 149608 82050 149620
rect 112346 149608 112352 149620
rect 112404 149608 112410 149660
rect 78582 149540 78588 149592
rect 78640 149580 78646 149592
rect 113082 149580 113088 149592
rect 78640 149552 113088 149580
rect 78640 149540 78646 149552
rect 113082 149540 113088 149552
rect 113140 149540 113146 149592
rect 75178 149472 75184 149524
rect 75236 149512 75242 149524
rect 112990 149512 112996 149524
rect 75236 149484 112996 149512
rect 75236 149472 75242 149484
rect 112990 149472 112996 149484
rect 113048 149472 113054 149524
rect 71682 149404 71688 149456
rect 71740 149444 71746 149456
rect 112898 149444 112904 149456
rect 71740 149416 112904 149444
rect 71740 149404 71746 149416
rect 112898 149404 112904 149416
rect 112956 149404 112962 149456
rect 26970 149336 26976 149388
rect 27028 149376 27034 149388
rect 117038 149376 117044 149388
rect 27028 149348 117044 149376
rect 27028 149336 27034 149348
rect 117038 149336 117044 149348
rect 117096 149336 117102 149388
rect 92290 149268 92296 149320
rect 92348 149308 92354 149320
rect 92348 149280 93854 149308
rect 92348 149268 92354 149280
rect 93826 149104 93854 149280
rect 102502 149268 102508 149320
rect 102560 149268 102566 149320
rect 102686 149268 102692 149320
rect 102744 149268 102750 149320
rect 102870 149268 102876 149320
rect 102928 149308 102934 149320
rect 116210 149308 116216 149320
rect 102928 149280 116216 149308
rect 102928 149268 102934 149280
rect 116210 149268 116216 149280
rect 116268 149268 116274 149320
rect 102520 149172 102548 149268
rect 102704 149240 102732 149268
rect 116486 149240 116492 149252
rect 102704 149212 116492 149240
rect 116486 149200 116492 149212
rect 116544 149200 116550 149252
rect 116026 149172 116032 149184
rect 102520 149144 116032 149172
rect 116026 149132 116032 149144
rect 116084 149132 116090 149184
rect 114094 149104 114100 149116
rect 93826 149076 96614 149104
rect 96586 148764 96614 149076
rect 106246 149076 114100 149104
rect 106246 148764 106274 149076
rect 114094 149064 114100 149076
rect 114152 149064 114158 149116
rect 109586 148996 109592 149048
rect 109644 149036 109650 149048
rect 115934 149036 115940 149048
rect 109644 149008 115940 149036
rect 109644 148996 109650 149008
rect 115934 148996 115940 149008
rect 115992 148996 115998 149048
rect 96586 148736 106274 148764
rect 110322 147568 110328 147620
rect 110380 147608 110386 147620
rect 116118 147608 116124 147620
rect 110380 147580 116124 147608
rect 110380 147568 110386 147580
rect 116118 147568 116124 147580
rect 116176 147568 116182 147620
rect 114094 140700 114100 140752
rect 114152 140740 114158 140752
rect 115934 140740 115940 140752
rect 114152 140712 115940 140740
rect 114152 140700 114158 140712
rect 115934 140700 115940 140712
rect 115992 140700 115998 140752
rect 114002 137912 114008 137964
rect 114060 137952 114066 137964
rect 116394 137952 116400 137964
rect 114060 137924 116400 137952
rect 114060 137912 114066 137924
rect 116394 137912 116400 137924
rect 116452 137912 116458 137964
rect 113910 136552 113916 136604
rect 113968 136592 113974 136604
rect 115934 136592 115940 136604
rect 113968 136564 115940 136592
rect 113968 136552 113974 136564
rect 115934 136552 115940 136564
rect 115992 136552 115998 136604
rect 112346 133832 112352 133884
rect 112404 133872 112410 133884
rect 116118 133872 116124 133884
rect 112404 133844 116124 133872
rect 112404 133832 112410 133844
rect 116118 133832 116124 133844
rect 116176 133832 116182 133884
rect 113082 132404 113088 132456
rect 113140 132444 113146 132456
rect 116118 132444 116124 132456
rect 113140 132416 116124 132444
rect 113140 132404 113146 132416
rect 116118 132404 116124 132416
rect 116176 132404 116182 132456
rect 112990 131044 112996 131096
rect 113048 131084 113054 131096
rect 116118 131084 116124 131096
rect 113048 131056 116124 131084
rect 113048 131044 113054 131056
rect 116118 131044 116124 131056
rect 116176 131044 116182 131096
rect 112898 128256 112904 128308
rect 112956 128296 112962 128308
rect 116118 128296 116124 128308
rect 112956 128268 116124 128296
rect 112956 128256 112962 128268
rect 116118 128256 116124 128268
rect 116176 128256 116182 128308
rect 112806 126896 112812 126948
rect 112864 126936 112870 126948
rect 116026 126936 116032 126948
rect 112864 126908 116032 126936
rect 112864 126896 112870 126908
rect 116026 126896 116032 126908
rect 116084 126896 116090 126948
rect 112714 124108 112720 124160
rect 112772 124148 112778 124160
rect 116118 124148 116124 124160
rect 112772 124120 116124 124148
rect 112772 124108 112778 124120
rect 116118 124108 116124 124120
rect 116176 124108 116182 124160
rect 112622 122748 112628 122800
rect 112680 122788 112686 122800
rect 115934 122788 115940 122800
rect 112680 122760 115940 122788
rect 112680 122748 112686 122760
rect 115934 122748 115940 122760
rect 115992 122748 115998 122800
rect 112530 121388 112536 121440
rect 112588 121428 112594 121440
rect 116118 121428 116124 121440
rect 112588 121400 116124 121428
rect 112588 121388 112594 121400
rect 116118 121388 116124 121400
rect 116176 121388 116182 121440
rect 111610 118600 111616 118652
rect 111668 118640 111674 118652
rect 116118 118640 116124 118652
rect 111668 118612 116124 118640
rect 111668 118600 111674 118612
rect 116118 118600 116124 118612
rect 116176 118600 116182 118652
rect 116486 117988 116492 118040
rect 116544 118028 116550 118040
rect 117222 118028 117228 118040
rect 116544 118000 117228 118028
rect 116544 117988 116550 118000
rect 117222 117988 117228 118000
rect 117280 117988 117286 118040
rect 112438 117240 112444 117292
rect 112496 117280 112502 117292
rect 116118 117280 116124 117292
rect 112496 117252 116124 117280
rect 112496 117240 112502 117252
rect 116118 117240 116124 117252
rect 116176 117240 116182 117292
rect 111518 114452 111524 114504
rect 111576 114492 111582 114504
rect 116118 114492 116124 114504
rect 111576 114464 116124 114492
rect 111576 114452 111582 114464
rect 116118 114452 116124 114464
rect 116176 114452 116182 114504
rect 111426 113092 111432 113144
rect 111484 113132 111490 113144
rect 115934 113132 115940 113144
rect 111484 113104 115940 113132
rect 111484 113092 111490 113104
rect 115934 113092 115940 113104
rect 115992 113092 115998 113144
rect 111334 111732 111340 111784
rect 111392 111772 111398 111784
rect 116118 111772 116124 111784
rect 111392 111744 116124 111772
rect 111392 111732 111398 111744
rect 116118 111732 116124 111744
rect 116176 111732 116182 111784
rect 111242 108944 111248 108996
rect 111300 108984 111306 108996
rect 116118 108984 116124 108996
rect 111300 108956 116124 108984
rect 111300 108944 111306 108956
rect 116118 108944 116124 108956
rect 116176 108944 116182 108996
rect 111150 92420 111156 92472
rect 111208 92460 111214 92472
rect 116118 92460 116124 92472
rect 111208 92432 116124 92460
rect 111208 92420 111214 92432
rect 116118 92420 116124 92432
rect 116176 92420 116182 92472
rect 111058 89632 111064 89684
rect 111116 89672 111122 89684
rect 116118 89672 116124 89684
rect 111116 89644 116124 89672
rect 111116 89632 111122 89644
rect 116118 89632 116124 89644
rect 116176 89632 116182 89684
rect 113818 88272 113824 88324
rect 113876 88312 113882 88324
rect 116026 88312 116032 88324
rect 113876 88284 116032 88312
rect 113876 88272 113882 88284
rect 116026 88272 116032 88284
rect 116084 88272 116090 88324
rect 114462 87184 114468 87236
rect 114520 87224 114526 87236
rect 116486 87224 116492 87236
rect 114520 87196 116492 87224
rect 114520 87184 114526 87196
rect 116486 87184 116492 87196
rect 116544 87184 116550 87236
rect 113910 86912 113916 86964
rect 113968 86952 113974 86964
rect 116210 86952 116216 86964
rect 113968 86924 116216 86952
rect 113968 86912 113974 86924
rect 116210 86912 116216 86924
rect 116268 86912 116274 86964
rect 114002 83920 114008 83972
rect 114060 83960 114066 83972
rect 116578 83960 116584 83972
rect 114060 83932 116584 83960
rect 114060 83920 114066 83932
rect 116578 83920 116584 83932
rect 116636 83920 116642 83972
rect 114094 82764 114100 82816
rect 114152 82804 114158 82816
rect 116302 82804 116308 82816
rect 114152 82776 116308 82804
rect 114152 82764 114158 82776
rect 116302 82764 116308 82776
rect 116360 82764 116366 82816
rect 114186 79976 114192 80028
rect 114244 80016 114250 80028
rect 115934 80016 115940 80028
rect 114244 79988 115940 80016
rect 114244 79976 114250 79988
rect 115934 79976 115940 79988
rect 115992 79976 115998 80028
rect 114186 71748 114192 71800
rect 114244 71788 114250 71800
rect 116578 71788 116584 71800
rect 114244 71760 116584 71788
rect 114244 71748 114250 71760
rect 116578 71748 116584 71760
rect 116636 71748 116642 71800
rect 114094 69028 114100 69080
rect 114152 69068 114158 69080
rect 116302 69068 116308 69080
rect 114152 69040 116308 69068
rect 114152 69028 114158 69040
rect 116302 69028 116308 69040
rect 116360 69028 116366 69080
rect 114002 67600 114008 67652
rect 114060 67640 114066 67652
rect 116118 67640 116124 67652
rect 114060 67612 116124 67640
rect 114060 67600 114066 67612
rect 116118 67600 116124 67612
rect 116176 67600 116182 67652
rect 113910 66240 113916 66292
rect 113968 66280 113974 66292
rect 116578 66280 116584 66292
rect 113968 66252 116584 66280
rect 113968 66240 113974 66252
rect 116578 66240 116584 66252
rect 116636 66240 116642 66292
rect 114462 64540 114468 64592
rect 114520 64580 114526 64592
rect 116578 64580 116584 64592
rect 114520 64552 116584 64580
rect 114520 64540 114526 64552
rect 116578 64540 116584 64552
rect 116636 64540 116642 64592
rect 113818 63520 113824 63572
rect 113876 63560 113882 63572
rect 116210 63560 116216 63572
rect 113876 63532 116216 63560
rect 113876 63520 113882 63532
rect 116210 63520 116216 63532
rect 116268 63520 116274 63572
rect 109678 41420 109684 41472
rect 109736 41460 109742 41472
rect 116118 41460 116124 41472
rect 109736 41432 116124 41460
rect 109736 41420 109742 41432
rect 116118 41420 116124 41432
rect 116176 41420 116182 41472
rect 114094 38632 114100 38684
rect 114152 38672 114158 38684
rect 116394 38672 116400 38684
rect 114152 38644 116400 38672
rect 114152 38632 114158 38644
rect 116394 38632 116400 38644
rect 116452 38632 116458 38684
rect 116210 38496 116216 38548
rect 116268 38536 116274 38548
rect 116394 38536 116400 38548
rect 116268 38508 116400 38536
rect 116268 38496 116274 38508
rect 116394 38496 116400 38508
rect 116452 38496 116458 38548
rect 114186 37272 114192 37324
rect 114244 37312 114250 37324
rect 116210 37312 116216 37324
rect 114244 37284 116216 37312
rect 114244 37272 114250 37284
rect 116210 37272 116216 37284
rect 116268 37272 116274 37324
rect 111058 34484 111064 34536
rect 111116 34524 111122 34536
rect 116118 34524 116124 34536
rect 111116 34496 116124 34524
rect 111116 34484 111122 34496
rect 116118 34484 116124 34496
rect 116176 34484 116182 34536
rect 112438 33124 112444 33176
rect 112496 33164 112502 33176
rect 116118 33164 116124 33176
rect 112496 33136 116124 33164
rect 112496 33124 112502 33136
rect 116118 33124 116124 33136
rect 116176 33124 116182 33176
rect 112530 31764 112536 31816
rect 112588 31804 112594 31816
rect 116118 31804 116124 31816
rect 112588 31776 116124 31804
rect 112588 31764 112594 31776
rect 116118 31764 116124 31776
rect 116176 31764 116182 31816
rect 112622 28976 112628 29028
rect 112680 29016 112686 29028
rect 116118 29016 116124 29028
rect 112680 28988 116124 29016
rect 112680 28976 112686 28988
rect 116118 28976 116124 28988
rect 116176 28976 116182 29028
rect 112714 27616 112720 27668
rect 112772 27656 112778 27668
rect 116118 27656 116124 27668
rect 112772 27628 116124 27656
rect 112772 27616 112778 27628
rect 116118 27616 116124 27628
rect 116176 27616 116182 27668
rect 112806 24828 112812 24880
rect 112864 24868 112870 24880
rect 116118 24868 116124 24880
rect 112864 24840 116124 24868
rect 112864 24828 112870 24840
rect 116118 24828 116124 24840
rect 116176 24828 116182 24880
rect 111150 23468 111156 23520
rect 111208 23508 111214 23520
rect 116118 23508 116124 23520
rect 111208 23480 116124 23508
rect 111208 23468 111214 23480
rect 116118 23468 116124 23480
rect 116176 23468 116182 23520
rect 111242 22108 111248 22160
rect 111300 22148 111306 22160
rect 116026 22148 116032 22160
rect 111300 22120 116032 22148
rect 111300 22108 111306 22120
rect 116026 22108 116032 22120
rect 116084 22108 116090 22160
rect 116026 16464 116032 16516
rect 116084 16504 116090 16516
rect 116210 16504 116216 16516
rect 116084 16476 116216 16504
rect 116084 16464 116090 16476
rect 116210 16464 116216 16476
rect 116268 16464 116274 16516
rect 116210 11840 116216 11892
rect 116268 11840 116274 11892
rect 116228 11676 116256 11840
rect 116302 11676 116308 11688
rect 116228 11648 116308 11676
rect 116302 11636 116308 11648
rect 116360 11636 116366 11688
rect 116946 11364 116952 11416
rect 117004 11404 117010 11416
rect 117314 11404 117320 11416
rect 117004 11376 117320 11404
rect 117004 11364 117010 11376
rect 117314 11364 117320 11376
rect 117372 11364 117378 11416
rect 116946 5448 116952 5500
rect 117004 5488 117010 5500
rect 117130 5488 117136 5500
rect 117004 5460 117136 5488
rect 117004 5448 117010 5460
rect 117130 5448 117136 5460
rect 117188 5448 117194 5500
rect 116302 5312 116308 5364
rect 116360 5352 116366 5364
rect 116946 5352 116952 5364
rect 116360 5324 116952 5352
rect 116360 5312 116366 5324
rect 116946 5312 116952 5324
rect 117004 5312 117010 5364
rect 115934 5176 115940 5228
rect 115992 5216 115998 5228
rect 116302 5216 116308 5228
rect 115992 5188 116308 5216
rect 115992 5176 115998 5188
rect 116302 5176 116308 5188
rect 116360 5176 116366 5228
rect 115934 5040 115940 5092
rect 115992 5080 115998 5092
rect 116118 5080 116124 5092
rect 115992 5052 116124 5080
rect 115992 5040 115998 5052
rect 116118 5040 116124 5052
rect 116176 5040 116182 5092
rect 109770 4156 109776 4208
rect 109828 4196 109834 4208
rect 116118 4196 116124 4208
rect 109828 4168 116124 4196
rect 109828 4156 109834 4168
rect 116118 4156 116124 4168
rect 116176 4156 116182 4208
rect 111058 3924 111064 3936
rect 75886 3896 111064 3924
rect 71746 3828 73154 3856
rect 62776 3692 63172 3720
rect 53208 3624 62620 3652
rect 39684 3488 48314 3516
rect 32784 3080 38654 3108
rect 26206 3012 28994 3040
rect 2498 2864 2504 2916
rect 2556 2904 2562 2916
rect 26206 2904 26234 3012
rect 2556 2876 26234 2904
rect 2556 2864 2562 2876
rect 28966 2564 28994 3012
rect 32784 2644 32812 3080
rect 32766 2592 32772 2644
rect 32824 2592 32830 2644
rect 38626 2632 38654 3080
rect 39684 2644 39712 3488
rect 40328 3420 47532 3448
rect 40328 2644 40356 3420
rect 47504 2644 47532 3420
rect 39114 2632 39120 2644
rect 38626 2604 39120 2632
rect 39114 2592 39120 2604
rect 39172 2592 39178 2644
rect 39666 2592 39672 2644
rect 39724 2592 39730 2644
rect 40310 2592 40316 2644
rect 40368 2592 40374 2644
rect 47486 2592 47492 2644
rect 47544 2592 47550 2644
rect 48286 2632 48314 3488
rect 53208 2700 53236 3624
rect 49620 2672 53236 2700
rect 53300 3556 58756 3584
rect 49620 2644 49648 2672
rect 49142 2632 49148 2644
rect 48286 2604 49148 2632
rect 49142 2592 49148 2604
rect 49200 2592 49206 2644
rect 49602 2592 49608 2644
rect 49660 2592 49666 2644
rect 50890 2592 50896 2644
rect 50948 2632 50954 2644
rect 53006 2632 53012 2644
rect 50948 2604 53012 2632
rect 50948 2592 50954 2604
rect 53006 2592 53012 2604
rect 53064 2592 53070 2644
rect 28966 2536 42932 2564
rect 36354 2456 36360 2508
rect 36412 2496 36418 2508
rect 40310 2496 40316 2508
rect 36412 2468 40316 2496
rect 36412 2456 36418 2468
rect 40310 2456 40316 2468
rect 40368 2456 40374 2508
rect 42904 2496 42932 2536
rect 46290 2524 46296 2576
rect 46348 2564 46354 2576
rect 53300 2564 53328 3556
rect 53484 2944 58664 2972
rect 53484 2644 53512 2944
rect 58636 2644 58664 2944
rect 58728 2644 58756 3556
rect 62592 3244 62620 3624
rect 62408 3216 62620 3244
rect 62408 2644 62436 3216
rect 62776 2644 62804 3692
rect 63144 3652 63172 3692
rect 63144 3624 63494 3652
rect 63466 3516 63494 3624
rect 67284 3556 67496 3584
rect 63466 3488 64874 3516
rect 64846 3312 64874 3488
rect 67284 3380 67312 3556
rect 67468 3516 67496 3556
rect 67606 3556 70394 3584
rect 67606 3516 67634 3556
rect 67468 3488 67634 3516
rect 70366 3516 70394 3556
rect 71746 3516 71774 3828
rect 73126 3788 73154 3828
rect 73126 3760 74534 3788
rect 74506 3584 74534 3760
rect 75886 3584 75914 3896
rect 111058 3884 111064 3896
rect 111116 3884 111122 3936
rect 112438 3856 112444 3868
rect 74506 3556 75914 3584
rect 77956 3828 112444 3856
rect 70366 3488 71774 3516
rect 68986 3420 70394 3448
rect 68986 3380 69014 3420
rect 66226 3352 67312 3380
rect 67606 3352 69014 3380
rect 70366 3380 70394 3420
rect 74506 3420 75914 3448
rect 74506 3380 74534 3420
rect 70366 3352 71774 3380
rect 66226 3312 66254 3352
rect 64846 3284 66254 3312
rect 64156 3216 64736 3244
rect 64156 3108 64184 3216
rect 64708 3176 64736 3216
rect 64846 3216 66254 3244
rect 64846 3176 64874 3216
rect 64708 3148 64874 3176
rect 66226 3176 66254 3216
rect 67606 3176 67634 3352
rect 71746 3312 71774 3352
rect 73126 3352 74534 3380
rect 75886 3380 75914 3420
rect 75886 3352 77294 3380
rect 73126 3312 73154 3352
rect 71746 3284 73154 3312
rect 66226 3148 67634 3176
rect 63466 3080 64184 3108
rect 77266 3108 77294 3352
rect 77956 3176 77984 3828
rect 112438 3816 112444 3828
rect 112496 3816 112502 3868
rect 112530 3788 112536 3800
rect 78508 3760 112536 3788
rect 77956 3148 78260 3176
rect 77266 3080 78168 3108
rect 63466 2768 63494 3080
rect 63052 2740 63494 2768
rect 73126 2808 78076 2836
rect 63052 2644 63080 2740
rect 73126 2700 73154 2808
rect 63144 2672 73154 2700
rect 63144 2644 63172 2672
rect 78048 2644 78076 2808
rect 78140 2644 78168 3080
rect 53466 2592 53472 2644
rect 53524 2592 53530 2644
rect 53650 2592 53656 2644
rect 53708 2632 53714 2644
rect 57514 2632 57520 2644
rect 53708 2604 57520 2632
rect 53708 2592 53714 2604
rect 57514 2592 57520 2604
rect 57572 2592 57578 2644
rect 58618 2592 58624 2644
rect 58676 2592 58682 2644
rect 58710 2592 58716 2644
rect 58768 2592 58774 2644
rect 62390 2592 62396 2644
rect 62448 2592 62454 2644
rect 62758 2592 62764 2644
rect 62816 2592 62822 2644
rect 63034 2592 63040 2644
rect 63092 2592 63098 2644
rect 63126 2592 63132 2644
rect 63184 2592 63190 2644
rect 65518 2592 65524 2644
rect 65576 2632 65582 2644
rect 65576 2604 76788 2632
rect 65576 2592 65582 2604
rect 46348 2536 53328 2564
rect 46348 2524 46354 2536
rect 56226 2524 56232 2576
rect 56284 2564 56290 2576
rect 73982 2564 73988 2576
rect 56284 2536 73988 2564
rect 56284 2524 56290 2536
rect 73982 2524 73988 2536
rect 74040 2524 74046 2576
rect 74074 2524 74080 2576
rect 74132 2564 74138 2576
rect 76650 2564 76656 2576
rect 74132 2536 76656 2564
rect 74132 2524 74138 2536
rect 76650 2524 76656 2536
rect 76708 2524 76714 2576
rect 76760 2564 76788 2604
rect 78030 2592 78036 2644
rect 78088 2592 78094 2644
rect 78122 2592 78128 2644
rect 78180 2592 78186 2644
rect 78232 2564 78260 3148
rect 78508 2644 78536 3760
rect 112530 3748 112536 3760
rect 112588 3748 112594 3800
rect 112622 3720 112628 3732
rect 79704 3692 112628 3720
rect 79704 2644 79732 3692
rect 112622 3680 112628 3692
rect 112680 3680 112686 3732
rect 112714 3652 112720 3664
rect 81084 3624 112720 3652
rect 81084 3516 81112 3624
rect 112714 3612 112720 3624
rect 112772 3612 112778 3664
rect 112806 3584 112812 3596
rect 79796 3488 81112 3516
rect 81176 3556 112812 3584
rect 79796 2644 79824 3488
rect 81176 2644 81204 3556
rect 112806 3544 112812 3556
rect 112864 3544 112870 3596
rect 111150 3516 111156 3528
rect 81820 3488 82124 3516
rect 81820 3448 81848 3488
rect 81636 3420 81848 3448
rect 81636 3380 81664 3420
rect 81268 3352 81664 3380
rect 82096 3380 82124 3488
rect 82372 3488 111156 3516
rect 82372 3380 82400 3488
rect 111150 3476 111156 3488
rect 111208 3476 111214 3528
rect 111242 3448 111248 3460
rect 82096 3352 82400 3380
rect 82464 3420 111248 3448
rect 81268 2644 81296 3352
rect 82464 3312 82492 3420
rect 111242 3408 111248 3420
rect 111300 3408 111306 3460
rect 114186 3380 114192 3392
rect 82280 3284 82492 3312
rect 82786 3352 114192 3380
rect 81360 3216 82124 3244
rect 81360 2644 81388 3216
rect 82096 3176 82124 3216
rect 82280 3176 82308 3284
rect 82786 3244 82814 3352
rect 114186 3340 114192 3352
rect 114244 3340 114250 3392
rect 114094 3312 114100 3324
rect 82096 3148 82308 3176
rect 82372 3216 82814 3244
rect 84166 3284 114100 3312
rect 82372 3108 82400 3216
rect 84166 3176 84194 3284
rect 114094 3272 114100 3284
rect 114152 3272 114158 3324
rect 82556 3148 84194 3176
rect 96586 3148 104894 3176
rect 82556 3108 82584 3148
rect 96586 3108 96614 3148
rect 82096 3080 82400 3108
rect 82464 3080 82584 3108
rect 82786 3080 96614 3108
rect 82096 2644 82124 3080
rect 82464 2972 82492 3080
rect 82786 2972 82814 3080
rect 101508 3012 104296 3040
rect 101508 2972 101536 3012
rect 82188 2944 82492 2972
rect 82556 2944 82814 2972
rect 89686 2944 101536 2972
rect 82188 2644 82216 2944
rect 78490 2592 78496 2644
rect 78548 2592 78554 2644
rect 79686 2592 79692 2644
rect 79744 2592 79750 2644
rect 79778 2592 79784 2644
rect 79836 2592 79842 2644
rect 81158 2592 81164 2644
rect 81216 2592 81222 2644
rect 81250 2592 81256 2644
rect 81308 2592 81314 2644
rect 81342 2592 81348 2644
rect 81400 2592 81406 2644
rect 82078 2592 82084 2644
rect 82136 2592 82142 2644
rect 82170 2592 82176 2644
rect 82228 2592 82234 2644
rect 82262 2592 82268 2644
rect 82320 2632 82326 2644
rect 82556 2632 82584 2944
rect 89686 2904 89714 2944
rect 82320 2604 82584 2632
rect 82786 2876 89714 2904
rect 96586 2876 98224 2904
rect 82320 2592 82326 2604
rect 76760 2536 78260 2564
rect 79410 2524 79416 2576
rect 79468 2524 79474 2576
rect 79594 2524 79600 2576
rect 79652 2564 79658 2576
rect 82786 2564 82814 2876
rect 96586 2836 96614 2876
rect 79652 2536 82814 2564
rect 84166 2808 96614 2836
rect 79652 2524 79658 2536
rect 79428 2496 79456 2524
rect 42904 2468 79456 2496
rect 52914 2388 52920 2440
rect 52972 2428 52978 2440
rect 53650 2428 53656 2440
rect 52972 2400 53656 2428
rect 52972 2388 52978 2400
rect 53650 2388 53656 2400
rect 53708 2388 53714 2440
rect 59722 2388 59728 2440
rect 59780 2428 59786 2440
rect 65518 2428 65524 2440
rect 59780 2400 65524 2428
rect 59780 2388 59786 2400
rect 65518 2388 65524 2400
rect 65576 2388 65582 2440
rect 66346 2388 66352 2440
rect 66404 2428 66410 2440
rect 82078 2428 82084 2440
rect 66404 2400 82084 2428
rect 66404 2388 66410 2400
rect 82078 2388 82084 2400
rect 82136 2388 82142 2440
rect 81158 2360 81164 2372
rect 53484 2332 81164 2360
rect 53006 2252 53012 2304
rect 53064 2292 53070 2304
rect 53484 2292 53512 2332
rect 81158 2320 81164 2332
rect 81216 2320 81222 2372
rect 76558 2292 76564 2304
rect 53064 2264 53512 2292
rect 53576 2264 76564 2292
rect 53064 2252 53070 2264
rect 47486 2184 47492 2236
rect 47544 2224 47550 2236
rect 53576 2224 53604 2264
rect 76558 2252 76564 2264
rect 76616 2252 76622 2304
rect 76650 2252 76656 2304
rect 76708 2292 76714 2304
rect 84166 2292 84194 2808
rect 98196 2564 98224 2876
rect 104268 2768 104296 3012
rect 104866 2972 104894 3148
rect 109586 3000 109592 3052
rect 109644 3040 109650 3052
rect 117958 3040 117964 3052
rect 109644 3012 117964 3040
rect 109644 3000 109650 3012
rect 117958 3000 117964 3012
rect 118016 3000 118022 3052
rect 117682 2972 117688 2984
rect 104866 2944 117688 2972
rect 117682 2932 117688 2944
rect 117740 2932 117746 2984
rect 116118 2904 116124 2916
rect 104866 2876 116124 2904
rect 104866 2836 104894 2876
rect 116118 2864 116124 2876
rect 116176 2864 116182 2916
rect 104360 2808 104894 2836
rect 106246 2808 294736 2836
rect 104360 2768 104388 2808
rect 104268 2740 104388 2768
rect 98270 2592 98276 2644
rect 98328 2632 98334 2644
rect 106090 2632 106096 2644
rect 98328 2604 106096 2632
rect 98328 2592 98334 2604
rect 106090 2592 106096 2604
rect 106148 2592 106154 2644
rect 106246 2564 106274 2808
rect 294708 2632 294736 2808
rect 425808 2808 443684 2836
rect 425808 2644 425836 2808
rect 443656 2644 443684 2808
rect 491312 2808 493640 2836
rect 491312 2644 491340 2808
rect 493612 2644 493640 2808
rect 294782 2632 294788 2644
rect 294708 2604 294788 2632
rect 294782 2592 294788 2604
rect 294840 2592 294846 2644
rect 425790 2592 425796 2644
rect 425848 2592 425854 2644
rect 443638 2592 443644 2644
rect 443696 2592 443702 2644
rect 491294 2592 491300 2644
rect 491352 2592 491358 2644
rect 493594 2592 493600 2644
rect 493652 2592 493658 2644
rect 98196 2536 106274 2564
rect 109586 2456 109592 2508
rect 109644 2496 109650 2508
rect 116578 2496 116584 2508
rect 109644 2468 116584 2496
rect 109644 2456 109650 2468
rect 116578 2456 116584 2468
rect 116636 2456 116642 2508
rect 106182 2388 106188 2440
rect 106240 2428 106246 2440
rect 116670 2428 116676 2440
rect 106240 2400 116676 2428
rect 106240 2388 106246 2400
rect 116670 2388 116676 2400
rect 116728 2388 116734 2440
rect 102962 2320 102968 2372
rect 103020 2360 103026 2372
rect 116762 2360 116768 2372
rect 103020 2332 116768 2360
rect 103020 2320 103026 2332
rect 116762 2320 116768 2332
rect 116820 2320 116826 2372
rect 76708 2264 84194 2292
rect 76708 2252 76714 2264
rect 99650 2252 99656 2304
rect 99708 2292 99714 2304
rect 116854 2292 116860 2304
rect 99708 2264 116860 2292
rect 99708 2252 99714 2264
rect 116854 2252 116860 2264
rect 116912 2252 116918 2304
rect 47544 2196 53604 2224
rect 47544 2184 47550 2196
rect 58710 2184 58716 2236
rect 58768 2224 58774 2236
rect 63126 2224 63132 2236
rect 58768 2196 63132 2224
rect 58768 2184 58774 2196
rect 63126 2184 63132 2196
rect 63184 2184 63190 2236
rect 69658 2184 69664 2236
rect 69716 2224 69722 2236
rect 82170 2224 82176 2236
rect 69716 2196 82176 2224
rect 69716 2184 69722 2196
rect 82170 2184 82176 2196
rect 82228 2184 82234 2236
rect 96338 2184 96344 2236
rect 96396 2224 96402 2236
rect 117038 2224 117044 2236
rect 96396 2196 117044 2224
rect 96396 2184 96402 2196
rect 117038 2184 117044 2196
rect 117096 2184 117102 2236
rect 57514 2116 57520 2168
rect 57572 2156 57578 2168
rect 57572 2128 63494 2156
rect 57572 2116 57578 2128
rect 63466 2088 63494 2128
rect 76558 2116 76564 2168
rect 76616 2156 76622 2168
rect 81342 2156 81348 2168
rect 76616 2128 81348 2156
rect 76616 2116 76622 2128
rect 81342 2116 81348 2128
rect 81400 2116 81406 2168
rect 93026 2116 93032 2168
rect 93084 2156 93090 2168
rect 117222 2156 117228 2168
rect 93084 2128 117228 2156
rect 93084 2116 93090 2128
rect 117222 2116 117228 2128
rect 117280 2116 117286 2168
rect 78490 2088 78496 2100
rect 63466 2060 78496 2088
rect 78490 2048 78496 2060
rect 78548 2048 78554 2100
rect 89622 2048 89628 2100
rect 89680 2088 89686 2100
rect 117314 2088 117320 2100
rect 89680 2060 117320 2088
rect 89680 2048 89686 2060
rect 117314 2048 117320 2060
rect 117372 2048 117378 2100
rect 86402 1980 86408 2032
rect 86460 2020 86466 2032
rect 117130 2020 117136 2032
rect 86460 1992 117136 2020
rect 86460 1980 86466 1992
rect 117130 1980 117136 1992
rect 117188 1980 117194 2032
rect 82630 1912 82636 1964
rect 82688 1952 82694 1964
rect 116486 1952 116492 1964
rect 82688 1924 116492 1952
rect 82688 1912 82694 1924
rect 116486 1912 116492 1924
rect 116544 1912 116550 1964
rect 79318 1844 79324 1896
rect 79376 1884 79382 1896
rect 116394 1884 116400 1896
rect 79376 1856 116400 1884
rect 79376 1844 79382 1856
rect 116394 1844 116400 1856
rect 116452 1844 116458 1896
rect 72694 1776 72700 1828
rect 72752 1816 72758 1828
rect 109678 1816 109684 1828
rect 72752 1788 109684 1816
rect 72752 1776 72758 1788
rect 109678 1776 109684 1788
rect 109736 1776 109742 1828
rect 76006 1708 76012 1760
rect 76064 1748 76070 1760
rect 116210 1748 116216 1760
rect 76064 1720 116216 1748
rect 76064 1708 76070 1720
rect 116210 1708 116216 1720
rect 116268 1708 116274 1760
rect 32674 1640 32680 1692
rect 32732 1680 32738 1692
rect 116026 1680 116032 1692
rect 32732 1652 116032 1680
rect 32732 1640 32738 1652
rect 116026 1640 116032 1652
rect 116084 1640 116090 1692
rect 29270 1572 29276 1624
rect 29328 1612 29334 1624
rect 115934 1612 115940 1624
rect 29328 1584 115940 1612
rect 29328 1572 29334 1584
rect 115934 1572 115940 1584
rect 115992 1572 115998 1624
rect 25958 1504 25964 1556
rect 26016 1544 26022 1556
rect 116946 1544 116952 1556
rect 26016 1516 116952 1544
rect 26016 1504 26022 1516
rect 116946 1504 116952 1516
rect 117004 1504 117010 1556
rect 22646 1436 22652 1488
rect 22704 1476 22710 1488
rect 116302 1476 116308 1488
rect 22704 1448 116308 1476
rect 22704 1436 22710 1448
rect 116302 1436 116308 1448
rect 116360 1436 116366 1488
rect 117682 1436 117688 1488
rect 117740 1476 117746 1488
rect 143626 1476 143632 1488
rect 117740 1448 143632 1476
rect 117740 1436 117746 1448
rect 143626 1436 143632 1448
rect 143684 1436 143690 1488
rect 5994 1368 6000 1420
rect 6052 1408 6058 1420
rect 109770 1408 109776 1420
rect 6052 1380 109776 1408
rect 6052 1368 6058 1380
rect 109770 1368 109776 1380
rect 109828 1368 109834 1420
rect 117958 1368 117964 1420
rect 118016 1408 118022 1420
rect 193582 1408 193588 1420
rect 118016 1380 193588 1408
rect 118016 1368 118022 1380
rect 193582 1368 193588 1380
rect 193640 1368 193646 1420
rect 294782 1368 294788 1420
rect 294840 1408 294846 1420
rect 343634 1408 343640 1420
rect 294840 1380 343640 1408
rect 294840 1368 294846 1380
rect 343634 1368 343640 1380
rect 343692 1368 343698 1420
<< via1 >>
rect 83648 160012 83700 160064
rect 167000 160012 167052 160064
rect 170220 160012 170272 160064
rect 198924 160012 198976 160064
rect 211436 160012 211488 160064
rect 280344 160012 280396 160064
rect 281264 160012 281316 160064
rect 330668 160080 330720 160132
rect 327448 160012 327500 160064
rect 334164 160012 334216 160064
rect 334256 160012 334308 160064
rect 335360 160080 335412 160132
rect 335084 160012 335136 160064
rect 374736 160012 374788 160064
rect 378876 160012 378928 160064
rect 398104 160012 398156 160064
rect 404084 160012 404136 160064
rect 427360 160012 427412 160064
rect 25596 159944 25648 159996
rect 109132 159944 109184 159996
rect 117228 159944 117280 159996
rect 191748 159944 191800 159996
rect 198004 159944 198056 159996
rect 270132 159944 270184 159996
rect 271236 159944 271288 159996
rect 272800 159944 272852 159996
rect 275376 159944 275428 159996
rect 329104 159944 329156 159996
rect 329196 159944 329248 159996
rect 370228 159944 370280 159996
rect 374644 159944 374696 159996
rect 388444 159944 388496 159996
rect 389824 159944 389876 159996
rect 413836 159944 413888 159996
rect 70124 159876 70176 159928
rect 148784 159876 148836 159928
rect 148876 159876 148928 159928
rect 56692 159808 56744 159860
rect 136548 159808 136600 159860
rect 136640 159808 136692 159860
rect 63408 159740 63460 159792
rect 146852 159740 146904 159792
rect 18880 159672 18932 159724
rect 107108 159672 107160 159724
rect 109684 159672 109736 159724
rect 137560 159672 137612 159724
rect 139952 159672 140004 159724
rect 147036 159808 147088 159860
rect 150532 159808 150584 159860
rect 147312 159740 147364 159792
rect 148876 159740 148928 159792
rect 152464 159876 152516 159928
rect 160100 159876 160152 159928
rect 160192 159876 160244 159928
rect 188344 159876 188396 159928
rect 191288 159876 191340 159928
rect 264888 159876 264940 159928
rect 268660 159876 268712 159928
rect 324044 159876 324096 159928
rect 328368 159876 328420 159928
rect 369492 159876 369544 159928
rect 372160 159876 372212 159928
rect 396172 159876 396224 159928
rect 403256 159876 403308 159928
rect 416596 159876 416648 159928
rect 450360 159876 450412 159928
rect 457168 159876 457220 159928
rect 458732 159876 458784 159928
rect 465080 159876 465132 159928
rect 478972 159876 479024 159928
rect 484584 159876 484636 159928
rect 150716 159808 150768 159860
rect 174636 159808 174688 159860
rect 49976 159604 50028 159656
rect 143264 159604 143316 159656
rect 143356 159604 143408 159656
rect 146668 159604 146720 159656
rect 32312 159536 32364 159588
rect 126428 159536 126480 159588
rect 126612 159536 126664 159588
rect 146208 159536 146260 159588
rect 146944 159604 146996 159656
rect 149060 159604 149112 159656
rect 153384 159740 153436 159792
rect 153476 159740 153528 159792
rect 180708 159808 180760 159860
rect 184572 159808 184624 159860
rect 259828 159808 259880 159860
rect 261944 159808 261996 159860
rect 318984 159808 319036 159860
rect 320824 159808 320876 159860
rect 357532 159808 357584 159860
rect 177856 159740 177908 159792
rect 253940 159740 253992 159792
rect 255228 159740 255280 159792
rect 313740 159740 313792 159792
rect 314108 159740 314160 159792
rect 357992 159808 358044 159860
rect 376300 159808 376352 159860
rect 406200 159808 406252 159860
rect 467196 159808 467248 159860
rect 473360 159808 473412 159860
rect 357808 159740 357860 159792
rect 365352 159740 365404 159792
rect 365444 159740 365496 159792
rect 395528 159740 395580 159792
rect 396540 159740 396592 159792
rect 413652 159740 413704 159792
rect 424324 159740 424376 159792
rect 442724 159740 442776 159792
rect 471428 159740 471480 159792
rect 477684 159740 477736 159792
rect 149336 159672 149388 159724
rect 164148 159672 164200 159724
rect 167736 159672 167788 159724
rect 245844 159672 245896 159724
rect 248512 159672 248564 159724
rect 160100 159604 160152 159656
rect 161020 159604 161072 159656
rect 240324 159604 240376 159656
rect 241796 159604 241848 159656
rect 302424 159604 302476 159656
rect 308220 159672 308272 159724
rect 347688 159672 347740 159724
rect 347780 159672 347832 159724
rect 378784 159672 378836 159724
rect 379704 159672 379756 159724
rect 405832 159672 405884 159724
rect 409972 159672 410024 159724
rect 417884 159672 417936 159724
rect 420920 159672 420972 159724
rect 440332 159672 440384 159724
rect 308588 159604 308640 159656
rect 309048 159604 309100 159656
rect 354864 159604 354916 159656
rect 355232 159604 355284 159656
rect 362960 159604 363012 159656
rect 369584 159604 369636 159656
rect 401048 159604 401100 159656
rect 414204 159604 414256 159656
rect 435088 159604 435140 159656
rect 459652 159604 459704 159656
rect 466460 159604 466512 159656
rect 468024 159604 468076 159656
rect 476028 159604 476080 159656
rect 157156 159536 157208 159588
rect 157616 159536 157668 159588
rect 239312 159536 239364 159588
rect 250996 159536 251048 159588
rect 310612 159536 310664 159588
rect 315764 159536 315816 159588
rect 358912 159536 358964 159588
rect 362868 159536 362920 159588
rect 394792 159536 394844 159588
rect 399024 159536 399076 159588
rect 408500 159536 408552 159588
rect 410800 159536 410852 159588
rect 432512 159536 432564 159588
rect 448704 159536 448756 159588
rect 456064 159536 456116 159588
rect 460480 159536 460532 159588
rect 466644 159536 466696 159588
rect 470508 159536 470560 159588
rect 476120 159536 476172 159588
rect 479800 159536 479852 159588
rect 485228 159536 485280 159588
rect 43260 159468 43312 159520
rect 137376 159468 137428 159520
rect 137468 159468 137520 159520
rect 146760 159468 146812 159520
rect 36544 159400 36596 159452
rect 135168 159400 135220 159452
rect 136548 159400 136600 159452
rect 144092 159400 144144 159452
rect 144184 159400 144236 159452
rect 225052 159468 225104 159520
rect 231676 159468 231728 159520
rect 295524 159468 295576 159520
rect 295616 159468 295668 159520
rect 339224 159468 339276 159520
rect 339316 159468 339368 159520
rect 349804 159468 349856 159520
rect 147220 159400 147272 159452
rect 150440 159400 150492 159452
rect 150900 159400 150952 159452
rect 234160 159400 234212 159452
rect 234988 159400 235040 159452
rect 298008 159400 298060 159452
rect 301504 159400 301556 159452
rect 347964 159400 348016 159452
rect 348056 159400 348108 159452
rect 354220 159468 354272 159520
rect 358636 159468 358688 159520
rect 392768 159468 392820 159520
rect 407488 159468 407540 159520
rect 429936 159468 429988 159520
rect 449532 159468 449584 159520
rect 455788 159468 455840 159520
rect 457076 159468 457128 159520
rect 464160 159468 464212 159520
rect 468852 159468 468904 159520
rect 474832 159468 474884 159520
rect 477316 159468 477368 159520
rect 483296 159468 483348 159520
rect 518072 159468 518124 159520
rect 522672 159468 522724 159520
rect 351092 159400 351144 159452
rect 355600 159400 355652 159452
rect 356152 159400 356204 159452
rect 390836 159400 390888 159452
rect 427636 159400 427688 159452
rect 445392 159400 445444 159452
rect 451188 159400 451240 159452
rect 456800 159400 456852 159452
rect 6276 159332 6328 159384
rect 122656 159332 122708 159384
rect 123116 159332 123168 159384
rect 146852 159332 146904 159384
rect 146944 159332 146996 159384
rect 223580 159332 223632 159384
rect 224960 159332 225012 159384
rect 290648 159332 290700 159384
rect 294788 159332 294840 159384
rect 76932 159264 76984 159316
rect 152464 159264 152516 159316
rect 163504 159264 163556 159316
rect 196992 159264 197044 159316
rect 201408 159264 201460 159316
rect 212632 159264 212684 159316
rect 214012 159264 214064 159316
rect 281540 159264 281592 159316
rect 282092 159264 282144 159316
rect 327448 159264 327500 159316
rect 327540 159264 327592 159316
rect 330576 159264 330628 159316
rect 330668 159264 330720 159316
rect 333704 159264 333756 159316
rect 335360 159264 335412 159316
rect 338304 159264 338356 159316
rect 93676 159196 93728 159248
rect 86960 159128 87012 159180
rect 169760 159128 169812 159180
rect 180340 159196 180392 159248
rect 183560 159196 183612 159248
rect 187056 159196 187108 159248
rect 216680 159196 216732 159248
rect 218244 159196 218296 159248
rect 285404 159196 285456 159248
rect 287980 159196 288032 159248
rect 338396 159196 338448 159248
rect 338672 159332 338724 159384
rect 339500 159332 339552 159384
rect 339592 159332 339644 159384
rect 342444 159332 342496 159384
rect 346032 159332 346084 159384
rect 382832 159332 382884 159384
rect 392308 159332 392360 159384
rect 403440 159332 403492 159384
rect 417516 159332 417568 159384
rect 437664 159332 437716 159384
rect 447876 159332 447928 159384
rect 338580 159264 338632 159316
rect 374092 159264 374144 159316
rect 378048 159264 378100 159316
rect 388352 159264 388404 159316
rect 388996 159264 389048 159316
rect 403900 159264 403952 159316
rect 453764 159332 453816 159384
rect 459652 159332 459704 159384
rect 469680 159332 469732 159384
rect 477408 159332 477460 159384
rect 478144 159332 478196 159384
rect 483940 159332 483992 159384
rect 518716 159332 518768 159384
rect 523500 159332 523552 159384
rect 456892 159264 456944 159316
rect 457904 159264 457956 159316
rect 464528 159264 464580 159316
rect 342352 159196 342404 159248
rect 342720 159196 342772 159248
rect 343824 159196 343876 159248
rect 349804 159196 349856 159248
rect 377956 159196 378008 159248
rect 385592 159196 385644 159248
rect 399852 159196 399904 159248
rect 461308 159196 461360 159248
rect 468024 159196 468076 159248
rect 176660 159128 176712 159180
rect 181444 159128 181496 159180
rect 100484 159060 100536 159112
rect 183100 159060 183152 159112
rect 193128 159128 193180 159180
rect 193772 159128 193824 159180
rect 220636 159128 220688 159180
rect 224132 159128 224184 159180
rect 288348 159128 288400 159180
rect 288900 159128 288952 159180
rect 339408 159128 339460 159180
rect 341892 159128 341944 159180
rect 378232 159128 378284 159180
rect 395712 159128 395764 159180
rect 405372 159128 405424 159180
rect 462136 159128 462188 159180
rect 467932 159128 467984 159180
rect 183744 159060 183796 159112
rect 203800 159060 203852 159112
rect 203892 159060 203944 159112
rect 210516 159060 210568 159112
rect 210608 159060 210660 159112
rect 215300 159060 215352 159112
rect 220728 159060 220780 159112
rect 278688 159060 278740 159112
rect 278780 159060 278832 159112
rect 279884 159060 279936 159112
rect 280068 159060 280120 159112
rect 282920 159060 282972 159112
rect 283012 159060 283064 159112
rect 284208 159060 284260 159112
rect 284668 159060 284720 159112
rect 285864 159060 285916 159112
rect 302332 159060 302384 159112
rect 349712 159060 349764 159112
rect 351920 159060 351972 159112
rect 385500 159060 385552 159112
rect 386420 159060 386472 159112
rect 387708 159060 387760 159112
rect 412548 159060 412600 159112
rect 413928 159060 413980 159112
rect 462964 159060 463016 159112
rect 469220 159060 469272 159112
rect 472256 159060 472308 159112
rect 479432 159060 479484 159112
rect 107200 158992 107252 159044
rect 73528 158924 73580 158976
rect 107568 158924 107620 158976
rect 119804 158924 119856 158976
rect 126612 158924 126664 158976
rect 96252 158856 96304 158908
rect 120540 158856 120592 158908
rect 120632 158856 120684 158908
rect 121184 158856 121236 158908
rect 124036 158856 124088 158908
rect 181444 158924 181496 158976
rect 183652 158992 183704 159044
rect 185584 158924 185636 158976
rect 102968 158720 103020 158772
rect 125508 158788 125560 158840
rect 127808 158856 127860 158908
rect 130752 158856 130804 158908
rect 195152 158856 195204 158908
rect 197176 158924 197228 158976
rect 200672 158992 200724 159044
rect 227720 158992 227772 159044
rect 230848 158992 230900 159044
rect 295156 158992 295208 159044
rect 200396 158856 200448 158908
rect 203800 158856 203852 158908
rect 204904 158856 204956 158908
rect 210516 158856 210568 158908
rect 213736 158856 213788 158908
rect 106372 158720 106424 158772
rect 127348 158788 127400 158840
rect 130844 158788 130896 158840
rect 133236 158788 133288 158840
rect 126520 158720 126572 158772
rect 137192 158720 137244 158772
rect 137376 158788 137428 158840
rect 147312 158788 147364 158840
rect 147588 158788 147640 158840
rect 149060 158788 149112 158840
rect 149152 158788 149204 158840
rect 156052 158788 156104 158840
rect 156788 158788 156840 158840
rect 194508 158788 194560 158840
rect 194692 158788 194744 158840
rect 203708 158788 203760 158840
rect 208124 158788 208176 158840
rect 211988 158788 212040 158840
rect 217324 158924 217376 158976
rect 220452 158924 220504 158976
rect 238392 158924 238444 158976
rect 242440 158924 242492 158976
rect 299480 158992 299532 159044
rect 307392 158992 307444 159044
rect 353208 158992 353260 159044
rect 355600 158992 355652 159044
rect 382556 158992 382608 159044
rect 383108 158992 383160 159044
rect 411444 158992 411496 159044
rect 455420 158992 455472 159044
rect 463332 158992 463384 159044
rect 473912 158992 473964 159044
rect 480260 158992 480312 159044
rect 480628 158992 480680 159044
rect 485872 158992 485924 159044
rect 507124 158992 507176 159044
rect 508412 158992 508464 159044
rect 214748 158856 214800 158908
rect 305368 158924 305420 158976
rect 310704 158924 310756 158976
rect 313188 158924 313240 158976
rect 314936 158924 314988 158976
rect 357440 158924 357492 158976
rect 357532 158924 357584 158976
rect 363512 158924 363564 158976
rect 158720 158720 158772 158772
rect 171140 158720 171192 158772
rect 172612 158720 172664 158772
rect 173624 158720 173676 158772
rect 197360 158720 197412 158772
rect 207296 158720 207348 158772
rect 214564 158720 214616 158772
rect 214840 158788 214892 158840
rect 221464 158788 221516 158840
rect 221556 158788 221608 158840
rect 224776 158788 224828 158840
rect 231308 158788 231360 158840
rect 237564 158788 237616 158840
rect 244280 158788 244332 158840
rect 298100 158856 298152 158908
rect 300308 158856 300360 158908
rect 305644 158856 305696 158908
rect 307300 158856 307352 158908
rect 312452 158856 312504 158908
rect 313464 158856 313516 158908
rect 365168 158924 365220 158976
rect 365352 158924 365404 158976
rect 378692 158924 378744 158976
rect 386236 158924 386288 158976
rect 391480 158924 391532 158976
rect 394332 158924 394384 158976
rect 409144 158924 409196 158976
rect 410892 158924 410944 158976
rect 416688 158924 416740 158976
rect 419540 158924 419592 158976
rect 420092 158924 420144 158976
rect 423588 158924 423640 158976
rect 454592 158924 454644 158976
rect 461860 158924 461912 158976
rect 466368 158924 466420 158976
rect 472532 158924 472584 158976
rect 475568 158924 475620 158976
rect 482008 158924 482060 158976
rect 261116 158788 261168 158840
rect 317144 158788 317196 158840
rect 317420 158788 317472 158840
rect 318432 158788 318484 158840
rect 319168 158788 319220 158840
rect 321560 158788 321612 158840
rect 322480 158788 322532 158840
rect 222108 158720 222160 158772
rect 240876 158720 240928 158772
rect 243360 158720 243412 158772
rect 254400 158720 254452 158772
rect 255412 158720 255464 158772
rect 258540 158720 258592 158772
rect 261024 158720 261076 158772
rect 264428 158720 264480 158772
rect 267648 158720 267700 158772
rect 267832 158720 267884 158772
rect 320272 158720 320324 158772
rect 321652 158720 321704 158772
rect 355232 158788 355284 158840
rect 330576 158720 330628 158772
rect 361304 158788 361356 158840
rect 384764 158856 384816 158908
rect 389640 158856 389692 158908
rect 446128 158856 446180 158908
rect 453948 158856 454000 158908
rect 456248 158856 456300 158908
rect 462964 158856 463016 158908
rect 463792 158856 463844 158908
rect 471244 158856 471296 158908
rect 474740 158856 474792 158908
rect 481364 158856 481416 158908
rect 481456 158856 481508 158908
rect 486424 158856 486476 158908
rect 508412 158856 508464 158908
rect 510068 158856 510120 158908
rect 367192 158720 367244 158772
rect 367928 158720 367980 158772
rect 378692 158720 378744 158772
rect 384948 158788 385000 158840
rect 404912 158788 404964 158840
rect 405648 158788 405700 158840
rect 452016 158788 452068 158840
rect 458180 158788 458232 158840
rect 464620 158788 464672 158840
rect 471612 158788 471664 158840
rect 476396 158788 476448 158840
rect 481640 158788 481692 158840
rect 499948 158788 500000 158840
rect 500592 158788 500644 158840
rect 506296 158788 506348 158840
rect 507584 158788 507636 158840
rect 385316 158720 385368 158772
rect 388076 158720 388128 158772
rect 390376 158720 390428 158772
rect 405740 158720 405792 158772
rect 409144 158720 409196 158772
rect 413376 158720 413428 158772
rect 419632 158720 419684 158772
rect 435180 158720 435232 158772
rect 435824 158720 435876 158772
rect 452844 158720 452896 158772
rect 459560 158720 459612 158772
rect 465540 158720 465592 158772
rect 472440 158720 472492 158772
rect 473084 158720 473136 158772
rect 478972 158720 479024 158772
rect 482284 158720 482336 158772
rect 487252 158720 487304 158772
rect 504456 158720 504508 158772
rect 505008 158720 505060 158772
rect 505836 158720 505888 158772
rect 506480 158720 506532 158772
rect 509700 158720 509752 158772
rect 511724 158720 511776 158772
rect 514944 158720 514996 158772
rect 518532 158720 518584 158772
rect 81072 158652 81124 158704
rect 180800 158652 180852 158704
rect 180892 158652 180944 158704
rect 181904 158652 181956 158704
rect 181996 158652 182048 158704
rect 256792 158652 256844 158704
rect 67640 158584 67692 158636
rect 170312 158584 170364 158636
rect 171968 158584 172020 158636
rect 250076 158584 250128 158636
rect 71044 158516 71096 158568
rect 172704 158516 172756 158568
rect 178684 158516 178736 158568
rect 255320 158516 255372 158568
rect 74356 158448 74408 158500
rect 175188 158448 175240 158500
rect 175280 158448 175332 158500
rect 252560 158448 252612 158500
rect 64236 158380 64288 158432
rect 167552 158380 167604 158432
rect 168564 158380 168616 158432
rect 247592 158380 247644 158432
rect 60924 158312 60976 158364
rect 164332 158312 164384 158364
rect 165252 158312 165304 158364
rect 245016 158312 245068 158364
rect 54208 158244 54260 158296
rect 160284 158244 160336 158296
rect 161848 158244 161900 158296
rect 242072 158244 242124 158296
rect 50804 158176 50856 158228
rect 157708 158176 157760 158228
rect 158444 158176 158496 158228
rect 238852 158176 238904 158228
rect 256884 158176 256936 158228
rect 315028 158176 315080 158228
rect 47492 158108 47544 158160
rect 155040 158108 155092 158160
rect 155132 158108 155184 158160
rect 237380 158108 237432 158160
rect 246764 158108 246816 158160
rect 306932 158108 306984 158160
rect 37372 158040 37424 158092
rect 146392 158040 146444 158092
rect 148416 158040 148468 158092
rect 231860 158040 231912 158092
rect 233332 158040 233384 158092
rect 297088 158040 297140 158092
rect 300676 158040 300728 158092
rect 348424 158040 348476 158092
rect 388 157972 440 158024
rect 118884 157972 118936 158024
rect 131580 157972 131632 158024
rect 218244 157972 218296 158024
rect 240048 157972 240100 158024
rect 302240 157972 302292 158024
rect 77760 157904 77812 157956
rect 84476 157836 84528 157888
rect 175924 157836 175976 157888
rect 176200 157904 176252 157956
rect 182272 157904 182324 157956
rect 185400 157904 185452 157956
rect 259460 157904 259512 157956
rect 178040 157836 178092 157888
rect 181536 157836 181588 157888
rect 188528 157836 188580 157888
rect 188804 157836 188856 157888
rect 263048 157836 263100 157888
rect 87788 157768 87840 157820
rect 181628 157768 181680 157820
rect 181812 157768 181864 157820
rect 190644 157768 190696 157820
rect 195520 157768 195572 157820
rect 267740 157768 267792 157820
rect 91192 157700 91244 157752
rect 181260 157700 181312 157752
rect 181904 157700 181956 157752
rect 94596 157632 94648 157684
rect 181536 157632 181588 157684
rect 181720 157632 181772 157684
rect 185400 157632 185452 157684
rect 190460 157700 190512 157752
rect 263784 157700 263836 157752
rect 236092 157632 236144 157684
rect 97908 157564 97960 157616
rect 193220 157564 193272 157616
rect 197360 157564 197412 157616
rect 251456 157564 251508 157616
rect 111340 157496 111392 157548
rect 203432 157496 203484 157548
rect 204904 157496 204956 157548
rect 258080 157496 258132 157548
rect 114744 157428 114796 157480
rect 206560 157428 206612 157480
rect 141700 157360 141752 157412
rect 227076 157360 227128 157412
rect 55864 157292 55916 157344
rect 161572 157292 161624 157344
rect 52460 157224 52512 157276
rect 158996 157224 159048 157276
rect 160100 157224 160152 157276
rect 204904 157292 204956 157344
rect 204996 157292 205048 157344
rect 273260 157292 273312 157344
rect 192116 157224 192168 157276
rect 265164 157224 265216 157276
rect 290556 157224 290608 157276
rect 339960 157224 340012 157276
rect 45744 157156 45796 157208
rect 153752 157156 153804 157208
rect 166908 157156 166960 157208
rect 246304 157156 246356 157208
rect 280436 157156 280488 157208
rect 332692 157156 332744 157208
rect 39028 157088 39080 157140
rect 143724 157088 143776 157140
rect 35716 157020 35768 157072
rect 145472 157088 145524 157140
rect 151728 157088 151780 157140
rect 234804 157088 234856 157140
rect 273720 157088 273772 157140
rect 327908 157088 327960 157140
rect 145288 157020 145340 157072
rect 229652 157020 229704 157072
rect 277124 157020 277176 157072
rect 330484 157020 330536 157072
rect 24768 156952 24820 157004
rect 137192 156952 137244 157004
rect 139124 156952 139176 157004
rect 225144 156952 225196 157004
rect 270316 156952 270368 157004
rect 325332 156952 325384 157004
rect 18052 156884 18104 156936
rect 132500 156884 132552 156936
rect 134892 156884 134944 156936
rect 213828 156884 213880 156936
rect 213920 156884 213972 156936
rect 223120 156884 223172 156936
rect 226616 156884 226668 156936
rect 291936 156884 291988 156936
rect 21364 156816 21416 156868
rect 135260 156816 135312 156868
rect 135812 156816 135864 156868
rect 222568 156816 222620 156868
rect 230020 156816 230072 156868
rect 294052 156816 294104 156868
rect 297272 156816 297324 156868
rect 345848 156816 345900 156868
rect 11244 156748 11296 156800
rect 127532 156748 127584 156800
rect 128176 156748 128228 156800
rect 216772 156748 216824 156800
rect 219900 156748 219952 156800
rect 285680 156748 285732 156800
rect 287152 156748 287204 156800
rect 338120 156748 338172 156800
rect 14648 156680 14700 156732
rect 130108 156680 130160 156732
rect 132408 156680 132460 156732
rect 219992 156680 220044 156732
rect 223212 156680 223264 156732
rect 289360 156680 289412 156732
rect 293868 156680 293920 156732
rect 343272 156680 343324 156732
rect 344376 156680 344428 156732
rect 381820 156680 381872 156732
rect 2044 156612 2096 156664
rect 120448 156612 120500 156664
rect 121460 156612 121512 156664
rect 201316 156612 201368 156664
rect 143724 156544 143776 156596
rect 147680 156544 147732 156596
rect 158720 156544 158772 156596
rect 219900 156612 219952 156664
rect 220084 156612 220136 156664
rect 281632 156612 281684 156664
rect 283840 156612 283892 156664
rect 335544 156612 335596 156664
rect 337660 156612 337712 156664
rect 375564 156612 375616 156664
rect 72700 156476 72752 156528
rect 174452 156476 174504 156528
rect 174636 156476 174688 156528
rect 79416 156408 79468 156460
rect 179604 156408 179656 156460
rect 198832 156476 198884 156528
rect 270500 156544 270552 156596
rect 204904 156476 204956 156528
rect 213920 156476 213972 156528
rect 214564 156476 214616 156528
rect 273904 156476 273956 156528
rect 92848 156340 92900 156392
rect 189816 156340 189868 156392
rect 101312 156272 101364 156324
rect 196256 156272 196308 156324
rect 201316 156408 201368 156460
rect 211620 156408 211672 156460
rect 202236 156340 202288 156392
rect 204996 156340 205048 156392
rect 209780 156340 209832 156392
rect 279056 156408 279108 156460
rect 216496 156340 216548 156392
rect 283104 156340 283156 156392
rect 230940 156272 230992 156324
rect 108028 156204 108080 156256
rect 200304 156204 200356 156256
rect 203064 156204 203116 156256
rect 214564 156204 214616 156256
rect 222108 156204 222160 156256
rect 269212 156204 269264 156256
rect 118148 156136 118200 156188
rect 209136 156136 209188 156188
rect 213184 156136 213236 156188
rect 220084 156136 220136 156188
rect 220636 156136 220688 156188
rect 266912 156136 266964 156188
rect 124864 156068 124916 156120
rect 213920 156068 213972 156120
rect 219900 156068 219952 156120
rect 220544 156068 220596 156120
rect 227720 156068 227772 156120
rect 272064 156068 272116 156120
rect 138296 156000 138348 156052
rect 224500 156000 224552 156052
rect 59268 155932 59320 155984
rect 164148 155932 164200 155984
rect 164240 155932 164292 155984
rect 228364 155932 228416 155984
rect 60096 155864 60148 155916
rect 85488 155864 85540 155916
rect 88708 155864 88760 155916
rect 186780 155864 186832 155916
rect 189632 155864 189684 155916
rect 263692 155864 263744 155916
rect 303160 155864 303212 155916
rect 350356 155864 350408 155916
rect 12164 155796 12216 155848
rect 109684 155796 109736 155848
rect 112260 155796 112312 155848
rect 204628 155796 204680 155848
rect 206468 155796 206520 155848
rect 276020 155796 276072 155848
rect 293040 155796 293092 155848
rect 342628 155796 342680 155848
rect 53380 155728 53432 155780
rect 76748 155728 76800 155780
rect 81900 155728 81952 155780
rect 181444 155728 181496 155780
rect 186228 155728 186280 155780
rect 260840 155728 260892 155780
rect 296444 155728 296496 155780
rect 345204 155728 345256 155780
rect 33140 155660 33192 155712
rect 60004 155660 60056 155712
rect 71872 155660 71924 155712
rect 173072 155660 173124 155712
rect 176292 155660 176344 155712
rect 46572 155592 46624 155644
rect 75092 155592 75144 155644
rect 75184 155592 75236 155644
rect 176384 155592 176436 155644
rect 177120 155660 177172 155712
rect 254032 155660 254084 155712
rect 289728 155660 289780 155712
rect 339592 155660 339644 155712
rect 253388 155592 253440 155644
rect 267004 155592 267056 155644
rect 322112 155592 322164 155644
rect 39856 155524 39908 155576
rect 71780 155524 71832 155576
rect 78588 155524 78640 155576
rect 178960 155524 179012 155576
rect 179512 155524 179564 155576
rect 255872 155524 255924 155576
rect 263600 155524 263652 155576
rect 320180 155524 320232 155576
rect 340972 155524 341024 155576
rect 378140 155524 378192 155576
rect 28908 155456 28960 155508
rect 56232 155456 56284 155508
rect 62580 155456 62632 155508
rect 165620 155456 165672 155508
rect 169392 155456 169444 155508
rect 247132 155456 247184 155508
rect 260288 155456 260340 155508
rect 317604 155456 317656 155508
rect 333428 155456 333480 155508
rect 373448 155456 373500 155508
rect 7932 155388 7984 155440
rect 122012 155388 122064 155440
rect 4528 155320 4580 155372
rect 121920 155320 121972 155372
rect 8760 155252 8812 155304
rect 125600 155388 125652 155440
rect 134064 155388 134116 155440
rect 137468 155388 137520 155440
rect 142528 155388 142580 155440
rect 227720 155388 227772 155440
rect 250168 155388 250220 155440
rect 309876 155388 309928 155440
rect 330116 155388 330168 155440
rect 369860 155388 369912 155440
rect 122288 155320 122340 155372
rect 211252 155320 211304 155372
rect 213828 155320 213880 155372
rect 125692 155252 125744 155304
rect 214840 155252 214892 155304
rect 216680 155320 216732 155372
rect 261392 155320 261444 155372
rect 263600 155320 263652 155372
rect 263784 155320 263836 155372
rect 316592 155320 316644 155372
rect 360660 155320 360712 155372
rect 221924 155252 221976 155304
rect 243452 155252 243504 155304
rect 304724 155252 304776 155304
rect 309968 155252 310020 155304
rect 354680 155252 354732 155304
rect 373816 155252 373868 155304
rect 403164 155252 403216 155304
rect 5356 155184 5408 155236
rect 123024 155184 123076 155236
rect 129004 155184 129056 155236
rect 217416 155184 217468 155236
rect 236736 155184 236788 155236
rect 299664 155184 299716 155236
rect 299756 155184 299808 155236
rect 347780 155184 347832 155236
rect 367100 155184 367152 155236
rect 399116 155184 399168 155236
rect 401600 155184 401652 155236
rect 425520 155184 425572 155236
rect 86132 155116 86184 155168
rect 183560 155116 183612 155168
rect 186688 155116 186740 155168
rect 95424 155048 95476 155100
rect 186320 155048 186372 155100
rect 186504 155048 186556 155100
rect 191748 155048 191800 155100
rect 192944 155116 192996 155168
rect 266084 155116 266136 155168
rect 306564 155116 306616 155168
rect 352932 155116 352984 155168
rect 194968 155048 195020 155100
rect 196348 155048 196400 155100
rect 268844 155048 268896 155100
rect 98736 154980 98788 155032
rect 186228 154980 186280 155032
rect 186596 154980 186648 155032
rect 194324 154980 194376 155032
rect 199660 154980 199712 155032
rect 271420 154980 271472 155032
rect 80244 154912 80296 154964
rect 86868 154912 86920 154964
rect 99564 154912 99616 154964
rect 186320 154912 186372 154964
rect 188344 154912 188396 154964
rect 240692 154912 240744 154964
rect 253572 154912 253624 154964
rect 312452 154912 312504 154964
rect 107108 154844 107160 154896
rect 133328 154844 133380 154896
rect 145840 154844 145892 154896
rect 229192 154844 229244 154896
rect 231308 154844 231360 154896
rect 277124 154844 277176 154896
rect 110512 154776 110564 154828
rect 128360 154776 128412 154828
rect 149244 154776 149296 154828
rect 232872 154776 232924 154828
rect 122012 154708 122064 154760
rect 124956 154708 125008 154760
rect 155960 154708 156012 154760
rect 238024 154708 238076 154760
rect 118976 154640 119028 154692
rect 124404 154640 124456 154692
rect 146208 154640 146260 154692
rect 121920 154572 121972 154624
rect 122380 154572 122432 154624
rect 44916 154504 44968 154556
rect 146484 154504 146536 154556
rect 41604 154436 41656 154488
rect 150624 154504 150676 154556
rect 162676 154640 162728 154692
rect 243084 154640 243136 154692
rect 159364 154572 159416 154624
rect 240140 154572 240192 154624
rect 156788 154504 156840 154556
rect 157340 154504 157392 154556
rect 225788 154504 225840 154556
rect 232504 154504 232556 154556
rect 296444 154504 296496 154556
rect 357348 154504 357400 154556
rect 391480 154504 391532 154556
rect 34796 154368 34848 154420
rect 145380 154368 145432 154420
rect 38476 154300 38528 154352
rect 145104 154300 145156 154352
rect 30656 154232 30708 154284
rect 137100 154232 137152 154284
rect 185124 154436 185176 154488
rect 191288 154436 191340 154488
rect 200120 154436 200172 154488
rect 225880 154436 225932 154488
rect 291292 154436 291344 154488
rect 353668 154436 353720 154488
rect 388904 154436 388956 154488
rect 400772 154436 400824 154488
rect 424876 154436 424928 154488
rect 23940 154164 23992 154216
rect 137008 154164 137060 154216
rect 13820 154096 13872 154148
rect 10416 154028 10468 154080
rect 120632 154028 120684 154080
rect 121552 154096 121604 154148
rect 188436 154368 188488 154420
rect 191472 154368 191524 154420
rect 202696 154368 202748 154420
rect 208952 154368 209004 154420
rect 278412 154368 278464 154420
rect 279976 154368 280028 154420
rect 332416 154368 332468 154420
rect 350264 154368 350316 154420
rect 386328 154368 386380 154420
rect 398196 154368 398248 154420
rect 423036 154368 423088 154420
rect 146944 154300 146996 154352
rect 191288 154300 191340 154352
rect 191380 154300 191432 154352
rect 202052 154300 202104 154352
rect 205548 154300 205600 154352
rect 275836 154300 275888 154352
rect 276204 154300 276256 154352
rect 329840 154300 329892 154352
rect 346860 154300 346912 154352
rect 383752 154300 383804 154352
rect 390652 154300 390704 154352
rect 417148 154300 417200 154352
rect 129464 154028 129516 154080
rect 129556 154028 129608 154080
rect 7104 153960 7156 154012
rect 118608 153960 118660 154012
rect 118700 153960 118752 154012
rect 1216 153892 1268 153944
rect 119804 153892 119856 153944
rect 124312 153960 124364 154012
rect 124404 153960 124456 154012
rect 120724 153892 120776 153944
rect 126888 153892 126940 153944
rect 127808 153960 127860 154012
rect 146852 154096 146904 154148
rect 137560 154028 137612 154080
rect 185216 154232 185268 154284
rect 185308 154232 185360 154284
rect 258540 154232 258592 154284
rect 266176 154232 266228 154284
rect 322020 154232 322072 154284
rect 343548 154232 343600 154284
rect 381176 154232 381228 154284
rect 393964 154232 394016 154284
rect 419724 154232 419776 154284
rect 147128 154164 147180 154216
rect 156604 154164 156656 154216
rect 156696 154164 156748 154216
rect 163504 154164 163556 154216
rect 165068 154164 165120 154216
rect 168656 154164 168708 154216
rect 172796 154164 172848 154216
rect 250812 154164 250864 154216
rect 252652 154164 252704 154216
rect 311716 154164 311768 154216
rect 326712 154164 326764 154216
rect 368296 154164 368348 154216
rect 387616 154164 387668 154216
rect 414572 154164 414624 154216
rect 147036 154096 147088 154148
rect 153200 154096 153252 154148
rect 153384 154096 153436 154148
rect 166264 154096 166316 154148
rect 166356 154096 166408 154148
rect 245660 154096 245712 154148
rect 245936 154096 245988 154148
rect 306656 154096 306708 154148
rect 323308 154096 323360 154148
rect 365720 154096 365772 154148
rect 383936 154096 383988 154148
rect 411996 154096 412048 154148
rect 152648 154028 152700 154080
rect 235448 154028 235500 154080
rect 242624 154028 242676 154080
rect 304080 154028 304132 154080
rect 319996 154028 320048 154080
rect 363236 154028 363288 154080
rect 370412 154028 370464 154080
rect 401692 154028 401744 154080
rect 137652 153960 137704 154012
rect 142344 153960 142396 154012
rect 145104 153960 145156 154012
rect 148140 153960 148192 154012
rect 150348 153960 150400 154012
rect 233516 153960 233568 154012
rect 235908 153960 235960 154012
rect 299020 153960 299072 154012
rect 313280 153960 313332 154012
rect 357900 153960 357952 154012
rect 363696 153960 363748 154012
rect 396540 153960 396592 154012
rect 397368 153960 397420 154012
rect 422300 153960 422352 154012
rect 209780 153892 209832 153944
rect 215668 153892 215720 153944
rect 283656 153892 283708 153944
rect 284208 153892 284260 153944
rect 334900 153892 334952 153944
rect 336832 153892 336884 153944
rect 3976 153824 4028 153876
rect 113824 153824 113876 153876
rect 115572 153824 115624 153876
rect 118516 153824 118568 153876
rect 118608 153824 118660 153876
rect 118700 153824 118752 153876
rect 125508 153824 125560 153876
rect 129556 153824 129608 153876
rect 129924 153824 129976 153876
rect 218060 153824 218112 153876
rect 219348 153824 219400 153876
rect 286140 153824 286192 153876
rect 286324 153824 286376 153876
rect 337476 153824 337528 153876
rect 340144 153892 340196 153944
rect 378600 153892 378652 153944
rect 380808 153892 380860 153944
rect 409420 153892 409472 153944
rect 376024 153824 376076 153876
rect 377220 153824 377272 153876
rect 406844 153824 406896 153876
rect 48320 153756 48372 153808
rect 155776 153756 155828 153808
rect 156604 153756 156656 153808
rect 212908 153756 212960 153808
rect 222384 153756 222436 153808
rect 288716 153756 288768 153808
rect 360384 153756 360436 153808
rect 394056 153756 394108 153808
rect 58348 153688 58400 153740
rect 156696 153688 156748 153740
rect 156788 153688 156840 153740
rect 210424 153688 210476 153740
rect 229100 153688 229152 153740
rect 293868 153688 293920 153740
rect 65156 153620 65208 153672
rect 165068 153620 165120 153672
rect 166264 153620 166316 153672
rect 215484 153620 215536 153672
rect 239220 153620 239272 153672
rect 301596 153620 301648 153672
rect 82820 153552 82872 153604
rect 182088 153552 182140 153604
rect 182916 153552 182968 153604
rect 185032 153552 185084 153604
rect 185124 153552 185176 153604
rect 188344 153552 188396 153604
rect 188436 153552 188488 153604
rect 197544 153552 197596 153604
rect 198924 153552 198976 153604
rect 248880 153552 248932 153604
rect 249708 153552 249760 153604
rect 309232 153552 309284 153604
rect 102140 153484 102192 153536
rect 196900 153484 196952 153536
rect 196992 153484 197044 153536
rect 199384 153484 199436 153536
rect 108856 153416 108908 153468
rect 191380 153416 191432 153468
rect 194508 153416 194560 153468
rect 200396 153484 200448 153536
rect 256516 153484 256568 153536
rect 238668 153416 238720 153468
rect 105452 153348 105504 153400
rect 199476 153348 199528 153400
rect 199568 153348 199620 153400
rect 243728 153348 243780 153400
rect 256056 153348 256108 153400
rect 314384 153484 314436 153536
rect 262772 153416 262824 153468
rect 319536 153416 319588 153468
rect 259552 153348 259604 153400
rect 316960 153348 317012 153400
rect 113824 153280 113876 153332
rect 118424 153280 118476 153332
rect 120724 153280 120776 153332
rect 207204 153280 207256 153332
rect 272892 153280 272944 153332
rect 327264 153280 327316 153332
rect 119436 153212 119488 153264
rect 207848 153212 207900 153264
rect 269488 153212 269540 153264
rect 324688 153212 324740 153264
rect 118516 153144 118568 153196
rect 120724 153144 120776 153196
rect 123484 153144 123536 153196
rect 205916 153144 205968 153196
rect 225052 153144 225104 153196
rect 229008 153144 229060 153196
rect 234436 153144 234488 153196
rect 297732 153144 297784 153196
rect 300308 153144 300360 153196
rect 342260 153144 342312 153196
rect 342352 153144 342404 153196
rect 343916 153144 343968 153196
rect 345296 153144 345348 153196
rect 345756 153144 345808 153196
rect 349436 153144 349488 153196
rect 385592 153144 385644 153196
rect 390376 153144 390428 153196
rect 415216 153144 415268 153196
rect 415860 153144 415912 153196
rect 433064 153212 433116 153264
rect 103796 153076 103848 153128
rect 198188 153076 198240 153128
rect 215300 153076 215352 153128
rect 279700 153076 279752 153128
rect 279884 153076 279936 153128
rect 331772 153076 331824 153128
rect 332600 153076 332652 153128
rect 372804 153076 372856 153128
rect 372988 153076 373040 153128
rect 403624 153076 403676 153128
rect 408500 153076 408552 153128
rect 415124 153076 415176 153128
rect 415308 153076 415360 153128
rect 435732 153144 435784 153196
rect 435824 153144 435876 153196
rect 86868 153008 86920 153060
rect 180248 153008 180300 153060
rect 181168 153008 181220 153060
rect 257252 153008 257304 153060
rect 257712 153008 257764 153060
rect 315672 153008 315724 153060
rect 317144 153008 317196 153060
rect 318248 153008 318300 153060
rect 318432 153008 318484 153060
rect 361304 153008 361356 153060
rect 367192 153008 367244 153060
rect 368940 153008 368992 153060
rect 369032 153008 369084 153060
rect 397184 153008 397236 153060
rect 398104 153008 398156 153060
rect 408132 153008 408184 153060
rect 411628 153008 411680 153060
rect 433156 153076 433208 153128
rect 433248 153076 433300 153128
rect 436376 153076 436428 153128
rect 437296 153144 437348 153196
rect 452476 153144 452528 153196
rect 453948 153144 454000 153196
rect 459468 153144 459520 153196
rect 461860 153144 461912 153196
rect 465908 153144 465960 153196
rect 466460 153144 466512 153196
rect 469772 153144 469824 153196
rect 471244 153144 471296 153196
rect 472992 153144 473044 153196
rect 474832 153144 474884 153196
rect 476856 153144 476908 153196
rect 485688 153144 485740 153196
rect 489644 153144 489696 153196
rect 490748 153144 490800 153196
rect 493508 153144 493560 153196
rect 494060 153144 494112 153196
rect 496084 153144 496136 153196
rect 496636 153144 496688 153196
rect 498016 153144 498068 153196
rect 498292 153144 498344 153196
rect 499304 153144 499356 153196
rect 500960 153144 501012 153196
rect 501880 153144 501932 153196
rect 511632 153144 511684 153196
rect 513748 153144 513800 153196
rect 514208 153144 514260 153196
rect 517428 153144 517480 153196
rect 438492 153076 438544 153128
rect 438584 153076 438636 153128
rect 453764 153076 453816 153128
rect 456892 153076 456944 153128
rect 460756 153076 460808 153128
rect 462964 153076 463016 153128
rect 467196 153076 467248 153128
rect 471612 153076 471664 153128
rect 473636 153076 473688 153128
rect 476120 153076 476172 153128
rect 478144 153076 478196 153128
rect 484860 153076 484912 153128
rect 489000 153076 489052 153128
rect 489920 153076 489972 153128
rect 492864 153076 492916 153128
rect 493232 153076 493284 153128
rect 495440 153076 495492 153128
rect 495808 153076 495860 153128
rect 497372 153076 497424 153128
rect 497464 153076 497516 153128
rect 498660 153076 498712 153128
rect 510988 153076 511040 153128
rect 513472 153076 513524 153128
rect 513564 153076 513616 153128
rect 516140 153076 516192 153128
rect 432696 153008 432748 153060
rect 449256 153008 449308 153060
rect 463332 153008 463384 153060
rect 466552 153008 466604 153060
rect 466644 153008 466696 153060
rect 470416 153008 470468 153060
rect 472440 153008 472492 153060
rect 474280 153008 474332 153060
rect 484032 153008 484084 153060
rect 488356 153008 488408 153060
rect 492404 153008 492456 153060
rect 494796 153008 494848 153060
rect 495256 153008 495308 153060
rect 496636 153008 496688 153060
rect 512276 153008 512328 153060
rect 514852 153008 514904 153060
rect 97080 152940 97132 152992
rect 193036 152940 193088 152992
rect 203708 152940 203760 152992
rect 267556 152940 267608 152992
rect 267648 152940 267700 152992
rect 320916 152940 320968 152992
rect 325884 152940 325936 152992
rect 367652 152940 367704 152992
rect 368756 152940 368808 152992
rect 400404 152940 400456 152992
rect 407028 152940 407080 152992
rect 429200 152940 429252 152992
rect 429292 152940 429344 152992
rect 446680 152940 446732 152992
rect 459560 152940 459612 152992
rect 464620 152940 464672 152992
rect 465080 152940 465132 152992
rect 469128 152940 469180 152992
rect 472532 152940 472584 152992
rect 474924 152940 474976 152992
rect 483204 152940 483256 152992
rect 487804 152940 487856 152992
rect 491576 152940 491628 152992
rect 494152 152940 494204 152992
rect 512920 152940 512972 152992
rect 515956 152940 516008 152992
rect 90364 152872 90416 152924
rect 187884 152872 187936 152924
rect 187976 152872 188028 152924
rect 262404 152872 262456 152924
rect 270868 152872 270920 152924
rect 321468 152872 321520 152924
rect 321560 152872 321612 152924
rect 323492 152872 323544 152924
rect 324228 152872 324280 152924
rect 366364 152872 366416 152924
rect 366456 152872 366508 152924
rect 398472 152872 398524 152924
rect 402428 152872 402480 152924
rect 426164 152872 426216 152924
rect 426256 152872 426308 152924
rect 427176 152872 427228 152924
rect 430488 152872 430540 152924
rect 447324 152872 447376 152924
rect 464160 152872 464212 152924
rect 467840 152872 467892 152924
rect 473360 152872 473412 152924
rect 475568 152872 475620 152924
rect 66812 152804 66864 152856
rect 169944 152804 169996 152856
rect 174544 152804 174596 152856
rect 252100 152804 252152 152856
rect 252192 152804 252244 152856
rect 311164 152804 311216 152856
rect 318708 152804 318760 152856
rect 361948 152804 362000 152856
rect 362040 152804 362092 152856
rect 395436 152804 395488 152856
rect 395528 152804 395580 152856
rect 397828 152804 397880 152856
rect 400128 152804 400180 152856
rect 424232 152804 424284 152856
rect 425152 152804 425204 152856
rect 443460 152804 443512 152856
rect 444472 152804 444524 152856
rect 458272 152804 458324 152856
rect 464528 152804 464580 152856
rect 468392 152804 468444 152856
rect 510344 152804 510396 152856
rect 512000 152804 512052 152856
rect 26424 152736 26476 152788
rect 139124 152736 139176 152788
rect 22192 152668 22244 152720
rect 135904 152668 135956 152720
rect 137468 152668 137520 152720
rect 143540 152736 143592 152788
rect 139400 152668 139452 152720
rect 141700 152668 141752 152720
rect 141792 152668 141844 152720
rect 151912 152736 151964 152788
rect 154304 152736 154356 152788
rect 236736 152736 236788 152788
rect 240324 152736 240376 152788
rect 241888 152736 241940 152788
rect 247684 152736 247736 152788
rect 307944 152736 307996 152788
rect 311808 152736 311860 152788
rect 356796 152736 356848 152788
rect 357440 152736 357492 152788
rect 359372 152736 359424 152788
rect 359556 152736 359608 152788
rect 393412 152736 393464 152788
rect 394884 152736 394936 152788
rect 420368 152736 420420 152788
rect 421748 152736 421800 152788
rect 433340 152736 433392 152788
rect 433432 152736 433484 152788
rect 438952 152736 439004 152788
rect 442816 152736 442868 152788
rect 456984 152736 457036 152788
rect 143816 152668 143868 152720
rect 221280 152668 221332 152720
rect 224776 152668 224828 152720
rect 288072 152668 288124 152720
rect 288348 152668 288400 152720
rect 290004 152668 290056 152720
rect 291384 152668 291436 152720
rect 341340 152668 341392 152720
rect 342444 152668 342496 152720
rect 344560 152668 344612 152720
rect 15476 152600 15528 152652
rect 130752 152600 130804 152652
rect 130844 152600 130896 152652
rect 216128 152600 216180 152652
rect 220452 152600 220504 152652
rect 284852 152600 284904 152652
rect 19708 152532 19760 152584
rect 133972 152532 134024 152584
rect 135168 152532 135220 152584
rect 138572 152532 138624 152584
rect 140780 152532 140832 152584
rect 226432 152532 226484 152584
rect 228272 152532 228324 152584
rect 293224 152600 293276 152652
rect 336188 152600 336240 152652
rect 336280 152600 336332 152652
rect 345388 152600 345440 152652
rect 2872 152464 2924 152516
rect 121092 152464 121144 152516
rect 121184 152464 121236 152516
rect 211068 152464 211120 152516
rect 211988 152464 212040 152516
rect 277768 152464 277820 152516
rect 285864 152464 285916 152516
rect 299388 152532 299440 152584
rect 347136 152668 347188 152720
rect 349068 152668 349120 152720
rect 352380 152668 352432 152720
rect 352472 152668 352524 152720
rect 382464 152668 382516 152720
rect 382556 152668 382608 152720
rect 386972 152668 387024 152720
rect 387708 152668 387760 152720
rect 413928 152668 413980 152720
rect 414020 152668 414072 152720
rect 427084 152668 427136 152720
rect 427176 152668 427228 152720
rect 431592 152668 431644 152720
rect 434628 152668 434680 152720
rect 450544 152668 450596 152720
rect 458180 152668 458232 152720
rect 463976 152668 464028 152720
rect 345572 152600 345624 152652
rect 375380 152600 375432 152652
rect 375472 152600 375524 152652
rect 405556 152600 405608 152652
rect 405648 152600 405700 152652
rect 428004 152600 428056 152652
rect 428464 152600 428516 152652
rect 446036 152600 446088 152652
rect 446956 152600 447008 152652
rect 345664 152532 345716 152584
rect 352288 152532 352340 152584
rect 352380 152532 352432 152584
rect 385040 152532 385092 152584
rect 385500 152532 385552 152584
rect 387616 152532 387668 152584
rect 393136 152532 393188 152584
rect 419080 152532 419132 152584
rect 419264 152532 419316 152584
rect 433432 152532 433484 152584
rect 433524 152532 433576 152584
rect 291844 152464 291896 152516
rect 336832 152464 336884 152516
rect 339500 152464 339552 152516
rect 377312 152464 377364 152516
rect 378232 152464 378284 152516
rect 379888 152464 379940 152516
rect 382188 152464 382240 152516
rect 410708 152464 410760 152516
rect 56232 152396 56284 152448
rect 141056 152396 141108 152448
rect 144092 152396 144144 152448
rect 60004 152328 60056 152380
rect 144276 152328 144328 152380
rect 149060 152396 149112 152448
rect 231584 152396 231636 152448
rect 245108 152396 245160 152448
rect 306012 152396 306064 152448
rect 307300 152396 307352 152448
rect 345664 152396 345716 152448
rect 345756 152396 345808 152448
rect 346676 152396 346728 152448
rect 162216 152328 162268 152380
rect 164424 152328 164476 152380
rect 244372 152328 244424 152380
rect 255412 152328 255464 152380
rect 313096 152328 313148 152380
rect 313188 152328 313240 152380
rect 356152 152396 356204 152448
rect 354496 152328 354548 152380
rect 389548 152396 389600 152448
rect 389640 152396 389692 152448
rect 412640 152396 412692 152448
rect 364524 152328 364576 152380
rect 369032 152328 369084 152380
rect 371332 152328 371384 152380
rect 402336 152328 402388 152380
rect 405832 152328 405884 152380
rect 408776 152328 408828 152380
rect 409144 152328 409196 152380
rect 76748 152260 76800 152312
rect 159640 152260 159692 152312
rect 172612 152260 172664 152312
rect 249524 152260 249576 152312
rect 265348 152260 265400 152312
rect 270868 152260 270920 152312
rect 272524 152260 272576 152312
rect 316316 152260 316368 152312
rect 320272 152260 320324 152312
rect 323400 152260 323452 152312
rect 323492 152260 323544 152312
rect 330392 152260 330444 152312
rect 330944 152260 330996 152312
rect 371516 152260 371568 152312
rect 381360 152260 381412 152312
rect 410064 152260 410116 152312
rect 410892 152328 410944 152380
rect 431224 152464 431276 152516
rect 431316 152464 431368 152516
rect 436744 152464 436796 152516
rect 418436 152396 418488 152448
rect 438308 152464 438360 152516
rect 438492 152532 438544 152584
rect 440976 152532 441028 152584
rect 441436 152532 441488 152584
rect 455696 152532 455748 152584
rect 459652 152600 459704 152652
rect 465264 152600 465316 152652
rect 460112 152532 460164 152584
rect 449900 152464 449952 152516
rect 437756 152396 437808 152448
rect 453120 152396 453172 152448
rect 428648 152328 428700 152380
rect 431040 152328 431092 152380
rect 447968 152328 448020 152380
rect 423588 152260 423640 152312
rect 426256 152260 426308 152312
rect 426348 152260 426400 152312
rect 431316 152260 431368 152312
rect 85488 152192 85540 152244
rect 164792 152192 164844 152244
rect 167000 152192 167052 152244
rect 182732 152192 182784 152244
rect 183100 152192 183152 152244
rect 195612 152192 195664 152244
rect 75092 152124 75144 152176
rect 154488 152124 154540 152176
rect 156052 152124 156104 152176
rect 172520 152124 172572 152176
rect 176660 152124 176712 152176
rect 190460 152124 190512 152176
rect 195152 152124 195204 152176
rect 218704 152192 218756 152244
rect 221464 152192 221516 152244
rect 282920 152192 282972 152244
rect 285496 152192 285548 152244
rect 291844 152192 291896 152244
rect 292488 152192 292540 152244
rect 341984 152192 342036 152244
rect 342260 152192 342312 152244
rect 346492 152192 346544 152244
rect 346584 152192 346636 152244
rect 380532 152192 380584 152244
rect 384948 152192 385000 152244
rect 392124 152192 392176 152244
rect 394332 152192 394384 152244
rect 417792 152192 417844 152244
rect 417884 152192 417936 152244
rect 421748 152192 421800 152244
rect 423404 152192 423456 152244
rect 442172 152260 442224 152312
rect 431500 152192 431552 152244
rect 441528 152192 441580 152244
rect 441988 152192 442040 152244
rect 456340 152260 456392 152312
rect 443644 152192 443696 152244
rect 457628 152192 457680 152244
rect 71780 152056 71832 152108
rect 149428 152056 149480 152108
rect 150440 152056 150492 152108
rect 167368 152056 167420 152108
rect 169760 152056 169812 152108
rect 185308 152056 185360 152108
rect 193128 152056 193180 152108
rect 213552 152124 213604 152176
rect 213736 152124 213788 152176
rect 274548 152124 274600 152176
rect 277952 152124 278004 152176
rect 331128 152124 331180 152176
rect 331864 152124 331916 152176
rect 372160 152124 372212 152176
rect 388352 152124 388404 152176
rect 407488 152124 407540 152176
rect 415124 152124 415176 152176
rect 423588 152124 423640 152176
rect 427084 152124 427136 152176
rect 433800 152124 433852 152176
rect 436744 152124 436796 152176
rect 444104 152124 444156 152176
rect 445668 152124 445720 152176
rect 458824 152124 458876 152176
rect 516692 152124 516744 152176
rect 520280 152124 520332 152176
rect 195888 152056 195940 152108
rect 208492 152056 208544 152108
rect 109684 151988 109736 152040
rect 128176 151988 128228 152040
rect 128360 151988 128412 152040
rect 203340 151988 203392 152040
rect 212632 151988 212684 152040
rect 272708 152056 272760 152108
rect 272800 152056 272852 152108
rect 325976 152056 326028 152108
rect 330392 152056 330444 152108
rect 362592 152056 362644 152108
rect 388444 152056 388496 152108
rect 404912 152056 404964 152108
rect 405372 152056 405424 152108
rect 421012 152056 421064 152108
rect 242440 151988 242492 152040
rect 300952 151988 301004 152040
rect 304816 151988 304868 152040
rect 351644 151988 351696 152040
rect 352748 151988 352800 152040
rect 388260 151988 388312 152040
rect 403440 151988 403492 152040
rect 418436 151988 418488 152040
rect 426808 152056 426860 152108
rect 426900 152056 426952 152108
rect 444748 152056 444800 152108
rect 515496 152056 515548 152108
rect 518992 152056 519044 152108
rect 107568 151920 107620 151972
rect 175096 151920 175148 151972
rect 185584 151920 185636 151972
rect 200764 151920 200816 151972
rect 243360 151920 243412 151972
rect 302884 151920 302936 151972
rect 30196 151852 30248 151904
rect 74540 151852 74592 151904
rect 109132 151852 109184 151904
rect 138480 151852 138532 151904
rect 138572 151852 138624 151904
rect 146852 151852 146904 151904
rect 33600 151784 33652 151836
rect 84200 151784 84252 151836
rect 105820 151784 105872 151836
rect 110328 151784 110380 151836
rect 113916 151784 113968 151836
rect 123484 151784 123536 151836
rect 138020 151784 138072 151836
rect 141792 151784 141844 151836
rect 143264 151784 143316 151836
rect 157064 151852 157116 151904
rect 160192 151852 160244 151904
rect 177672 151852 177724 151904
rect 191656 151852 191708 151904
rect 195888 151852 195940 151904
rect 272616 151852 272668 151904
rect 326620 151920 326672 151972
rect 325056 151852 325108 151904
rect 343824 151852 343876 151904
rect 346584 151852 346636 151904
rect 346676 151852 346728 151904
rect 352472 151852 352524 151904
rect 261024 151784 261076 151836
rect 272524 151784 272576 151836
rect 283012 151784 283064 151836
rect 287428 151784 287480 151836
rect 303988 151784 304040 151836
rect 351000 151784 351052 151836
rect 362960 151920 363012 151972
rect 364524 151920 364576 151972
rect 386236 151920 386288 151972
rect 399760 151920 399812 151972
rect 399852 151920 399904 151972
rect 355324 151852 355376 151904
rect 390192 151852 390244 151904
rect 367008 151784 367060 151836
rect 378784 151784 378836 151836
rect 384396 151784 384448 151836
rect 385316 151784 385368 151836
rect 394700 151784 394752 151836
rect 396172 151784 396224 151836
rect 402980 151784 403032 151836
rect 413836 151920 413888 151972
rect 416504 151920 416556 151972
rect 416596 151920 416648 151972
rect 422576 151988 422628 152040
rect 431500 151988 431552 152040
rect 431592 151988 431644 152040
rect 439596 151988 439648 152040
rect 419540 151920 419592 151972
rect 437020 151920 437072 151972
rect 439412 151920 439464 151972
rect 454408 151988 454460 152040
rect 456800 151988 456852 152040
rect 463332 151988 463384 152040
rect 486516 151988 486568 152040
rect 490288 151988 490340 152040
rect 515956 151988 516008 152040
rect 519912 151988 519964 152040
rect 403900 151852 403952 151904
rect 415860 151852 415912 151904
rect 413284 151784 413336 151836
rect 413652 151784 413704 151836
rect 421656 151852 421708 151904
rect 421748 151852 421800 151904
rect 431868 151852 431920 151904
rect 433340 151852 433392 151904
rect 419632 151784 419684 151836
rect 434444 151784 434496 151836
rect 436100 151852 436152 151904
rect 451832 151920 451884 151972
rect 456064 151920 456116 151972
rect 461400 151920 461452 151972
rect 469220 151920 469272 151972
rect 472348 151920 472400 151972
rect 487344 151920 487396 151972
rect 490932 151920 490984 151972
rect 507676 151920 507728 151972
rect 509240 151920 509292 151972
rect 517428 151920 517480 151972
rect 521568 151920 521620 151972
rect 440884 151852 440936 151904
rect 440976 151852 441028 151904
rect 451188 151852 451240 151904
rect 457168 151852 457220 151904
rect 462688 151852 462740 151904
rect 468024 151852 468076 151904
rect 471060 151852 471112 151904
rect 489092 151852 489144 151904
rect 492220 151852 492272 151904
rect 499488 151852 499540 151904
rect 499948 151852 500000 151904
rect 440240 151784 440292 151836
rect 455052 151784 455104 151836
rect 455788 151784 455840 151836
rect 462044 151784 462096 151836
rect 467932 151784 467984 151836
rect 471704 151784 471756 151836
rect 488448 151784 488500 151836
rect 491576 151784 491628 151836
rect 509056 151784 509108 151836
rect 510896 151784 510948 151836
rect 84200 151376 84252 151428
rect 117228 151376 117280 151428
rect 74540 151308 74592 151360
rect 117136 151308 117188 151360
rect 68008 151240 68060 151292
rect 112812 151240 112864 151292
rect 64512 151172 64564 151224
rect 112720 151172 112772 151224
rect 61108 151104 61160 151156
rect 112628 151104 112680 151156
rect 57704 151036 57756 151088
rect 112536 151036 112588 151088
rect 54208 150968 54260 151020
rect 111616 150968 111668 151020
rect 50804 150900 50856 150952
rect 112444 150900 112496 150952
rect 47308 150832 47360 150884
rect 111524 150832 111576 150884
rect 43904 150764 43956 150816
rect 111432 150764 111484 150816
rect 40500 150696 40552 150748
rect 111340 150696 111392 150748
rect 37004 150628 37056 150680
rect 111248 150628 111300 150680
rect 19800 150560 19852 150612
rect 116860 150560 116912 150612
rect 16396 150492 16448 150544
rect 116768 150492 116820 150544
rect 2688 150424 2740 150476
rect 111064 150424 111116 150476
rect 118424 150152 118476 150204
rect 121782 150152 121834 150204
rect 135444 150152 135496 150204
rect 136594 150152 136646 150204
rect 146392 150152 146444 150204
rect 147542 150152 147594 150204
rect 147680 150152 147732 150204
rect 148830 150152 148882 150204
rect 164332 150152 164384 150204
rect 165482 150152 165534 150204
rect 165620 150152 165672 150204
rect 166770 150152 166822 150204
rect 171140 150152 171192 150204
rect 171922 150152 171974 150204
rect 182272 150152 182324 150204
rect 183422 150152 183474 150204
rect 183560 150152 183612 150204
rect 184710 150152 184762 150204
rect 200304 150152 200356 150204
rect 201454 150152 201506 150204
rect 204260 150152 204312 150204
rect 205318 150152 205370 150204
rect 211252 150152 211304 150204
rect 212310 150152 212362 150204
rect 218244 150152 218296 150204
rect 219394 150152 219446 150204
rect 229192 150152 229244 150204
rect 230342 150152 230394 150204
rect 238852 150152 238904 150204
rect 240002 150152 240054 150204
rect 245844 150152 245896 150204
rect 246994 150152 247046 150204
rect 247132 150152 247184 150204
rect 248282 150152 248334 150204
rect 253940 150152 253992 150204
rect 254722 150152 254774 150204
rect 256792 150152 256844 150204
rect 257942 150152 257994 150204
rect 258080 150152 258132 150204
rect 259230 150152 259282 150204
rect 259460 150152 259512 150204
rect 260518 150152 260570 150204
rect 263600 150152 263652 150204
rect 264382 150152 264434 150204
rect 281540 150152 281592 150204
rect 282322 150152 282374 150204
rect 283104 150152 283156 150204
rect 284254 150152 284306 150204
rect 285680 150152 285732 150204
rect 286830 150152 286882 150204
rect 299480 150152 299532 150204
rect 300354 150152 300406 150204
rect 302424 150152 302476 150204
rect 303574 150152 303626 150204
rect 347964 150152 348016 150204
rect 349114 150152 349166 150204
rect 354680 150152 354732 150204
rect 355554 150152 355606 150204
rect 358912 150152 358964 150204
rect 360062 150152 360114 150204
rect 369860 150152 369912 150204
rect 370918 150152 370970 150204
rect 375564 150152 375616 150204
rect 376714 150152 376766 150204
rect 378140 150152 378192 150204
rect 379290 150152 379342 150204
rect 394884 150152 394936 150204
rect 396034 150152 396086 150204
rect 403164 150152 403216 150204
rect 404314 150152 404366 150204
rect 477684 150152 477736 150204
rect 478834 150152 478886 150204
rect 478972 150152 479024 150204
rect 480122 150152 480174 150204
rect 481640 150152 481692 150204
rect 482698 150152 482750 150204
rect 6368 150016 6420 150068
rect 111156 150016 111208 150068
rect 23388 149948 23440 150000
rect 116952 149948 117004 150000
rect 13360 149880 13412 149932
rect 116676 149880 116728 149932
rect 9588 149812 9640 149864
rect 116584 149812 116636 149864
rect 88984 149744 89036 149796
rect 114008 149744 114060 149796
rect 85488 149676 85540 149728
rect 113916 149676 113968 149728
rect 81992 149608 82044 149660
rect 112352 149608 112404 149660
rect 78588 149540 78640 149592
rect 113088 149540 113140 149592
rect 75184 149472 75236 149524
rect 112996 149472 113048 149524
rect 71688 149404 71740 149456
rect 112904 149404 112956 149456
rect 26976 149336 27028 149388
rect 117044 149336 117096 149388
rect 92296 149268 92348 149320
rect 102508 149268 102560 149320
rect 102692 149268 102744 149320
rect 102876 149268 102928 149320
rect 116216 149268 116268 149320
rect 116492 149200 116544 149252
rect 116032 149132 116084 149184
rect 114100 149064 114152 149116
rect 109592 148996 109644 149048
rect 115940 148996 115992 149048
rect 110328 147568 110380 147620
rect 116124 147568 116176 147620
rect 114100 140700 114152 140752
rect 115940 140700 115992 140752
rect 114008 137912 114060 137964
rect 116400 137912 116452 137964
rect 113916 136552 113968 136604
rect 115940 136552 115992 136604
rect 112352 133832 112404 133884
rect 116124 133832 116176 133884
rect 113088 132404 113140 132456
rect 116124 132404 116176 132456
rect 112996 131044 113048 131096
rect 116124 131044 116176 131096
rect 112904 128256 112956 128308
rect 116124 128256 116176 128308
rect 112812 126896 112864 126948
rect 116032 126896 116084 126948
rect 112720 124108 112772 124160
rect 116124 124108 116176 124160
rect 112628 122748 112680 122800
rect 115940 122748 115992 122800
rect 112536 121388 112588 121440
rect 116124 121388 116176 121440
rect 111616 118600 111668 118652
rect 116124 118600 116176 118652
rect 116492 117988 116544 118040
rect 117228 117988 117280 118040
rect 112444 117240 112496 117292
rect 116124 117240 116176 117292
rect 111524 114452 111576 114504
rect 116124 114452 116176 114504
rect 111432 113092 111484 113144
rect 115940 113092 115992 113144
rect 111340 111732 111392 111784
rect 116124 111732 116176 111784
rect 111248 108944 111300 108996
rect 116124 108944 116176 108996
rect 111156 92420 111208 92472
rect 116124 92420 116176 92472
rect 111064 89632 111116 89684
rect 116124 89632 116176 89684
rect 113824 88272 113876 88324
rect 116032 88272 116084 88324
rect 114468 87184 114520 87236
rect 116492 87184 116544 87236
rect 113916 86912 113968 86964
rect 116216 86912 116268 86964
rect 114008 83920 114060 83972
rect 116584 83920 116636 83972
rect 114100 82764 114152 82816
rect 116308 82764 116360 82816
rect 114192 79976 114244 80028
rect 115940 79976 115992 80028
rect 114192 71748 114244 71800
rect 116584 71748 116636 71800
rect 114100 69028 114152 69080
rect 116308 69028 116360 69080
rect 114008 67600 114060 67652
rect 116124 67600 116176 67652
rect 113916 66240 113968 66292
rect 116584 66240 116636 66292
rect 114468 64540 114520 64592
rect 116584 64540 116636 64592
rect 113824 63520 113876 63572
rect 116216 63520 116268 63572
rect 109684 41420 109736 41472
rect 116124 41420 116176 41472
rect 114100 38632 114152 38684
rect 116400 38632 116452 38684
rect 116216 38496 116268 38548
rect 116400 38496 116452 38548
rect 114192 37272 114244 37324
rect 116216 37272 116268 37324
rect 111064 34484 111116 34536
rect 116124 34484 116176 34536
rect 112444 33124 112496 33176
rect 116124 33124 116176 33176
rect 112536 31764 112588 31816
rect 116124 31764 116176 31816
rect 112628 28976 112680 29028
rect 116124 28976 116176 29028
rect 112720 27616 112772 27668
rect 116124 27616 116176 27668
rect 112812 24828 112864 24880
rect 116124 24828 116176 24880
rect 111156 23468 111208 23520
rect 116124 23468 116176 23520
rect 111248 22108 111300 22160
rect 116032 22108 116084 22160
rect 116032 16464 116084 16516
rect 116216 16464 116268 16516
rect 116216 11840 116268 11892
rect 116308 11636 116360 11688
rect 116952 11364 117004 11416
rect 117320 11364 117372 11416
rect 116952 5448 117004 5500
rect 117136 5448 117188 5500
rect 116308 5312 116360 5364
rect 116952 5312 117004 5364
rect 115940 5176 115992 5228
rect 116308 5176 116360 5228
rect 115940 5040 115992 5092
rect 116124 5040 116176 5092
rect 109776 4156 109828 4208
rect 116124 4156 116176 4208
rect 2504 2864 2556 2916
rect 32772 2592 32824 2644
rect 39120 2592 39172 2644
rect 39672 2592 39724 2644
rect 40316 2592 40368 2644
rect 47492 2592 47544 2644
rect 49148 2592 49200 2644
rect 49608 2592 49660 2644
rect 50896 2592 50948 2644
rect 53012 2592 53064 2644
rect 36360 2456 36412 2508
rect 40316 2456 40368 2508
rect 46296 2524 46348 2576
rect 111064 3884 111116 3936
rect 112444 3816 112496 3868
rect 53472 2592 53524 2644
rect 53656 2592 53708 2644
rect 57520 2592 57572 2644
rect 58624 2592 58676 2644
rect 58716 2592 58768 2644
rect 62396 2592 62448 2644
rect 62764 2592 62816 2644
rect 63040 2592 63092 2644
rect 63132 2592 63184 2644
rect 65524 2592 65576 2644
rect 56232 2524 56284 2576
rect 73988 2524 74040 2576
rect 74080 2524 74132 2576
rect 76656 2524 76708 2576
rect 78036 2592 78088 2644
rect 78128 2592 78180 2644
rect 112536 3748 112588 3800
rect 112628 3680 112680 3732
rect 112720 3612 112772 3664
rect 112812 3544 112864 3596
rect 111156 3476 111208 3528
rect 111248 3408 111300 3460
rect 114192 3340 114244 3392
rect 114100 3272 114152 3324
rect 78496 2592 78548 2644
rect 79692 2592 79744 2644
rect 79784 2592 79836 2644
rect 81164 2592 81216 2644
rect 81256 2592 81308 2644
rect 81348 2592 81400 2644
rect 82084 2592 82136 2644
rect 82176 2592 82228 2644
rect 82268 2592 82320 2644
rect 79416 2524 79468 2576
rect 79600 2524 79652 2576
rect 52920 2388 52972 2440
rect 53656 2388 53708 2440
rect 59728 2388 59780 2440
rect 65524 2388 65576 2440
rect 66352 2388 66404 2440
rect 82084 2388 82136 2440
rect 53012 2252 53064 2304
rect 81164 2320 81216 2372
rect 47492 2184 47544 2236
rect 76564 2252 76616 2304
rect 76656 2252 76708 2304
rect 109592 3000 109644 3052
rect 117964 3000 118016 3052
rect 117688 2932 117740 2984
rect 116124 2864 116176 2916
rect 98276 2592 98328 2644
rect 106096 2592 106148 2644
rect 294788 2592 294840 2644
rect 425796 2592 425848 2644
rect 443644 2592 443696 2644
rect 491300 2592 491352 2644
rect 493600 2592 493652 2644
rect 109592 2456 109644 2508
rect 116584 2456 116636 2508
rect 106188 2388 106240 2440
rect 116676 2388 116728 2440
rect 102968 2320 103020 2372
rect 116768 2320 116820 2372
rect 99656 2252 99708 2304
rect 116860 2252 116912 2304
rect 58716 2184 58768 2236
rect 63132 2184 63184 2236
rect 69664 2184 69716 2236
rect 82176 2184 82228 2236
rect 96344 2184 96396 2236
rect 117044 2184 117096 2236
rect 57520 2116 57572 2168
rect 76564 2116 76616 2168
rect 81348 2116 81400 2168
rect 93032 2116 93084 2168
rect 117228 2116 117280 2168
rect 78496 2048 78548 2100
rect 89628 2048 89680 2100
rect 117320 2048 117372 2100
rect 86408 1980 86460 2032
rect 117136 1980 117188 2032
rect 82636 1912 82688 1964
rect 116492 1912 116544 1964
rect 79324 1844 79376 1896
rect 116400 1844 116452 1896
rect 72700 1776 72752 1828
rect 109684 1776 109736 1828
rect 76012 1708 76064 1760
rect 116216 1708 116268 1760
rect 32680 1640 32732 1692
rect 116032 1640 116084 1692
rect 29276 1572 29328 1624
rect 115940 1572 115992 1624
rect 25964 1504 26016 1556
rect 116952 1504 117004 1556
rect 22652 1436 22704 1488
rect 116308 1436 116360 1488
rect 117688 1436 117740 1488
rect 143632 1436 143684 1488
rect 6000 1368 6052 1420
rect 109776 1368 109828 1420
rect 117964 1368 118016 1420
rect 193588 1368 193640 1420
rect 294788 1368 294840 1420
rect 343640 1368 343692 1420
<< metal2 >>
rect 386 163200 442 164400
rect 1214 163200 1270 164400
rect 2042 163200 2098 164400
rect 2870 163200 2926 164400
rect 3698 163200 3754 164400
rect 3804 163254 4016 163282
rect 400 158030 428 163200
rect 388 158024 440 158030
rect 388 157966 440 157972
rect 1228 153950 1256 163200
rect 2056 156670 2084 163200
rect 2044 156664 2096 156670
rect 2044 156606 2096 156612
rect 1216 153944 1268 153950
rect 1216 153886 1268 153892
rect 2884 152522 2912 163200
rect 3712 163146 3740 163200
rect 3804 163146 3832 163254
rect 3712 163118 3832 163146
rect 3988 153882 4016 163254
rect 4526 163200 4582 164400
rect 5354 163200 5410 164400
rect 6274 163200 6330 164400
rect 7102 163200 7158 164400
rect 7930 163200 7986 164400
rect 8758 163200 8814 164400
rect 9586 163200 9642 164400
rect 10414 163200 10470 164400
rect 11242 163200 11298 164400
rect 12162 163200 12218 164400
rect 12990 163200 13046 164400
rect 13818 163200 13874 164400
rect 14646 163200 14702 164400
rect 15474 163200 15530 164400
rect 16302 163200 16358 164400
rect 17130 163200 17186 164400
rect 18050 163200 18106 164400
rect 18878 163200 18934 164400
rect 19706 163200 19762 164400
rect 20534 163200 20590 164400
rect 21362 163200 21418 164400
rect 22190 163200 22246 164400
rect 23018 163200 23074 164400
rect 23938 163200 23994 164400
rect 24766 163200 24822 164400
rect 25594 163200 25650 164400
rect 26422 163200 26478 164400
rect 27250 163200 27306 164400
rect 28078 163200 28134 164400
rect 28906 163200 28962 164400
rect 29826 163200 29882 164400
rect 30654 163200 30710 164400
rect 31482 163200 31538 164400
rect 32310 163200 32366 164400
rect 33138 163200 33194 164400
rect 33966 163200 34022 164400
rect 34794 163200 34850 164400
rect 35714 163200 35770 164400
rect 36542 163200 36598 164400
rect 37370 163200 37426 164400
rect 38198 163200 38254 164400
rect 38304 163254 38516 163282
rect 4540 155378 4568 163200
rect 4528 155372 4580 155378
rect 4528 155314 4580 155320
rect 5368 155242 5396 163200
rect 6288 159390 6316 163200
rect 6276 159384 6328 159390
rect 6276 159326 6328 159332
rect 5356 155236 5408 155242
rect 5356 155178 5408 155184
rect 7116 154018 7144 163200
rect 7944 155446 7972 163200
rect 7932 155440 7984 155446
rect 7932 155382 7984 155388
rect 8772 155310 8800 163200
rect 8760 155304 8812 155310
rect 8760 155246 8812 155252
rect 7104 154012 7156 154018
rect 7104 153954 7156 153960
rect 3976 153876 4028 153882
rect 3976 153818 4028 153824
rect 2872 152516 2924 152522
rect 2872 152458 2924 152464
rect 9600 152425 9628 163200
rect 10428 154086 10456 163200
rect 11256 156806 11284 163200
rect 11244 156800 11296 156806
rect 11244 156742 11296 156748
rect 12176 155854 12204 163200
rect 12164 155848 12216 155854
rect 12164 155790 12216 155796
rect 10416 154080 10468 154086
rect 10416 154022 10468 154028
rect 13004 152561 13032 163200
rect 13832 154154 13860 163200
rect 14660 156738 14688 163200
rect 14648 156732 14700 156738
rect 14648 156674 14700 156680
rect 13820 154148 13872 154154
rect 13820 154090 13872 154096
rect 15488 152658 15516 163200
rect 16316 159497 16344 163200
rect 16302 159488 16358 159497
rect 16302 159423 16358 159432
rect 17144 153921 17172 163200
rect 18064 156942 18092 163200
rect 18892 159730 18920 163200
rect 18880 159724 18932 159730
rect 18880 159666 18932 159672
rect 18052 156936 18104 156942
rect 18052 156878 18104 156884
rect 17130 153912 17186 153921
rect 17130 153847 17186 153856
rect 15476 152652 15528 152658
rect 15476 152594 15528 152600
rect 19720 152590 19748 163200
rect 20548 153785 20576 163200
rect 21376 156874 21404 163200
rect 21364 156868 21416 156874
rect 21364 156810 21416 156816
rect 20534 153776 20590 153785
rect 20534 153711 20590 153720
rect 22204 152726 22232 163200
rect 23032 159361 23060 163200
rect 23018 159352 23074 159361
rect 23018 159287 23074 159296
rect 23952 154222 23980 163200
rect 24780 157010 24808 163200
rect 25608 160002 25636 163200
rect 25596 159996 25648 160002
rect 25596 159938 25648 159944
rect 24768 157004 24820 157010
rect 24768 156946 24820 156952
rect 23940 154216 23992 154222
rect 23940 154158 23992 154164
rect 26436 152794 26464 163200
rect 27264 154057 27292 163200
rect 28092 156777 28120 163200
rect 28078 156768 28134 156777
rect 28078 156703 28134 156712
rect 28920 155514 28948 163200
rect 29840 159633 29868 163200
rect 29826 159624 29882 159633
rect 29826 159559 29882 159568
rect 28908 155508 28960 155514
rect 28908 155450 28960 155456
rect 30668 154290 30696 163200
rect 31496 156641 31524 163200
rect 32324 159594 32352 163200
rect 32312 159588 32364 159594
rect 32312 159530 32364 159536
rect 31482 156632 31538 156641
rect 31482 156567 31538 156576
rect 33152 155718 33180 163200
rect 33980 158001 34008 163200
rect 33966 157992 34022 158001
rect 33966 157927 34022 157936
rect 33140 155712 33192 155718
rect 33140 155654 33192 155660
rect 34808 154426 34836 163200
rect 35728 157078 35756 163200
rect 36556 159458 36584 163200
rect 36544 159452 36596 159458
rect 36544 159394 36596 159400
rect 37384 158098 37412 163200
rect 38212 163146 38240 163200
rect 38304 163146 38332 163254
rect 38212 163118 38332 163146
rect 37372 158092 37424 158098
rect 37372 158034 37424 158040
rect 35716 157072 35768 157078
rect 35716 157014 35768 157020
rect 34796 154420 34848 154426
rect 34796 154362 34848 154368
rect 38488 154358 38516 163254
rect 39026 163200 39082 164400
rect 39854 163200 39910 164400
rect 40682 163200 40738 164400
rect 41602 163200 41658 164400
rect 42430 163200 42486 164400
rect 43258 163200 43314 164400
rect 44086 163200 44142 164400
rect 44914 163200 44970 164400
rect 45742 163200 45798 164400
rect 46570 163200 46626 164400
rect 47490 163200 47546 164400
rect 48318 163200 48374 164400
rect 49146 163200 49202 164400
rect 49974 163200 50030 164400
rect 50802 163200 50858 164400
rect 51630 163200 51686 164400
rect 52458 163200 52514 164400
rect 53378 163200 53434 164400
rect 54206 163200 54262 164400
rect 55034 163200 55090 164400
rect 55862 163200 55918 164400
rect 56690 163200 56746 164400
rect 57518 163200 57574 164400
rect 58346 163200 58402 164400
rect 59266 163200 59322 164400
rect 60094 163200 60150 164400
rect 60922 163200 60978 164400
rect 61750 163200 61806 164400
rect 62578 163200 62634 164400
rect 63406 163200 63462 164400
rect 64234 163200 64290 164400
rect 65154 163200 65210 164400
rect 65982 163200 66038 164400
rect 66810 163200 66866 164400
rect 67638 163200 67694 164400
rect 68466 163200 68522 164400
rect 69294 163200 69350 164400
rect 70122 163200 70178 164400
rect 71042 163200 71098 164400
rect 71870 163200 71926 164400
rect 72698 163200 72754 164400
rect 73526 163200 73582 164400
rect 74354 163200 74410 164400
rect 75182 163200 75238 164400
rect 76010 163200 76066 164400
rect 76930 163200 76986 164400
rect 77758 163200 77814 164400
rect 78586 163200 78642 164400
rect 79414 163200 79470 164400
rect 80242 163200 80298 164400
rect 81070 163200 81126 164400
rect 81898 163200 81954 164400
rect 82818 163200 82874 164400
rect 83646 163200 83702 164400
rect 84474 163200 84530 164400
rect 85302 163200 85358 164400
rect 86130 163200 86186 164400
rect 86958 163200 87014 164400
rect 87786 163200 87842 164400
rect 88706 163200 88762 164400
rect 89534 163200 89590 164400
rect 90362 163200 90418 164400
rect 91190 163200 91246 164400
rect 92018 163200 92074 164400
rect 92846 163200 92902 164400
rect 93674 163200 93730 164400
rect 94594 163200 94650 164400
rect 95422 163200 95478 164400
rect 96250 163200 96306 164400
rect 97078 163200 97134 164400
rect 97906 163200 97962 164400
rect 98734 163200 98790 164400
rect 99562 163200 99618 164400
rect 100482 163200 100538 164400
rect 101310 163200 101366 164400
rect 102138 163200 102194 164400
rect 102966 163200 103022 164400
rect 103794 163200 103850 164400
rect 104622 163200 104678 164400
rect 105450 163200 105506 164400
rect 106370 163200 106426 164400
rect 107198 163200 107254 164400
rect 108026 163200 108082 164400
rect 108854 163200 108910 164400
rect 109682 163200 109738 164400
rect 110510 163200 110566 164400
rect 111338 163200 111394 164400
rect 112258 163200 112314 164400
rect 113086 163200 113142 164400
rect 113914 163200 113970 164400
rect 114742 163200 114798 164400
rect 115570 163200 115626 164400
rect 116398 163200 116454 164400
rect 117226 163200 117282 164400
rect 118146 163200 118202 164400
rect 118974 163200 119030 164400
rect 119802 163200 119858 164400
rect 120630 163200 120686 164400
rect 121458 163200 121514 164400
rect 122286 163200 122342 164400
rect 123114 163200 123170 164400
rect 124034 163200 124090 164400
rect 124862 163200 124918 164400
rect 125690 163200 125746 164400
rect 126518 163200 126574 164400
rect 127346 163200 127402 164400
rect 128174 163200 128230 164400
rect 129002 163200 129058 164400
rect 129922 163200 129978 164400
rect 130750 163200 130806 164400
rect 131578 163200 131634 164400
rect 132406 163200 132462 164400
rect 133234 163200 133290 164400
rect 134062 163200 134118 164400
rect 134890 163200 134946 164400
rect 135810 163200 135866 164400
rect 136638 163200 136694 164400
rect 137466 163200 137522 164400
rect 138294 163200 138350 164400
rect 139122 163200 139178 164400
rect 139950 163200 140006 164400
rect 140778 163200 140834 164400
rect 141698 163200 141754 164400
rect 142526 163200 142582 164400
rect 143354 163200 143410 164400
rect 144182 163200 144238 164400
rect 145010 163200 145066 164400
rect 145116 163254 145328 163282
rect 39040 157146 39068 163200
rect 39028 157140 39080 157146
rect 39028 157082 39080 157088
rect 39868 155582 39896 163200
rect 40696 158273 40724 163200
rect 40682 158264 40738 158273
rect 40682 158199 40738 158208
rect 39856 155576 39908 155582
rect 39856 155518 39908 155524
rect 41616 154494 41644 163200
rect 42444 156913 42472 163200
rect 43272 159526 43300 163200
rect 43260 159520 43312 159526
rect 43260 159462 43312 159468
rect 44100 158137 44128 163200
rect 44086 158128 44142 158137
rect 44086 158063 44142 158072
rect 42430 156904 42486 156913
rect 42430 156839 42486 156848
rect 44928 154562 44956 163200
rect 45756 157214 45784 163200
rect 45744 157208 45796 157214
rect 45744 157150 45796 157156
rect 46584 155650 46612 163200
rect 47504 158166 47532 163200
rect 47492 158160 47544 158166
rect 47492 158102 47544 158108
rect 46572 155644 46624 155650
rect 46572 155586 46624 155592
rect 44916 154556 44968 154562
rect 44916 154498 44968 154504
rect 41604 154488 41656 154494
rect 41604 154430 41656 154436
rect 38476 154352 38528 154358
rect 38476 154294 38528 154300
rect 30656 154284 30708 154290
rect 30656 154226 30708 154232
rect 27250 154048 27306 154057
rect 27250 153983 27306 153992
rect 48332 153814 48360 163200
rect 49160 157049 49188 163200
rect 49988 159662 50016 163200
rect 49976 159656 50028 159662
rect 49976 159598 50028 159604
rect 50816 158234 50844 163200
rect 50804 158228 50856 158234
rect 50804 158170 50856 158176
rect 49146 157040 49202 157049
rect 49146 156975 49202 156984
rect 51644 154193 51672 163200
rect 52472 157282 52500 163200
rect 52460 157276 52512 157282
rect 52460 157218 52512 157224
rect 53392 155786 53420 163200
rect 54220 158302 54248 163200
rect 54208 158296 54260 158302
rect 54208 158238 54260 158244
rect 53380 155780 53432 155786
rect 53380 155722 53432 155728
rect 55048 154329 55076 163200
rect 55876 157350 55904 163200
rect 56704 159866 56732 163200
rect 56692 159860 56744 159866
rect 56692 159802 56744 159808
rect 57532 158409 57560 163200
rect 57518 158400 57574 158409
rect 57518 158335 57574 158344
rect 55864 157344 55916 157350
rect 55864 157286 55916 157292
rect 56232 155508 56284 155514
rect 56232 155450 56284 155456
rect 55034 154320 55090 154329
rect 55034 154255 55090 154264
rect 51630 154184 51686 154193
rect 51630 154119 51686 154128
rect 48320 153808 48372 153814
rect 48320 153750 48372 153756
rect 26424 152788 26476 152794
rect 26424 152730 26476 152736
rect 22192 152720 22244 152726
rect 22192 152662 22244 152668
rect 19708 152584 19760 152590
rect 12990 152552 13046 152561
rect 19708 152526 19760 152532
rect 12990 152487 13046 152496
rect 56244 152454 56272 155450
rect 58360 153746 58388 163200
rect 59280 155990 59308 163200
rect 59268 155984 59320 155990
rect 59268 155926 59320 155932
rect 60108 155922 60136 163200
rect 60936 158370 60964 163200
rect 60924 158364 60976 158370
rect 60924 158306 60976 158312
rect 60096 155916 60148 155922
rect 60096 155858 60148 155864
rect 60004 155712 60056 155718
rect 60004 155654 60056 155660
rect 58348 153740 58400 153746
rect 58348 153682 58400 153688
rect 56232 152448 56284 152454
rect 9586 152416 9642 152425
rect 56232 152390 56284 152396
rect 60016 152386 60044 155654
rect 61764 155281 61792 163200
rect 62592 155514 62620 163200
rect 63420 159798 63448 163200
rect 63408 159792 63460 159798
rect 63408 159734 63460 159740
rect 64248 158438 64276 163200
rect 64236 158432 64288 158438
rect 64236 158374 64288 158380
rect 62580 155508 62632 155514
rect 62580 155450 62632 155456
rect 61750 155272 61806 155281
rect 61750 155207 61806 155216
rect 65168 153678 65196 163200
rect 65996 157185 66024 163200
rect 65982 157176 66038 157185
rect 65982 157111 66038 157120
rect 65156 153672 65208 153678
rect 65156 153614 65208 153620
rect 66824 152862 66852 163200
rect 67652 158642 67680 163200
rect 67640 158636 67692 158642
rect 67640 158578 67692 158584
rect 68480 155417 68508 163200
rect 69308 155553 69336 163200
rect 70136 159934 70164 163200
rect 70124 159928 70176 159934
rect 70124 159870 70176 159876
rect 71056 158574 71084 163200
rect 71044 158568 71096 158574
rect 71044 158510 71096 158516
rect 71884 155718 71912 163200
rect 72712 156534 72740 163200
rect 73540 158982 73568 163200
rect 73528 158976 73580 158982
rect 73528 158918 73580 158924
rect 74368 158506 74396 163200
rect 74356 158500 74408 158506
rect 74356 158442 74408 158448
rect 72700 156528 72752 156534
rect 72700 156470 72752 156476
rect 71872 155712 71924 155718
rect 71872 155654 71924 155660
rect 75196 155650 75224 163200
rect 76024 155689 76052 163200
rect 76944 159322 76972 163200
rect 76932 159316 76984 159322
rect 76932 159258 76984 159264
rect 77772 157962 77800 163200
rect 77760 157956 77812 157962
rect 77760 157898 77812 157904
rect 76748 155780 76800 155786
rect 76748 155722 76800 155728
rect 76010 155680 76066 155689
rect 75092 155644 75144 155650
rect 75092 155586 75144 155592
rect 75184 155644 75236 155650
rect 76010 155615 76066 155624
rect 75184 155586 75236 155592
rect 71780 155576 71832 155582
rect 69294 155544 69350 155553
rect 71780 155518 71832 155524
rect 69294 155479 69350 155488
rect 68466 155408 68522 155417
rect 68466 155343 68522 155352
rect 66812 152856 66864 152862
rect 66812 152798 66864 152804
rect 9586 152351 9642 152360
rect 60004 152380 60056 152386
rect 60004 152322 60056 152328
rect 71792 152114 71820 155518
rect 75104 152182 75132 155586
rect 76760 152318 76788 155722
rect 78600 155582 78628 163200
rect 79428 156466 79456 163200
rect 79416 156460 79468 156466
rect 79416 156402 79468 156408
rect 78588 155576 78640 155582
rect 78588 155518 78640 155524
rect 80256 154970 80284 163200
rect 81084 158710 81112 163200
rect 81072 158704 81124 158710
rect 81072 158646 81124 158652
rect 81912 155786 81940 163200
rect 81900 155780 81952 155786
rect 81900 155722 81952 155728
rect 80244 154964 80296 154970
rect 80244 154906 80296 154912
rect 82832 153610 82860 163200
rect 83660 160070 83688 163200
rect 83648 160064 83700 160070
rect 83648 160006 83700 160012
rect 84488 157894 84516 163200
rect 84476 157888 84528 157894
rect 84476 157830 84528 157836
rect 85316 155825 85344 163200
rect 85488 155916 85540 155922
rect 85488 155858 85540 155864
rect 85302 155816 85358 155825
rect 85302 155751 85358 155760
rect 82820 153604 82872 153610
rect 82820 153546 82872 153552
rect 76748 152312 76800 152318
rect 76748 152254 76800 152260
rect 85500 152250 85528 155858
rect 86144 155174 86172 163200
rect 86972 159186 87000 163200
rect 86960 159180 87012 159186
rect 86960 159122 87012 159128
rect 87800 157826 87828 163200
rect 87788 157820 87840 157826
rect 87788 157762 87840 157768
rect 88720 155922 88748 163200
rect 89548 158794 89576 163200
rect 89548 158766 89760 158794
rect 88708 155916 88760 155922
rect 88708 155858 88760 155864
rect 86132 155168 86184 155174
rect 86132 155110 86184 155116
rect 86868 154964 86920 154970
rect 86868 154906 86920 154912
rect 86880 153066 86908 154906
rect 89732 154465 89760 158766
rect 89718 154456 89774 154465
rect 89718 154391 89774 154400
rect 86868 153060 86920 153066
rect 86868 153002 86920 153008
rect 90376 152930 90404 163200
rect 91204 157758 91232 163200
rect 91192 157752 91244 157758
rect 91192 157694 91244 157700
rect 92032 155961 92060 163200
rect 92860 156398 92888 163200
rect 93688 159254 93716 163200
rect 93676 159248 93728 159254
rect 93676 159190 93728 159196
rect 94608 157690 94636 163200
rect 94596 157684 94648 157690
rect 94596 157626 94648 157632
rect 92848 156392 92900 156398
rect 92848 156334 92900 156340
rect 92018 155952 92074 155961
rect 92018 155887 92074 155896
rect 95436 155106 95464 163200
rect 96264 158914 96292 163200
rect 96252 158908 96304 158914
rect 96252 158850 96304 158856
rect 95424 155100 95476 155106
rect 95424 155042 95476 155048
rect 97092 152998 97120 163200
rect 97920 157622 97948 163200
rect 97908 157616 97960 157622
rect 97908 157558 97960 157564
rect 98748 155038 98776 163200
rect 98736 155032 98788 155038
rect 98736 154974 98788 154980
rect 99576 154970 99604 163200
rect 100496 159118 100524 163200
rect 100484 159112 100536 159118
rect 100484 159054 100536 159060
rect 101324 156330 101352 163200
rect 101312 156324 101364 156330
rect 101312 156266 101364 156272
rect 99564 154964 99616 154970
rect 99564 154906 99616 154912
rect 102152 153542 102180 163200
rect 102980 158778 103008 163200
rect 102968 158772 103020 158778
rect 102968 158714 103020 158720
rect 102140 153536 102192 153542
rect 102140 153478 102192 153484
rect 103808 153134 103836 163200
rect 104636 158545 104664 163200
rect 104622 158536 104678 158545
rect 104622 158471 104678 158480
rect 105464 153406 105492 163200
rect 106384 158778 106412 163200
rect 107108 159724 107160 159730
rect 107108 159666 107160 159672
rect 106372 158772 106424 158778
rect 106372 158714 106424 158720
rect 107120 154902 107148 159666
rect 107212 159050 107240 163200
rect 107200 159044 107252 159050
rect 107200 158986 107252 158992
rect 107568 158976 107620 158982
rect 107568 158918 107620 158924
rect 107108 154896 107160 154902
rect 107108 154838 107160 154844
rect 105452 153400 105504 153406
rect 105452 153342 105504 153348
rect 103796 153128 103848 153134
rect 103796 153070 103848 153076
rect 97080 152992 97132 152998
rect 97080 152934 97132 152940
rect 90364 152924 90416 152930
rect 90364 152866 90416 152872
rect 85488 152244 85540 152250
rect 85488 152186 85540 152192
rect 75092 152176 75144 152182
rect 75092 152118 75144 152124
rect 71780 152108 71832 152114
rect 71780 152050 71832 152056
rect 107580 151978 107608 158918
rect 108040 156262 108068 163200
rect 108028 156256 108080 156262
rect 108028 156198 108080 156204
rect 108868 153474 108896 163200
rect 109132 159996 109184 160002
rect 109132 159938 109184 159944
rect 108856 153468 108908 153474
rect 108856 153410 108908 153416
rect 107568 151972 107620 151978
rect 107568 151914 107620 151920
rect 109144 151910 109172 159938
rect 109696 159730 109724 163200
rect 109684 159724 109736 159730
rect 109684 159666 109736 159672
rect 109684 155848 109736 155854
rect 109684 155790 109736 155796
rect 109696 152046 109724 155790
rect 110524 154834 110552 163200
rect 111352 157554 111380 163200
rect 111340 157548 111392 157554
rect 111340 157490 111392 157496
rect 112272 155854 112300 163200
rect 113100 157321 113128 163200
rect 113086 157312 113142 157321
rect 113086 157247 113142 157256
rect 112260 155848 112312 155854
rect 112260 155790 112312 155796
rect 110512 154828 110564 154834
rect 110512 154770 110564 154776
rect 113824 153876 113876 153882
rect 113824 153818 113876 153824
rect 113836 153338 113864 153818
rect 113824 153332 113876 153338
rect 113824 153274 113876 153280
rect 109684 152040 109736 152046
rect 109684 151982 109736 151988
rect 30196 151904 30248 151910
rect 30196 151846 30248 151852
rect 74540 151904 74592 151910
rect 74540 151846 74592 151852
rect 109132 151904 109184 151910
rect 109132 151846 109184 151852
rect 19800 150612 19852 150618
rect 19800 150554 19852 150560
rect 16396 150544 16448 150550
rect 16396 150486 16448 150492
rect 2688 150476 2740 150482
rect 2688 150418 2740 150424
rect 2700 149940 2728 150418
rect 6368 150068 6420 150074
rect 6368 150010 6420 150016
rect 6380 149954 6408 150010
rect 6118 149926 6408 149954
rect 13018 149938 13400 149954
rect 16408 149940 16436 150486
rect 19812 149940 19840 150554
rect 23388 150000 23440 150006
rect 23322 149948 23388 149954
rect 23322 149942 23440 149948
rect 13018 149932 13412 149938
rect 13018 149926 13360 149932
rect 23322 149926 23428 149942
rect 30208 149940 30236 151846
rect 33600 151836 33652 151842
rect 33600 151778 33652 151784
rect 33612 149940 33640 151778
rect 74552 151366 74580 151846
rect 113928 151842 113956 163200
rect 114756 157486 114784 163200
rect 114744 157480 114796 157486
rect 114744 157422 114796 157428
rect 115584 153882 115612 163200
rect 115572 153876 115624 153882
rect 115572 153818 115624 153824
rect 116412 153649 116440 163200
rect 117240 160002 117268 163200
rect 117228 159996 117280 160002
rect 117228 159938 117280 159944
rect 118160 156194 118188 163200
rect 118884 158024 118936 158030
rect 118884 157966 118936 157972
rect 118148 156188 118200 156194
rect 118148 156130 118200 156136
rect 118608 154012 118660 154018
rect 118608 153954 118660 153960
rect 118700 154012 118752 154018
rect 118700 153954 118752 153960
rect 118620 153882 118648 153954
rect 118712 153882 118740 153954
rect 118516 153876 118568 153882
rect 118516 153818 118568 153824
rect 118608 153876 118660 153882
rect 118608 153818 118660 153824
rect 118700 153876 118752 153882
rect 118700 153818 118752 153824
rect 116398 153640 116454 153649
rect 116398 153575 116454 153584
rect 118424 153332 118476 153338
rect 118424 153274 118476 153280
rect 84200 151836 84252 151842
rect 84200 151778 84252 151784
rect 105820 151836 105872 151842
rect 105820 151778 105872 151784
rect 110328 151836 110380 151842
rect 110328 151778 110380 151784
rect 113916 151836 113968 151842
rect 113916 151778 113968 151784
rect 84212 151434 84240 151778
rect 84200 151428 84252 151434
rect 84200 151370 84252 151376
rect 74540 151360 74592 151366
rect 74540 151302 74592 151308
rect 68008 151292 68060 151298
rect 68008 151234 68060 151240
rect 64512 151224 64564 151230
rect 64512 151166 64564 151172
rect 61108 151156 61160 151162
rect 61108 151098 61160 151104
rect 57704 151088 57756 151094
rect 57704 151030 57756 151036
rect 54208 151020 54260 151026
rect 54208 150962 54260 150968
rect 50804 150952 50856 150958
rect 50804 150894 50856 150900
rect 47308 150884 47360 150890
rect 47308 150826 47360 150832
rect 43904 150816 43956 150822
rect 43904 150758 43956 150764
rect 40500 150748 40552 150754
rect 40500 150690 40552 150696
rect 37004 150680 37056 150686
rect 37004 150622 37056 150628
rect 37016 149940 37044 150622
rect 40512 149940 40540 150690
rect 43916 149940 43944 150758
rect 47320 149940 47348 150826
rect 50816 149940 50844 150894
rect 54220 149940 54248 150962
rect 57716 149940 57744 151030
rect 61120 149940 61148 151098
rect 64524 149940 64552 151166
rect 68020 149940 68048 151234
rect 105832 149940 105860 151778
rect 13360 149874 13412 149880
rect 9588 149864 9640 149870
rect 9522 149812 9588 149818
rect 9522 149806 9640 149812
rect 9522 149790 9628 149806
rect 88642 149802 89024 149818
rect 88642 149796 89036 149802
rect 88642 149790 88984 149796
rect 88984 149738 89036 149744
rect 85488 149728 85540 149734
rect 81742 149666 82032 149682
rect 85238 149676 85488 149682
rect 85238 149670 85540 149676
rect 81742 149660 82044 149666
rect 81742 149654 81992 149660
rect 85238 149654 85528 149670
rect 81992 149602 82044 149608
rect 78588 149592 78640 149598
rect 74842 149530 75224 149546
rect 78338 149540 78588 149546
rect 95790 149560 95846 149569
rect 78338 149534 78640 149540
rect 74842 149524 75236 149530
rect 74842 149518 75184 149524
rect 78338 149518 78628 149534
rect 95542 149518 95790 149546
rect 95790 149495 95846 149504
rect 102690 149560 102746 149569
rect 102690 149495 102746 149504
rect 75184 149466 75236 149472
rect 71688 149456 71740 149462
rect 26726 149394 27016 149410
rect 71438 149404 71688 149410
rect 99286 149424 99342 149433
rect 71438 149398 71740 149404
rect 26726 149388 27028 149394
rect 26726 149382 26976 149388
rect 71438 149382 71728 149398
rect 92046 149382 92336 149410
rect 98946 149382 99286 149410
rect 26976 149330 27028 149336
rect 92308 149326 92336 149382
rect 102350 149382 102548 149410
rect 99286 149359 99342 149368
rect 102520 149326 102548 149382
rect 102704 149326 102732 149495
rect 102874 149424 102930 149433
rect 109250 149382 109632 149410
rect 102874 149359 102930 149368
rect 102888 149326 102916 149359
rect 92296 149320 92348 149326
rect 92296 149262 92348 149268
rect 102508 149320 102560 149326
rect 102508 149262 102560 149268
rect 102692 149320 102744 149326
rect 102692 149262 102744 149268
rect 102876 149320 102928 149326
rect 102876 149262 102928 149268
rect 109604 149054 109632 149382
rect 109592 149048 109644 149054
rect 109592 148990 109644 148996
rect 110340 147626 110368 151778
rect 117228 151428 117280 151434
rect 117228 151370 117280 151376
rect 117136 151360 117188 151366
rect 117136 151302 117188 151308
rect 112812 151292 112864 151298
rect 112812 151234 112864 151240
rect 112720 151224 112772 151230
rect 112720 151166 112772 151172
rect 112628 151156 112680 151162
rect 112628 151098 112680 151104
rect 112536 151088 112588 151094
rect 112536 151030 112588 151036
rect 111616 151020 111668 151026
rect 111616 150962 111668 150968
rect 111524 150884 111576 150890
rect 111524 150826 111576 150832
rect 111432 150816 111484 150822
rect 111432 150758 111484 150764
rect 111340 150748 111392 150754
rect 111340 150690 111392 150696
rect 111248 150680 111300 150686
rect 111248 150622 111300 150628
rect 111064 150476 111116 150482
rect 111064 150418 111116 150424
rect 110328 147620 110380 147626
rect 110328 147562 110380 147568
rect 111076 89690 111104 150418
rect 111156 150068 111208 150074
rect 111156 150010 111208 150016
rect 111168 92478 111196 150010
rect 111260 109002 111288 150622
rect 111352 111790 111380 150690
rect 111444 113150 111472 150758
rect 111536 114510 111564 150826
rect 111628 118658 111656 150962
rect 112444 150952 112496 150958
rect 112444 150894 112496 150900
rect 112352 149660 112404 149666
rect 112352 149602 112404 149608
rect 112364 133890 112392 149602
rect 112352 133884 112404 133890
rect 112352 133826 112404 133832
rect 111616 118652 111668 118658
rect 111616 118594 111668 118600
rect 112456 117298 112484 150894
rect 112548 121446 112576 151030
rect 112640 122806 112668 151098
rect 112732 124166 112760 151166
rect 112824 126954 112852 151234
rect 116860 150612 116912 150618
rect 116860 150554 116912 150560
rect 116768 150544 116820 150550
rect 116768 150486 116820 150492
rect 116676 149932 116728 149938
rect 116676 149874 116728 149880
rect 116584 149864 116636 149870
rect 116584 149806 116636 149812
rect 114008 149796 114060 149802
rect 114008 149738 114060 149744
rect 113916 149728 113968 149734
rect 113916 149670 113968 149676
rect 113088 149592 113140 149598
rect 113088 149534 113140 149540
rect 112996 149524 113048 149530
rect 112996 149466 113048 149472
rect 112904 149456 112956 149462
rect 112904 149398 112956 149404
rect 112916 128314 112944 149398
rect 113008 131102 113036 149466
rect 113100 132462 113128 149534
rect 113822 144256 113878 144265
rect 113822 144191 113878 144200
rect 113088 132456 113140 132462
rect 113088 132398 113140 132404
rect 112996 131096 113048 131102
rect 112996 131038 113048 131044
rect 112904 128308 112956 128314
rect 112904 128250 112956 128256
rect 112812 126948 112864 126954
rect 112812 126890 112864 126896
rect 112720 124160 112772 124166
rect 112720 124102 112772 124108
rect 112628 122800 112680 122806
rect 112628 122742 112680 122748
rect 112536 121440 112588 121446
rect 112536 121382 112588 121388
rect 112444 117292 112496 117298
rect 112444 117234 112496 117240
rect 111524 114504 111576 114510
rect 111524 114446 111576 114452
rect 111432 113144 111484 113150
rect 111432 113086 111484 113092
rect 111340 111784 111392 111790
rect 111340 111726 111392 111732
rect 111248 108996 111300 109002
rect 111248 108938 111300 108944
rect 111156 92472 111208 92478
rect 111156 92414 111208 92420
rect 111064 89684 111116 89690
rect 111064 89626 111116 89632
rect 113836 88330 113864 144191
rect 113928 136610 113956 149670
rect 114020 137970 114048 149738
rect 116216 149320 116268 149326
rect 116216 149262 116268 149268
rect 116032 149184 116084 149190
rect 116032 149126 116084 149132
rect 114100 149116 114152 149122
rect 114100 149058 114152 149064
rect 114112 140758 114140 149058
rect 115940 149048 115992 149054
rect 115938 149016 115940 149025
rect 115992 149016 115994 149025
rect 115938 148951 115994 148960
rect 116044 145217 116072 149126
rect 116124 147620 116176 147626
rect 116124 147562 116176 147568
rect 116136 147121 116164 147562
rect 116122 147112 116178 147121
rect 116122 147047 116178 147056
rect 116030 145208 116086 145217
rect 116030 145143 116086 145152
rect 116228 143313 116256 149262
rect 116492 149252 116544 149258
rect 116492 149194 116544 149200
rect 116214 143304 116270 143313
rect 116214 143239 116270 143248
rect 116504 141409 116532 149194
rect 116490 141400 116546 141409
rect 116490 141335 116546 141344
rect 114100 140752 114152 140758
rect 114100 140694 114152 140700
rect 115940 140752 115992 140758
rect 115940 140694 115992 140700
rect 115952 139505 115980 140694
rect 115938 139496 115994 139505
rect 115938 139431 115994 139440
rect 114008 137964 114060 137970
rect 114008 137906 114060 137912
rect 116400 137964 116452 137970
rect 116400 137906 116452 137912
rect 116412 137601 116440 137906
rect 116398 137592 116454 137601
rect 116398 137527 116454 137536
rect 113916 136604 113968 136610
rect 113916 136546 113968 136552
rect 115940 136604 115992 136610
rect 115940 136546 115992 136552
rect 115952 135561 115980 136546
rect 115938 135552 115994 135561
rect 115938 135487 115994 135496
rect 116124 133884 116176 133890
rect 116124 133826 116176 133832
rect 116136 133657 116164 133826
rect 116122 133648 116178 133657
rect 116122 133583 116178 133592
rect 113914 132832 113970 132841
rect 113914 132767 113970 132776
rect 113824 88324 113876 88330
rect 113824 88266 113876 88272
rect 113928 86970 113956 132767
rect 116124 132456 116176 132462
rect 116124 132398 116176 132404
rect 116136 131753 116164 132398
rect 116122 131744 116178 131753
rect 116122 131679 116178 131688
rect 116124 131096 116176 131102
rect 116124 131038 116176 131044
rect 116136 129849 116164 131038
rect 116122 129840 116178 129849
rect 116122 129775 116178 129784
rect 116124 128308 116176 128314
rect 116124 128250 116176 128256
rect 116136 127945 116164 128250
rect 116122 127936 116178 127945
rect 116122 127871 116178 127880
rect 116032 126948 116084 126954
rect 116032 126890 116084 126896
rect 116044 126041 116072 126890
rect 116030 126032 116086 126041
rect 116030 125967 116086 125976
rect 116124 124160 116176 124166
rect 116122 124128 116124 124137
rect 116176 124128 116178 124137
rect 116122 124063 116178 124072
rect 115940 122800 115992 122806
rect 115940 122742 115992 122748
rect 115952 122233 115980 122742
rect 115938 122224 115994 122233
rect 115938 122159 115994 122168
rect 116124 121440 116176 121446
rect 114006 121408 114062 121417
rect 116124 121382 116176 121388
rect 114006 121343 114062 121352
rect 113916 86964 113968 86970
rect 113916 86906 113968 86912
rect 114020 83978 114048 121343
rect 116136 120193 116164 121382
rect 116122 120184 116178 120193
rect 116122 120119 116178 120128
rect 116124 118652 116176 118658
rect 116124 118594 116176 118600
rect 116136 118289 116164 118594
rect 116122 118280 116178 118289
rect 116122 118215 116178 118224
rect 116492 118040 116544 118046
rect 116492 117982 116544 117988
rect 116124 117292 116176 117298
rect 116124 117234 116176 117240
rect 116136 116385 116164 117234
rect 116122 116376 116178 116385
rect 116122 116311 116178 116320
rect 116124 114504 116176 114510
rect 116122 114472 116124 114481
rect 116176 114472 116178 114481
rect 116122 114407 116178 114416
rect 115940 113144 115992 113150
rect 115940 113086 115992 113092
rect 115952 112577 115980 113086
rect 115938 112568 115994 112577
rect 115938 112503 115994 112512
rect 116124 111784 116176 111790
rect 116124 111726 116176 111732
rect 116136 110673 116164 111726
rect 116122 110664 116178 110673
rect 116122 110599 116178 110608
rect 114098 110120 114154 110129
rect 114098 110055 114154 110064
rect 114008 83972 114060 83978
rect 114008 83914 114060 83920
rect 114112 82822 114140 110055
rect 116124 108996 116176 109002
rect 116124 108938 116176 108944
rect 116136 108769 116164 108938
rect 116122 108760 116178 108769
rect 116122 108695 116178 108704
rect 116504 106865 116532 117982
rect 116490 106856 116546 106865
rect 116490 106791 116546 106800
rect 114190 98696 114246 98705
rect 114190 98631 114246 98640
rect 114100 82816 114152 82822
rect 114100 82758 114152 82764
rect 114204 80034 114232 98631
rect 116596 93401 116624 149806
rect 116688 95305 116716 149874
rect 116780 97209 116808 150486
rect 116872 99113 116900 150554
rect 116952 150000 117004 150006
rect 116952 149942 117004 149948
rect 116964 101017 116992 149942
rect 117044 149388 117096 149394
rect 117044 149330 117096 149336
rect 117056 102921 117084 149330
rect 117148 104825 117176 151302
rect 117240 118046 117268 151370
rect 118436 150210 118464 153274
rect 118528 153202 118556 153818
rect 118516 153196 118568 153202
rect 118516 153138 118568 153144
rect 118424 150204 118476 150210
rect 118424 150146 118476 150152
rect 118896 149954 118924 157966
rect 118988 154698 119016 163200
rect 119816 158982 119844 163200
rect 119804 158976 119856 158982
rect 119804 158918 119856 158924
rect 120538 158944 120594 158953
rect 120644 158914 120672 163200
rect 120538 158879 120540 158888
rect 120592 158879 120594 158888
rect 120632 158908 120684 158914
rect 120540 158850 120592 158856
rect 120632 158850 120684 158856
rect 121184 158908 121236 158914
rect 121184 158850 121236 158856
rect 120448 156664 120500 156670
rect 120448 156606 120500 156612
rect 118976 154692 119028 154698
rect 118976 154634 119028 154640
rect 119804 153944 119856 153950
rect 119804 153886 119856 153892
rect 119434 153640 119490 153649
rect 119434 153575 119490 153584
rect 119448 153270 119476 153575
rect 119436 153264 119488 153270
rect 119436 153206 119488 153212
rect 119816 150090 119844 153886
rect 120460 150090 120488 156606
rect 120632 154080 120684 154086
rect 120684 154028 120764 154034
rect 120632 154022 120764 154028
rect 120644 154006 120764 154022
rect 120736 153950 120764 154006
rect 120724 153944 120776 153950
rect 120724 153886 120776 153892
rect 120724 153332 120776 153338
rect 120724 153274 120776 153280
rect 120736 153202 120764 153274
rect 120724 153196 120776 153202
rect 120724 153138 120776 153144
rect 121196 152522 121224 158850
rect 121472 156670 121500 163200
rect 121550 158944 121606 158953
rect 121550 158879 121606 158888
rect 121460 156664 121512 156670
rect 121460 156606 121512 156612
rect 121564 154154 121592 158879
rect 122012 155440 122064 155446
rect 122012 155382 122064 155388
rect 121920 155372 121972 155378
rect 121920 155314 121972 155320
rect 121932 154630 121960 155314
rect 122024 154766 122052 155382
rect 122300 155378 122328 163200
rect 123128 159390 123156 163200
rect 122656 159384 122708 159390
rect 122656 159326 122708 159332
rect 123116 159384 123168 159390
rect 123116 159326 123168 159332
rect 122668 159225 122696 159326
rect 122654 159216 122710 159225
rect 122654 159151 122710 159160
rect 122838 159216 122894 159225
rect 122838 159151 122894 159160
rect 122852 157334 122880 159151
rect 124048 158914 124076 163200
rect 124036 158908 124088 158914
rect 124036 158850 124088 158856
rect 122852 157306 123708 157334
rect 122288 155372 122340 155378
rect 122288 155314 122340 155320
rect 123024 155236 123076 155242
rect 123024 155178 123076 155184
rect 122012 154760 122064 154766
rect 122012 154702 122064 154708
rect 121920 154624 121972 154630
rect 121920 154566 121972 154572
rect 122380 154624 122432 154630
rect 122380 154566 122432 154572
rect 121552 154148 121604 154154
rect 121552 154090 121604 154096
rect 121092 152516 121144 152522
rect 121092 152458 121144 152464
rect 121184 152516 121236 152522
rect 121184 152458 121236 152464
rect 121104 150090 121132 152458
rect 121782 150204 121834 150210
rect 121782 150146 121834 150152
rect 119816 150062 119890 150090
rect 120460 150062 120534 150090
rect 121104 150062 121178 150090
rect 118896 149926 119324 149954
rect 119862 149940 119890 150062
rect 120506 149940 120534 150062
rect 121150 149940 121178 150062
rect 121794 149940 121822 150146
rect 122392 150090 122420 154566
rect 123036 150090 123064 155178
rect 123484 153196 123536 153202
rect 123484 153138 123536 153144
rect 123496 151842 123524 153138
rect 123484 151836 123536 151842
rect 123484 151778 123536 151784
rect 123680 150226 123708 157306
rect 124876 156126 124904 163200
rect 125508 158840 125560 158846
rect 125508 158782 125560 158788
rect 124864 156120 124916 156126
rect 124864 156062 124916 156068
rect 124956 154760 125008 154766
rect 124956 154702 125008 154708
rect 124404 154692 124456 154698
rect 124404 154634 124456 154640
rect 124416 154018 124444 154634
rect 124312 154012 124364 154018
rect 124312 153954 124364 153960
rect 124404 154012 124456 154018
rect 124404 153954 124456 153960
rect 123680 150198 123754 150226
rect 122392 150062 122466 150090
rect 123036 150062 123110 150090
rect 122438 149940 122466 150062
rect 123082 149940 123110 150062
rect 123726 149940 123754 150198
rect 124324 150090 124352 153954
rect 124968 150090 124996 154702
rect 125520 153882 125548 158782
rect 125600 155440 125652 155446
rect 125600 155382 125652 155388
rect 125508 153876 125560 153882
rect 125508 153818 125560 153824
rect 125612 150090 125640 155382
rect 125704 155310 125732 163200
rect 126428 159588 126480 159594
rect 126428 159530 126480 159536
rect 125692 155304 125744 155310
rect 125692 155246 125744 155252
rect 126440 152697 126468 159530
rect 126532 158778 126560 163200
rect 126612 159588 126664 159594
rect 126612 159530 126664 159536
rect 126624 158982 126652 159530
rect 127070 159488 127126 159497
rect 127070 159423 127126 159432
rect 126612 158976 126664 158982
rect 126612 158918 126664 158924
rect 126520 158772 126572 158778
rect 126520 158714 126572 158720
rect 126888 153944 126940 153950
rect 126888 153886 126940 153892
rect 126426 152688 126482 152697
rect 126426 152623 126482 152632
rect 126242 152416 126298 152425
rect 126242 152351 126298 152360
rect 126256 150090 126284 152351
rect 126900 150090 126928 153886
rect 127084 153105 127112 159423
rect 127360 158846 127388 163200
rect 127808 158908 127860 158914
rect 127808 158850 127860 158856
rect 127348 158840 127400 158846
rect 127348 158782 127400 158788
rect 127532 156800 127584 156806
rect 127532 156742 127584 156748
rect 127070 153096 127126 153105
rect 127070 153031 127126 153040
rect 127544 150090 127572 156742
rect 127820 154018 127848 158850
rect 128188 156806 128216 163200
rect 128176 156800 128228 156806
rect 128176 156742 128228 156748
rect 129016 155242 129044 163200
rect 129004 155236 129056 155242
rect 129004 155178 129056 155184
rect 128360 154828 128412 154834
rect 128360 154770 128412 154776
rect 127808 154012 127860 154018
rect 127808 153954 127860 153960
rect 128372 152046 128400 154770
rect 129464 154080 129516 154086
rect 129464 154022 129516 154028
rect 129556 154080 129608 154086
rect 129556 154022 129608 154028
rect 128818 152552 128874 152561
rect 128818 152487 128874 152496
rect 128176 152040 128228 152046
rect 128176 151982 128228 151988
rect 128360 152040 128412 152046
rect 128360 151982 128412 151988
rect 128188 150090 128216 151982
rect 128832 150226 128860 152487
rect 129476 150226 129504 154022
rect 129568 153882 129596 154022
rect 129936 153882 129964 163200
rect 130764 158914 130792 163200
rect 130752 158908 130804 158914
rect 130752 158850 130804 158856
rect 130844 158840 130896 158846
rect 130844 158782 130896 158788
rect 130108 156732 130160 156738
rect 130108 156674 130160 156680
rect 129556 153876 129608 153882
rect 129556 153818 129608 153824
rect 129924 153876 129976 153882
rect 129924 153818 129976 153824
rect 130120 150226 130148 156674
rect 130856 152658 130884 158782
rect 131592 158030 131620 163200
rect 131580 158024 131632 158030
rect 131580 157966 131632 157972
rect 132420 156738 132448 163200
rect 133248 158846 133276 163200
rect 133236 158840 133288 158846
rect 133236 158782 133288 158788
rect 132500 156936 132552 156942
rect 132500 156878 132552 156884
rect 132408 156732 132460 156738
rect 132408 156674 132460 156680
rect 132038 153912 132094 153921
rect 132038 153847 132094 153856
rect 131394 153096 131450 153105
rect 131394 153031 131450 153040
rect 130752 152652 130804 152658
rect 130752 152594 130804 152600
rect 130844 152652 130896 152658
rect 130844 152594 130896 152600
rect 130764 150226 130792 152594
rect 131408 150226 131436 153031
rect 132052 150226 132080 153847
rect 132512 151814 132540 156878
rect 134076 155446 134104 163200
rect 134904 156942 134932 163200
rect 135168 159452 135220 159458
rect 135168 159394 135220 159400
rect 134892 156936 134944 156942
rect 134892 156878 134944 156884
rect 134064 155440 134116 155446
rect 134064 155382 134116 155388
rect 133328 154896 133380 154902
rect 133328 154838 133380 154844
rect 132512 151786 132724 151814
rect 132696 150226 132724 151786
rect 133340 150226 133368 154838
rect 134614 153776 134670 153785
rect 134614 153711 134670 153720
rect 133972 152584 134024 152590
rect 133972 152526 134024 152532
rect 133984 150226 134012 152526
rect 134628 150226 134656 153711
rect 135180 152590 135208 159394
rect 135442 159352 135498 159361
rect 135442 159287 135498 159296
rect 135260 156868 135312 156874
rect 135260 156810 135312 156816
rect 135168 152584 135220 152590
rect 135168 152526 135220 152532
rect 135272 150226 135300 156810
rect 128832 150198 128906 150226
rect 129476 150198 129550 150226
rect 130120 150198 130194 150226
rect 130764 150198 130838 150226
rect 131408 150198 131482 150226
rect 132052 150198 132126 150226
rect 132696 150198 132770 150226
rect 133340 150198 133414 150226
rect 133984 150198 134058 150226
rect 134628 150198 134702 150226
rect 135272 150198 135346 150226
rect 135456 150210 135484 159287
rect 135824 156874 135852 163200
rect 136652 159866 136680 163200
rect 136548 159860 136600 159866
rect 136548 159802 136600 159808
rect 136640 159860 136692 159866
rect 136640 159802 136692 159808
rect 136560 159458 136588 159802
rect 137480 159526 137508 163200
rect 137560 159724 137612 159730
rect 137560 159666 137612 159672
rect 137376 159520 137428 159526
rect 137374 159488 137376 159497
rect 137468 159520 137520 159526
rect 137428 159488 137430 159497
rect 136548 159452 136600 159458
rect 137468 159462 137520 159468
rect 137374 159423 137430 159432
rect 136548 159394 136600 159400
rect 137376 158840 137428 158846
rect 137204 158788 137376 158794
rect 137204 158782 137428 158788
rect 137204 158778 137416 158782
rect 137192 158772 137416 158778
rect 137244 158766 137416 158772
rect 137192 158714 137244 158720
rect 137192 157004 137244 157010
rect 137192 156946 137244 156952
rect 135812 156868 135864 156874
rect 135812 156810 135864 156816
rect 137100 154284 137152 154290
rect 137100 154226 137152 154232
rect 137008 154216 137060 154222
rect 137008 154158 137060 154164
rect 135904 152720 135956 152726
rect 135904 152662 135956 152668
rect 135916 150226 135944 152662
rect 137020 151814 137048 154158
rect 137112 153921 137140 154226
rect 137098 153912 137154 153921
rect 137098 153847 137154 153856
rect 137204 151814 137232 156946
rect 137468 155440 137520 155446
rect 137468 155382 137520 155388
rect 137480 152726 137508 155382
rect 137572 154086 137600 159666
rect 138018 159488 138074 159497
rect 138018 159423 138074 159432
rect 137560 154080 137612 154086
rect 137560 154022 137612 154028
rect 137652 154012 137704 154018
rect 137652 153954 137704 153960
rect 137664 153921 137692 153954
rect 137650 153912 137706 153921
rect 137650 153847 137706 153856
rect 137468 152720 137520 152726
rect 137468 152662 137520 152668
rect 138032 151842 138060 159423
rect 138308 156058 138336 163200
rect 139136 157010 139164 163200
rect 139964 159730 139992 163200
rect 139952 159724 140004 159730
rect 139952 159666 140004 159672
rect 139398 159624 139454 159633
rect 139398 159559 139454 159568
rect 139124 157004 139176 157010
rect 139124 156946 139176 156952
rect 138296 156052 138348 156058
rect 138296 155994 138348 156000
rect 139124 152788 139176 152794
rect 139124 152730 139176 152736
rect 138572 152584 138624 152590
rect 138572 152526 138624 152532
rect 138584 151910 138612 152526
rect 138480 151904 138532 151910
rect 138480 151846 138532 151852
rect 138572 151904 138624 151910
rect 138572 151846 138624 151852
rect 138020 151836 138072 151842
rect 137020 151786 137140 151814
rect 137204 151786 137876 151814
rect 137112 150226 137140 151786
rect 137848 150226 137876 151786
rect 138020 151778 138072 151784
rect 138492 150226 138520 151846
rect 139136 150226 139164 152730
rect 139412 152726 139440 159559
rect 139950 156768 140006 156777
rect 139950 156703 140006 156712
rect 139766 154048 139822 154057
rect 139766 153983 139822 153992
rect 139400 152720 139452 152726
rect 139400 152662 139452 152668
rect 139780 150226 139808 153983
rect 139964 151814 139992 156703
rect 140792 152590 140820 163200
rect 141712 157418 141740 163200
rect 141700 157412 141752 157418
rect 141700 157354 141752 157360
rect 142540 155446 142568 163200
rect 143368 159662 143396 163200
rect 143264 159656 143316 159662
rect 143264 159598 143316 159604
rect 143356 159656 143408 159662
rect 143356 159598 143408 159604
rect 142986 156632 143042 156641
rect 142986 156567 143042 156576
rect 142528 155440 142580 155446
rect 142528 155382 142580 155388
rect 142344 154012 142396 154018
rect 142344 153954 142396 153960
rect 141700 152720 141752 152726
rect 141700 152662 141752 152668
rect 141792 152720 141844 152726
rect 141792 152662 141844 152668
rect 140780 152584 140832 152590
rect 140780 152526 140832 152532
rect 141056 152448 141108 152454
rect 141056 152390 141108 152396
rect 139964 151786 140452 151814
rect 140424 150226 140452 151786
rect 141068 150226 141096 152390
rect 141712 150226 141740 152662
rect 141804 151842 141832 152662
rect 141792 151836 141844 151842
rect 141792 151778 141844 151784
rect 142356 150226 142384 153954
rect 143000 150226 143028 156567
rect 143276 151842 143304 159598
rect 144196 159458 144224 163200
rect 145024 163146 145052 163200
rect 145116 163146 145144 163254
rect 145024 163118 145144 163146
rect 144092 159452 144144 159458
rect 144092 159394 144144 159400
rect 144184 159452 144236 159458
rect 144184 159394 144236 159400
rect 143724 157140 143776 157146
rect 143724 157082 143776 157088
rect 143736 156602 143764 157082
rect 143724 156596 143776 156602
rect 143724 156538 143776 156544
rect 143552 152794 143764 152810
rect 143540 152788 143764 152794
rect 143592 152782 143764 152788
rect 143540 152730 143592 152736
rect 143736 152708 143764 152782
rect 143816 152720 143868 152726
rect 143630 152688 143686 152697
rect 143736 152680 143816 152708
rect 143816 152662 143868 152668
rect 143630 152623 143686 152632
rect 143264 151836 143316 151842
rect 143264 151778 143316 151784
rect 143644 150226 143672 152623
rect 144104 152454 144132 159394
rect 144918 157992 144974 158001
rect 144918 157927 144974 157936
rect 144092 152448 144144 152454
rect 144092 152390 144144 152396
rect 144276 152380 144328 152386
rect 144276 152322 144328 152328
rect 144288 150226 144316 152322
rect 144932 150226 144960 157927
rect 145300 157078 145328 163254
rect 145838 163200 145894 164400
rect 146666 163200 146722 164400
rect 146772 163254 147076 163282
rect 145472 157140 145524 157146
rect 145472 157082 145524 157088
rect 145288 157072 145340 157078
rect 145288 157014 145340 157020
rect 145380 154420 145432 154426
rect 145380 154362 145432 154368
rect 145104 154352 145156 154358
rect 145104 154294 145156 154300
rect 145116 154018 145144 154294
rect 145104 154012 145156 154018
rect 145104 153954 145156 153960
rect 145392 150498 145420 154362
rect 145484 151814 145512 157082
rect 145852 154902 145880 163200
rect 146680 163146 146708 163200
rect 146772 163146 146800 163254
rect 146680 163118 146800 163146
rect 147048 159866 147076 163254
rect 147586 163200 147642 164400
rect 148414 163200 148470 164400
rect 149242 163200 149298 164400
rect 150070 163200 150126 164400
rect 150176 163254 150388 163282
rect 147036 159860 147088 159866
rect 147036 159802 147088 159808
rect 146852 159792 146904 159798
rect 147312 159792 147364 159798
rect 146904 159740 147260 159746
rect 146852 159734 147260 159740
rect 147312 159734 147364 159740
rect 146864 159718 147260 159734
rect 146668 159656 146720 159662
rect 146944 159656 146996 159662
rect 146720 159604 146944 159610
rect 146668 159598 146996 159604
rect 146208 159588 146260 159594
rect 146680 159582 146984 159598
rect 146208 159530 146260 159536
rect 145840 154896 145892 154902
rect 145840 154838 145892 154844
rect 146220 154698 146248 159530
rect 146760 159520 146812 159526
rect 146812 159468 146984 159474
rect 146760 159462 146984 159468
rect 146772 159446 146984 159462
rect 147232 159458 147260 159718
rect 146956 159390 146984 159446
rect 147220 159452 147272 159458
rect 147220 159394 147272 159400
rect 146852 159384 146904 159390
rect 146852 159326 146904 159332
rect 146944 159384 146996 159390
rect 146944 159326 146996 159332
rect 146864 158658 146892 159326
rect 147324 158846 147352 159734
rect 147600 158846 147628 163200
rect 147312 158840 147364 158846
rect 147312 158782 147364 158788
rect 147588 158840 147640 158846
rect 147588 158782 147640 158788
rect 146864 158630 147168 158658
rect 146392 158092 146444 158098
rect 146392 158034 146444 158040
rect 146208 154692 146260 154698
rect 146208 154634 146260 154640
rect 145484 151786 146248 151814
rect 145392 150470 145604 150498
rect 145576 150226 145604 150470
rect 146220 150226 146248 151786
rect 124324 150062 124398 150090
rect 124968 150062 125042 150090
rect 125612 150062 125686 150090
rect 126256 150062 126330 150090
rect 126900 150062 126974 150090
rect 127544 150062 127618 150090
rect 128188 150062 128262 150090
rect 124370 149940 124398 150062
rect 125014 149940 125042 150062
rect 125658 149940 125686 150062
rect 126302 149940 126330 150062
rect 126946 149940 126974 150062
rect 127590 149940 127618 150062
rect 128234 149940 128262 150062
rect 128878 149940 128906 150198
rect 129522 149940 129550 150198
rect 130166 149940 130194 150198
rect 130810 149940 130838 150198
rect 131454 149940 131482 150198
rect 132098 149940 132126 150198
rect 132742 149940 132770 150198
rect 133386 149940 133414 150198
rect 134030 149940 134058 150198
rect 134674 149940 134702 150198
rect 135318 149940 135346 150198
rect 135444 150204 135496 150210
rect 135916 150198 135990 150226
rect 135444 150146 135496 150152
rect 135962 149940 135990 150198
rect 136594 150204 136646 150210
rect 137112 150198 137278 150226
rect 137848 150198 137922 150226
rect 138492 150198 138566 150226
rect 139136 150198 139210 150226
rect 139780 150198 139854 150226
rect 140424 150198 140498 150226
rect 141068 150198 141142 150226
rect 141712 150198 141786 150226
rect 142356 150198 142430 150226
rect 143000 150198 143074 150226
rect 143644 150198 143718 150226
rect 144288 150198 144362 150226
rect 144932 150198 145006 150226
rect 145576 150198 145650 150226
rect 146220 150198 146294 150226
rect 146404 150210 146432 158034
rect 146484 154556 146536 154562
rect 146484 154498 146536 154504
rect 146496 154442 146524 154498
rect 146496 154414 147076 154442
rect 146944 154352 146996 154358
rect 146944 154294 146996 154300
rect 146956 154170 146984 154294
rect 146864 154154 146984 154170
rect 147048 154154 147076 154414
rect 147140 154222 147168 158630
rect 148428 158098 148456 163200
rect 148784 159928 148836 159934
rect 148784 159870 148836 159876
rect 148876 159928 148928 159934
rect 148876 159870 148928 159876
rect 149256 159882 149284 163200
rect 150084 163146 150112 163200
rect 150176 163146 150204 163254
rect 150084 163118 150204 163146
rect 148796 158930 148824 159870
rect 148888 159798 148916 159870
rect 149256 159854 149468 159882
rect 148876 159792 148928 159798
rect 148876 159734 148928 159740
rect 149336 159724 149388 159730
rect 149336 159666 149388 159672
rect 149060 159656 149112 159662
rect 149348 159610 149376 159666
rect 149112 159604 149376 159610
rect 149060 159598 149376 159604
rect 149072 159582 149376 159598
rect 148796 158902 149192 158930
rect 149164 158846 149192 158902
rect 149060 158840 149112 158846
rect 149060 158782 149112 158788
rect 149152 158840 149204 158846
rect 149152 158782 149204 158788
rect 148416 158092 148468 158098
rect 148416 158034 148468 158040
rect 147680 156596 147732 156602
rect 147680 156538 147732 156544
rect 147128 154216 147180 154222
rect 147128 154158 147180 154164
rect 146852 154148 146984 154154
rect 146904 154142 146984 154148
rect 147036 154148 147088 154154
rect 146852 154090 146904 154096
rect 147036 154090 147088 154096
rect 146852 151904 146904 151910
rect 146852 151846 146904 151852
rect 146864 150226 146892 151846
rect 136594 150146 136646 150152
rect 136606 149940 136634 150146
rect 137250 149940 137278 150198
rect 137894 149940 137922 150198
rect 138538 149940 138566 150198
rect 139182 149940 139210 150198
rect 139826 149940 139854 150198
rect 140470 149940 140498 150198
rect 141114 149940 141142 150198
rect 141758 149940 141786 150198
rect 142402 149940 142430 150198
rect 143046 149940 143074 150198
rect 143690 149940 143718 150198
rect 144334 149940 144362 150198
rect 144978 149940 145006 150198
rect 145622 149940 145650 150198
rect 146266 149940 146294 150198
rect 146392 150204 146444 150210
rect 146864 150198 146938 150226
rect 147692 150210 147720 156538
rect 148140 154012 148192 154018
rect 148140 153954 148192 153960
rect 148152 150226 148180 153954
rect 149072 152454 149100 158782
rect 149440 157334 149468 159854
rect 149610 158264 149666 158273
rect 149610 158199 149666 158208
rect 149256 157306 149468 157334
rect 149256 154834 149284 157306
rect 149244 154828 149296 154834
rect 149244 154770 149296 154776
rect 149060 152448 149112 152454
rect 149060 152390 149112 152396
rect 149428 152108 149480 152114
rect 149428 152050 149480 152056
rect 149440 150226 149468 152050
rect 149624 151814 149652 158199
rect 150360 154018 150388 163254
rect 150898 163200 150954 164400
rect 151726 163200 151782 164400
rect 152554 163200 152610 164400
rect 153474 163200 153530 164400
rect 154302 163200 154358 164400
rect 155130 163200 155186 164400
rect 155958 163200 156014 164400
rect 156786 163200 156842 164400
rect 157614 163200 157670 164400
rect 158442 163200 158498 164400
rect 159362 163200 159418 164400
rect 160190 163200 160246 164400
rect 161018 163200 161074 164400
rect 161846 163200 161902 164400
rect 162674 163200 162730 164400
rect 163502 163200 163558 164400
rect 164330 163200 164386 164400
rect 165250 163200 165306 164400
rect 166078 163200 166134 164400
rect 166184 163254 166396 163282
rect 150544 159866 150756 159882
rect 150532 159860 150768 159866
rect 150584 159854 150716 159860
rect 150532 159802 150584 159808
rect 150716 159802 150768 159808
rect 150912 159458 150940 163200
rect 150440 159452 150492 159458
rect 150440 159394 150492 159400
rect 150900 159452 150952 159458
rect 150900 159394 150952 159400
rect 150348 154012 150400 154018
rect 150348 153954 150400 153960
rect 150452 152114 150480 159394
rect 151740 157146 151768 163200
rect 152568 160290 152596 163200
rect 152568 160262 152688 160290
rect 152464 159928 152516 159934
rect 152464 159870 152516 159876
rect 152476 159322 152504 159870
rect 152464 159316 152516 159322
rect 152464 159258 152516 159264
rect 152554 158128 152610 158137
rect 152554 158063 152610 158072
rect 151728 157140 151780 157146
rect 151728 157082 151780 157088
rect 150714 156904 150770 156913
rect 150714 156839 150770 156848
rect 150624 154556 150676 154562
rect 150624 154498 150676 154504
rect 150440 152108 150492 152114
rect 150440 152050 150492 152056
rect 149624 151786 150020 151814
rect 149992 150226 150020 151786
rect 150636 150226 150664 154498
rect 150728 151814 150756 156839
rect 151912 152788 151964 152794
rect 151912 152730 151964 152736
rect 150728 151786 151308 151814
rect 151280 150226 151308 151786
rect 151924 150226 151952 152730
rect 152568 150226 152596 158063
rect 152660 154086 152688 160262
rect 153488 159798 153516 163200
rect 153384 159792 153436 159798
rect 153384 159734 153436 159740
rect 153476 159792 153528 159798
rect 153476 159734 153528 159740
rect 153396 154154 153424 159734
rect 153752 157208 153804 157214
rect 153752 157150 153804 157156
rect 153200 154148 153252 154154
rect 153200 154090 153252 154096
rect 153384 154148 153436 154154
rect 153384 154090 153436 154096
rect 152648 154080 152700 154086
rect 152648 154022 152700 154028
rect 153212 150226 153240 154090
rect 153764 151814 153792 157150
rect 154316 152794 154344 163200
rect 155144 158166 155172 163200
rect 155040 158160 155092 158166
rect 155040 158102 155092 158108
rect 155132 158160 155184 158166
rect 155132 158102 155184 158108
rect 154304 152788 154356 152794
rect 154304 152730 154356 152736
rect 154488 152176 154540 152182
rect 154488 152118 154540 152124
rect 153764 151786 153884 151814
rect 153856 150226 153884 151786
rect 154500 150226 154528 152118
rect 155052 151814 155080 158102
rect 155972 154766 156000 163200
rect 156800 158846 156828 163200
rect 157154 159624 157210 159633
rect 157154 159559 157156 159568
rect 157208 159559 157210 159568
rect 157338 159624 157394 159633
rect 157628 159594 157656 163200
rect 157338 159559 157394 159568
rect 157616 159588 157668 159594
rect 157156 159530 157208 159536
rect 156052 158840 156104 158846
rect 156052 158782 156104 158788
rect 156788 158840 156840 158846
rect 156788 158782 156840 158788
rect 155960 154760 156012 154766
rect 155960 154702 156012 154708
rect 155776 153808 155828 153814
rect 155776 153750 155828 153756
rect 155052 151786 155172 151814
rect 155144 150226 155172 151786
rect 155788 150226 155816 153750
rect 156064 152182 156092 158782
rect 156418 157040 156474 157049
rect 156418 156975 156474 156984
rect 156052 152176 156104 152182
rect 156052 152118 156104 152124
rect 156432 150226 156460 156975
rect 157352 154562 157380 159559
rect 157616 159530 157668 159536
rect 158456 158234 158484 163200
rect 158720 158772 158772 158778
rect 158720 158714 158772 158720
rect 157708 158228 157760 158234
rect 157708 158170 157760 158176
rect 158444 158228 158496 158234
rect 158444 158170 158496 158176
rect 156788 154556 156840 154562
rect 156788 154498 156840 154504
rect 157340 154556 157392 154562
rect 157340 154498 157392 154504
rect 156604 154216 156656 154222
rect 156604 154158 156656 154164
rect 156696 154216 156748 154222
rect 156696 154158 156748 154164
rect 156616 153814 156644 154158
rect 156604 153808 156656 153814
rect 156604 153750 156656 153756
rect 156708 153746 156736 154158
rect 156800 153746 156828 154498
rect 156696 153740 156748 153746
rect 156696 153682 156748 153688
rect 156788 153740 156840 153746
rect 156788 153682 156840 153688
rect 157064 151904 157116 151910
rect 157064 151846 157116 151852
rect 157076 150226 157104 151846
rect 157720 150226 157748 158170
rect 158732 156602 158760 158714
rect 158996 157276 159048 157282
rect 158996 157218 159048 157224
rect 158720 156596 158772 156602
rect 158720 156538 158772 156544
rect 158350 154184 158406 154193
rect 158350 154119 158406 154128
rect 158364 150226 158392 154119
rect 159008 150226 159036 157218
rect 159376 154630 159404 163200
rect 160204 159934 160232 163200
rect 160100 159928 160152 159934
rect 160100 159870 160152 159876
rect 160192 159928 160244 159934
rect 160192 159870 160244 159876
rect 160112 159746 160140 159870
rect 160112 159718 160232 159746
rect 160100 159656 160152 159662
rect 160100 159598 160152 159604
rect 160112 157282 160140 159598
rect 160100 157276 160152 157282
rect 160100 157218 160152 157224
rect 159364 154624 159416 154630
rect 159364 154566 159416 154572
rect 159640 152312 159692 152318
rect 159640 152254 159692 152260
rect 159652 150226 159680 152254
rect 160204 151910 160232 159718
rect 161032 159662 161060 163200
rect 161020 159656 161072 159662
rect 161020 159598 161072 159604
rect 161860 158302 161888 163200
rect 160284 158296 160336 158302
rect 160284 158238 160336 158244
rect 161848 158296 161900 158302
rect 161848 158238 161900 158244
rect 160192 151904 160244 151910
rect 160192 151846 160244 151852
rect 160296 150226 160324 158238
rect 161572 157344 161624 157350
rect 161572 157286 161624 157292
rect 160926 154320 160982 154329
rect 160926 154255 160982 154264
rect 160940 150226 160968 154255
rect 161584 150226 161612 157286
rect 162688 154698 162716 163200
rect 163516 159322 163544 163200
rect 164344 161474 164372 163200
rect 164344 161446 164464 161474
rect 164148 159724 164200 159730
rect 164148 159666 164200 159672
rect 163504 159316 163556 159322
rect 163504 159258 163556 159264
rect 162858 158400 162914 158409
rect 162858 158335 162914 158344
rect 162676 154692 162728 154698
rect 162676 154634 162728 154640
rect 162216 152380 162268 152386
rect 162216 152322 162268 152328
rect 162228 150226 162256 152322
rect 162872 150226 162900 158335
rect 164160 156074 164188 159666
rect 164332 158364 164384 158370
rect 164332 158306 164384 158312
rect 164160 156046 164280 156074
rect 164252 155990 164280 156046
rect 164148 155984 164200 155990
rect 164148 155926 164200 155932
rect 164240 155984 164292 155990
rect 164240 155926 164292 155932
rect 163504 154216 163556 154222
rect 163504 154158 163556 154164
rect 163516 150226 163544 154158
rect 164160 150226 164188 155926
rect 146392 150146 146444 150152
rect 146910 149940 146938 150198
rect 147542 150204 147594 150210
rect 147542 150146 147594 150152
rect 147680 150204 147732 150210
rect 148152 150198 148226 150226
rect 147680 150146 147732 150152
rect 147554 149940 147582 150146
rect 148198 149940 148226 150198
rect 148830 150204 148882 150210
rect 149440 150198 149514 150226
rect 149992 150198 150066 150226
rect 150636 150198 150710 150226
rect 151280 150198 151354 150226
rect 151924 150198 151998 150226
rect 152568 150198 152642 150226
rect 153212 150198 153286 150226
rect 153856 150198 153930 150226
rect 154500 150198 154574 150226
rect 155144 150198 155218 150226
rect 155788 150198 155862 150226
rect 156432 150198 156506 150226
rect 157076 150198 157150 150226
rect 157720 150198 157794 150226
rect 158364 150198 158438 150226
rect 159008 150198 159082 150226
rect 159652 150198 159726 150226
rect 160296 150198 160370 150226
rect 160940 150198 161014 150226
rect 161584 150198 161658 150226
rect 162228 150198 162302 150226
rect 162872 150198 162946 150226
rect 163516 150198 163590 150226
rect 164160 150198 164234 150226
rect 164344 150210 164372 158306
rect 164436 152386 164464 161446
rect 165264 158370 165292 163200
rect 166092 163146 166120 163200
rect 166184 163146 166212 163254
rect 166092 163118 166212 163146
rect 165252 158364 165304 158370
rect 165252 158306 165304 158312
rect 165620 155508 165672 155514
rect 165620 155450 165672 155456
rect 165068 154216 165120 154222
rect 165068 154158 165120 154164
rect 165080 153678 165108 154158
rect 165068 153672 165120 153678
rect 165068 153614 165120 153620
rect 164424 152380 164476 152386
rect 164424 152322 164476 152328
rect 164792 152244 164844 152250
rect 164792 152186 164844 152192
rect 164804 150226 164832 152186
rect 148830 150146 148882 150152
rect 148842 149940 148870 150146
rect 149486 149940 149514 150198
rect 150038 149940 150066 150198
rect 150682 149940 150710 150198
rect 151326 149940 151354 150198
rect 151970 149940 151998 150198
rect 152614 149940 152642 150198
rect 153258 149940 153286 150198
rect 153902 149940 153930 150198
rect 154546 149940 154574 150198
rect 155190 149940 155218 150198
rect 155834 149940 155862 150198
rect 156478 149940 156506 150198
rect 157122 149940 157150 150198
rect 157766 149940 157794 150198
rect 158410 149940 158438 150198
rect 159054 149940 159082 150198
rect 159698 149940 159726 150198
rect 160342 149940 160370 150198
rect 160986 149940 161014 150198
rect 161630 149940 161658 150198
rect 162274 149940 162302 150198
rect 162918 149940 162946 150198
rect 163562 149940 163590 150198
rect 164206 149940 164234 150198
rect 164332 150204 164384 150210
rect 164804 150198 164878 150226
rect 165632 150210 165660 155450
rect 166078 155272 166134 155281
rect 166078 155207 166134 155216
rect 166092 150226 166120 155207
rect 166368 154154 166396 163254
rect 166906 163200 166962 164400
rect 167734 163200 167790 164400
rect 168562 163200 168618 164400
rect 169390 163200 169446 164400
rect 170218 163200 170274 164400
rect 171138 163200 171194 164400
rect 171966 163200 172022 164400
rect 172794 163200 172850 164400
rect 173622 163200 173678 164400
rect 174450 163200 174506 164400
rect 175278 163200 175334 164400
rect 176106 163200 176162 164400
rect 177026 163200 177082 164400
rect 177854 163200 177910 164400
rect 178682 163200 178738 164400
rect 179510 163200 179566 164400
rect 180338 163200 180394 164400
rect 181166 163200 181222 164400
rect 181994 163200 182050 164400
rect 182914 163200 182970 164400
rect 183742 163200 183798 164400
rect 184570 163200 184626 164400
rect 185398 163200 185454 164400
rect 186226 163200 186282 164400
rect 187054 163200 187110 164400
rect 187882 163200 187938 164400
rect 188802 163200 188858 164400
rect 189630 163200 189686 164400
rect 190458 163200 190514 164400
rect 191286 163200 191342 164400
rect 192114 163200 192170 164400
rect 192942 163200 192998 164400
rect 193770 163200 193826 164400
rect 194690 163200 194746 164400
rect 195518 163200 195574 164400
rect 196346 163200 196402 164400
rect 197174 163200 197230 164400
rect 198002 163200 198058 164400
rect 198830 163200 198886 164400
rect 199658 163200 199714 164400
rect 200578 163200 200634 164400
rect 201406 163200 201462 164400
rect 202234 163200 202290 164400
rect 203062 163200 203118 164400
rect 203890 163200 203946 164400
rect 204718 163200 204774 164400
rect 205546 163200 205602 164400
rect 206466 163200 206522 164400
rect 207294 163200 207350 164400
rect 208122 163200 208178 164400
rect 208950 163200 209006 164400
rect 209778 163200 209834 164400
rect 210606 163200 210662 164400
rect 211434 163200 211490 164400
rect 212354 163200 212410 164400
rect 213182 163200 213238 164400
rect 214010 163200 214066 164400
rect 214838 163200 214894 164400
rect 215666 163200 215722 164400
rect 216494 163200 216550 164400
rect 217322 163200 217378 164400
rect 218242 163200 218298 164400
rect 219070 163200 219126 164400
rect 219176 163254 219388 163282
rect 166920 157214 166948 163200
rect 167000 160064 167052 160070
rect 167000 160006 167052 160012
rect 166908 157208 166960 157214
rect 166908 157150 166960 157156
rect 166264 154148 166316 154154
rect 166264 154090 166316 154096
rect 166356 154148 166408 154154
rect 166356 154090 166408 154096
rect 166276 153678 166304 154090
rect 166264 153672 166316 153678
rect 166264 153614 166316 153620
rect 167012 152250 167040 160006
rect 167748 159730 167776 163200
rect 167736 159724 167788 159730
rect 167736 159666 167788 159672
rect 168576 158438 168604 163200
rect 167552 158432 167604 158438
rect 167552 158374 167604 158380
rect 168564 158432 168616 158438
rect 168564 158374 168616 158380
rect 167000 152244 167052 152250
rect 167000 152186 167052 152192
rect 167368 152108 167420 152114
rect 167368 152050 167420 152056
rect 167380 150226 167408 152050
rect 167564 151814 167592 158374
rect 169298 157176 169354 157185
rect 169298 157111 169354 157120
rect 168656 154216 168708 154222
rect 168656 154158 168708 154164
rect 167564 151786 168052 151814
rect 168024 150226 168052 151786
rect 168668 150226 168696 154158
rect 169312 150226 169340 157111
rect 169404 155514 169432 163200
rect 170232 160070 170260 163200
rect 170220 160064 170272 160070
rect 170220 160006 170272 160012
rect 169760 159180 169812 159186
rect 169760 159122 169812 159128
rect 169392 155508 169444 155514
rect 169392 155450 169444 155456
rect 169772 152114 169800 159122
rect 171152 158778 171180 163200
rect 171140 158772 171192 158778
rect 171140 158714 171192 158720
rect 171980 158642 172008 163200
rect 172612 158772 172664 158778
rect 172612 158714 172664 158720
rect 170312 158636 170364 158642
rect 170312 158578 170364 158584
rect 171968 158636 172020 158642
rect 171968 158578 172020 158584
rect 169944 152856 169996 152862
rect 169944 152798 169996 152804
rect 169760 152108 169812 152114
rect 169760 152050 169812 152056
rect 169956 150226 169984 152798
rect 170324 151814 170352 158578
rect 171138 155544 171194 155553
rect 171138 155479 171194 155488
rect 170324 151786 170628 151814
rect 170600 150226 170628 151786
rect 164332 150146 164384 150152
rect 164850 149940 164878 150198
rect 165482 150204 165534 150210
rect 165482 150146 165534 150152
rect 165620 150204 165672 150210
rect 166092 150198 166166 150226
rect 165620 150146 165672 150152
rect 165494 149940 165522 150146
rect 166138 149940 166166 150198
rect 166770 150204 166822 150210
rect 167380 150198 167454 150226
rect 168024 150198 168098 150226
rect 168668 150198 168742 150226
rect 169312 150198 169386 150226
rect 169956 150198 170030 150226
rect 170600 150198 170674 150226
rect 171152 150210 171180 155479
rect 171230 155408 171286 155417
rect 171230 155343 171286 155352
rect 171244 150226 171272 155343
rect 172624 152318 172652 158714
rect 172704 158568 172756 158574
rect 172704 158510 172756 158516
rect 172612 152312 172664 152318
rect 172612 152254 172664 152260
rect 172520 152176 172572 152182
rect 172520 152118 172572 152124
rect 172532 150226 172560 152118
rect 172716 151814 172744 158510
rect 172808 154222 172836 163200
rect 173636 158778 173664 163200
rect 174464 161474 174492 163200
rect 174464 161446 174584 161474
rect 173624 158772 173676 158778
rect 173624 158714 173676 158720
rect 174452 156528 174504 156534
rect 174452 156470 174504 156476
rect 173072 155712 173124 155718
rect 173072 155654 173124 155660
rect 172796 154216 172848 154222
rect 172796 154158 172848 154164
rect 173084 151814 173112 155654
rect 172716 151786 173020 151814
rect 173084 151786 173848 151814
rect 172992 150498 173020 151786
rect 172992 150470 173204 150498
rect 173176 150226 173204 150470
rect 173820 150226 173848 151786
rect 174464 150226 174492 156470
rect 174556 152862 174584 161446
rect 174636 159860 174688 159866
rect 174636 159802 174688 159808
rect 174648 156534 174676 159802
rect 175292 158506 175320 163200
rect 176120 161474 176148 163200
rect 176120 161446 176332 161474
rect 175188 158500 175240 158506
rect 175188 158442 175240 158448
rect 175280 158500 175332 158506
rect 175280 158442 175332 158448
rect 175200 158386 175228 158442
rect 175200 158358 175320 158386
rect 174636 156528 174688 156534
rect 174636 156470 174688 156476
rect 174544 152856 174596 152862
rect 174544 152798 174596 152804
rect 175096 151972 175148 151978
rect 175096 151914 175148 151920
rect 175108 150226 175136 151914
rect 175292 151814 175320 158358
rect 176200 157956 176252 157962
rect 176200 157898 176252 157904
rect 175924 157888 175976 157894
rect 176212 157842 176240 157898
rect 175976 157836 176240 157842
rect 175924 157830 176240 157836
rect 175936 157814 176240 157830
rect 176304 155718 176332 161446
rect 176660 159180 176712 159186
rect 176660 159122 176712 159128
rect 176292 155712 176344 155718
rect 176292 155654 176344 155660
rect 176384 155644 176436 155650
rect 176384 155586 176436 155592
rect 175292 151786 175780 151814
rect 175752 150226 175780 151786
rect 176396 150226 176424 155586
rect 176672 152182 176700 159122
rect 177040 157334 177068 163200
rect 177868 159798 177896 163200
rect 177856 159792 177908 159798
rect 177856 159734 177908 159740
rect 178696 158574 178724 163200
rect 178684 158568 178736 158574
rect 178684 158510 178736 158516
rect 178040 157888 178092 157894
rect 178040 157830 178092 157836
rect 177040 157306 177160 157334
rect 177132 155718 177160 157306
rect 177120 155712 177172 155718
rect 177026 155680 177082 155689
rect 177120 155654 177172 155660
rect 177026 155615 177082 155624
rect 176660 152176 176712 152182
rect 176660 152118 176712 152124
rect 177040 150226 177068 155615
rect 177672 151904 177724 151910
rect 177672 151846 177724 151852
rect 177684 150226 177712 151846
rect 178052 151814 178080 157830
rect 179524 155582 179552 163200
rect 180352 159254 180380 163200
rect 180708 159860 180760 159866
rect 180708 159802 180760 159808
rect 180340 159248 180392 159254
rect 180340 159190 180392 159196
rect 180720 158794 180748 159802
rect 180720 158766 180932 158794
rect 180904 158710 180932 158766
rect 180800 158704 180852 158710
rect 180800 158646 180852 158652
rect 180892 158704 180944 158710
rect 180892 158646 180944 158652
rect 179604 156460 179656 156466
rect 179604 156402 179656 156408
rect 178960 155576 179012 155582
rect 178960 155518 179012 155524
rect 179512 155576 179564 155582
rect 179512 155518 179564 155524
rect 178052 151786 178356 151814
rect 178328 150226 178356 151786
rect 178972 150226 179000 155518
rect 179616 150226 179644 156402
rect 180248 153060 180300 153066
rect 180248 153002 180300 153008
rect 180260 150226 180288 153002
rect 180812 150226 180840 158646
rect 181180 153066 181208 163200
rect 181444 159180 181496 159186
rect 181444 159122 181496 159128
rect 181456 158982 181484 159122
rect 181444 158976 181496 158982
rect 181444 158918 181496 158924
rect 182008 158710 182036 163200
rect 181904 158704 181956 158710
rect 181904 158646 181956 158652
rect 181996 158704 182048 158710
rect 181996 158646 182048 158652
rect 181272 157950 181576 157978
rect 181272 157758 181300 157950
rect 181548 157894 181576 157950
rect 181536 157888 181588 157894
rect 181536 157830 181588 157836
rect 181628 157820 181680 157826
rect 181628 157762 181680 157768
rect 181812 157820 181864 157826
rect 181812 157762 181864 157768
rect 181260 157752 181312 157758
rect 181260 157694 181312 157700
rect 181640 157706 181668 157762
rect 181640 157690 181760 157706
rect 181536 157684 181588 157690
rect 181640 157684 181772 157690
rect 181640 157678 181720 157684
rect 181536 157626 181588 157632
rect 181720 157626 181772 157632
rect 181548 157570 181576 157626
rect 181824 157570 181852 157762
rect 181916 157758 181944 158646
rect 182272 157956 182324 157962
rect 182272 157898 182324 157904
rect 181904 157752 181956 157758
rect 181904 157694 181956 157700
rect 181548 157542 181852 157570
rect 181444 155780 181496 155786
rect 181444 155722 181496 155728
rect 181168 153060 181220 153066
rect 181168 153002 181220 153008
rect 181456 150226 181484 155722
rect 182088 153604 182140 153610
rect 182088 153546 182140 153552
rect 182100 150226 182128 153546
rect 166770 150146 166822 150152
rect 166782 149940 166810 150146
rect 167426 149940 167454 150198
rect 168070 149940 168098 150198
rect 168714 149940 168742 150198
rect 169358 149940 169386 150198
rect 170002 149940 170030 150198
rect 170646 149940 170674 150198
rect 171140 150204 171192 150210
rect 171244 150198 171318 150226
rect 171140 150146 171192 150152
rect 171290 149940 171318 150198
rect 171922 150204 171974 150210
rect 172532 150198 172606 150226
rect 173176 150198 173250 150226
rect 173820 150198 173894 150226
rect 174464 150198 174538 150226
rect 175108 150198 175182 150226
rect 175752 150198 175826 150226
rect 176396 150198 176470 150226
rect 177040 150198 177114 150226
rect 177684 150198 177758 150226
rect 178328 150198 178402 150226
rect 178972 150198 179046 150226
rect 179616 150198 179690 150226
rect 180260 150198 180334 150226
rect 180812 150198 180886 150226
rect 181456 150198 181530 150226
rect 182100 150198 182174 150226
rect 182284 150210 182312 157898
rect 182928 153610 182956 163200
rect 183560 159248 183612 159254
rect 183612 159208 183692 159236
rect 183560 159190 183612 159196
rect 183100 159112 183152 159118
rect 183100 159054 183152 159060
rect 182916 153604 182968 153610
rect 182916 153546 182968 153552
rect 183112 152250 183140 159054
rect 183664 159050 183692 159208
rect 183756 159118 183784 163200
rect 184584 159866 184612 163200
rect 184572 159860 184624 159866
rect 184572 159802 184624 159808
rect 183744 159112 183796 159118
rect 183744 159054 183796 159060
rect 183652 159044 183704 159050
rect 183652 158986 183704 158992
rect 185412 157962 185440 163200
rect 185584 158976 185636 158982
rect 185584 158918 185636 158924
rect 185400 157956 185452 157962
rect 185400 157898 185452 157904
rect 185400 157684 185452 157690
rect 185400 157626 185452 157632
rect 184018 155816 184074 155825
rect 184018 155751 184074 155760
rect 183560 155168 183612 155174
rect 183560 155110 183612 155116
rect 182732 152244 182784 152250
rect 182732 152186 182784 152192
rect 183100 152244 183152 152250
rect 183100 152186 183152 152192
rect 182744 150226 182772 152186
rect 171922 150146 171974 150152
rect 171934 149940 171962 150146
rect 172578 149940 172606 150198
rect 173222 149940 173250 150198
rect 173866 149940 173894 150198
rect 174510 149940 174538 150198
rect 175154 149940 175182 150198
rect 175798 149940 175826 150198
rect 176442 149940 176470 150198
rect 177086 149940 177114 150198
rect 177730 149940 177758 150198
rect 178374 149940 178402 150198
rect 179018 149940 179046 150198
rect 179662 149940 179690 150198
rect 180306 149940 180334 150198
rect 180858 149940 180886 150198
rect 181502 149940 181530 150198
rect 182146 149940 182174 150198
rect 182272 150204 182324 150210
rect 182744 150198 182818 150226
rect 183572 150210 183600 155110
rect 184032 150226 184060 155751
rect 185124 154488 185176 154494
rect 185124 154430 185176 154436
rect 185136 153610 185164 154430
rect 185214 154320 185270 154329
rect 185214 154255 185216 154264
rect 185268 154255 185270 154264
rect 185308 154284 185360 154290
rect 185216 154226 185268 154232
rect 185308 154226 185360 154232
rect 185320 153626 185348 154226
rect 185032 153604 185084 153610
rect 185032 153546 185084 153552
rect 185124 153604 185176 153610
rect 185124 153546 185176 153552
rect 185228 153598 185348 153626
rect 185044 153490 185072 153546
rect 185228 153490 185256 153598
rect 185044 153462 185256 153490
rect 185308 152108 185360 152114
rect 185308 152050 185360 152056
rect 185320 150226 185348 152050
rect 185412 151814 185440 157626
rect 185596 151978 185624 158918
rect 186240 155786 186268 163200
rect 187068 159254 187096 163200
rect 187896 161474 187924 163200
rect 187896 161446 188016 161474
rect 187056 159248 187108 159254
rect 187056 159190 187108 159196
rect 186780 155916 186832 155922
rect 186780 155858 186832 155864
rect 186228 155780 186280 155786
rect 186228 155722 186280 155728
rect 186688 155168 186740 155174
rect 186688 155110 186740 155116
rect 186320 155100 186372 155106
rect 186504 155100 186556 155106
rect 186372 155060 186504 155088
rect 186320 155042 186372 155048
rect 186504 155042 186556 155048
rect 186228 155032 186280 155038
rect 186226 155000 186228 155009
rect 186596 155032 186648 155038
rect 186280 155000 186282 155009
rect 186594 155000 186596 155009
rect 186648 155000 186650 155009
rect 186226 154935 186282 154944
rect 186320 154964 186372 154970
rect 186594 154935 186650 154944
rect 186320 154906 186372 154912
rect 186332 154850 186360 154906
rect 186700 154850 186728 155110
rect 186332 154822 186728 154850
rect 185584 151972 185636 151978
rect 185584 151914 185636 151920
rect 185412 151786 185992 151814
rect 185964 150226 185992 151786
rect 186792 150226 186820 155858
rect 187238 154456 187294 154465
rect 187238 154391 187294 154400
rect 182272 150146 182324 150152
rect 182790 149940 182818 150198
rect 183422 150204 183474 150210
rect 183422 150146 183474 150152
rect 183560 150204 183612 150210
rect 184032 150198 184106 150226
rect 183560 150146 183612 150152
rect 183434 149940 183462 150146
rect 184078 149940 184106 150198
rect 184710 150204 184762 150210
rect 185320 150198 185394 150226
rect 185964 150198 186038 150226
rect 184710 150146 184762 150152
rect 184722 149940 184750 150146
rect 185366 149940 185394 150198
rect 186010 149940 186038 150198
rect 186654 150198 186820 150226
rect 186654 149940 186682 150198
rect 187252 150090 187280 154391
rect 187988 152930 188016 161446
rect 188344 159928 188396 159934
rect 188344 159870 188396 159876
rect 188356 154970 188384 159870
rect 188816 157894 188844 163200
rect 188528 157888 188580 157894
rect 188528 157830 188580 157836
rect 188804 157888 188856 157894
rect 188804 157830 188856 157836
rect 188344 154964 188396 154970
rect 188344 154906 188396 154912
rect 188436 154420 188488 154426
rect 188436 154362 188488 154368
rect 188448 153610 188476 154362
rect 188344 153604 188396 153610
rect 188344 153546 188396 153552
rect 188436 153604 188488 153610
rect 188436 153546 188488 153552
rect 188356 153513 188384 153546
rect 188342 153504 188398 153513
rect 188342 153439 188398 153448
rect 187884 152924 187936 152930
rect 187884 152866 187936 152872
rect 187976 152924 188028 152930
rect 187976 152866 188028 152872
rect 187896 150090 187924 152866
rect 188540 150226 188568 157830
rect 189170 155952 189226 155961
rect 189644 155922 189672 163200
rect 190472 157758 190500 163200
rect 191300 159934 191328 163200
rect 191748 159996 191800 160002
rect 191748 159938 191800 159944
rect 191288 159928 191340 159934
rect 191288 159870 191340 159876
rect 190644 157820 190696 157826
rect 190644 157762 190696 157768
rect 190460 157752 190512 157758
rect 190460 157694 190512 157700
rect 190656 157334 190684 157762
rect 191760 157334 191788 159938
rect 190656 157306 191144 157334
rect 189816 156392 189868 156398
rect 189816 156334 189868 156340
rect 189170 155887 189226 155896
rect 189632 155916 189684 155922
rect 188540 150198 188614 150226
rect 187252 150062 187326 150090
rect 187896 150062 187970 150090
rect 187298 149940 187326 150062
rect 187942 149940 187970 150062
rect 188586 149940 188614 150198
rect 189184 150090 189212 155887
rect 189632 155858 189684 155864
rect 189828 150090 189856 156334
rect 190460 152176 190512 152182
rect 190460 152118 190512 152124
rect 190472 150090 190500 152118
rect 191116 150226 191144 157306
rect 191668 157306 191788 157334
rect 191288 154488 191340 154494
rect 191288 154430 191340 154436
rect 191300 154358 191328 154430
rect 191472 154420 191524 154426
rect 191472 154362 191524 154368
rect 191288 154352 191340 154358
rect 191288 154294 191340 154300
rect 191380 154352 191432 154358
rect 191484 154329 191512 154362
rect 191380 154294 191432 154300
rect 191470 154320 191526 154329
rect 191392 153474 191420 154294
rect 191470 154255 191526 154264
rect 191380 153468 191432 153474
rect 191380 153410 191432 153416
rect 191668 151910 191696 157306
rect 192128 157282 192156 163200
rect 192116 157276 192168 157282
rect 192116 157218 192168 157224
rect 192956 155174 192984 163200
rect 193784 159186 193812 163200
rect 193128 159180 193180 159186
rect 193128 159122 193180 159128
rect 193772 159180 193824 159186
rect 193772 159122 193824 159128
rect 192944 155168 192996 155174
rect 192944 155110 192996 155116
rect 191748 155100 191800 155106
rect 191748 155042 191800 155048
rect 191656 151904 191708 151910
rect 191656 151846 191708 151852
rect 191116 150198 191190 150226
rect 189184 150062 189258 150090
rect 189828 150062 189902 150090
rect 190472 150062 190546 150090
rect 189230 149940 189258 150062
rect 189874 149940 189902 150062
rect 190518 149940 190546 150062
rect 191162 149940 191190 150198
rect 191760 150090 191788 155042
rect 192390 153504 192446 153513
rect 192390 153439 192446 153448
rect 192404 150090 192432 153439
rect 193036 152992 193088 152998
rect 193036 152934 193088 152940
rect 193048 150090 193076 152934
rect 193140 152114 193168 159122
rect 194704 158846 194732 163200
rect 195152 158908 195204 158914
rect 195152 158850 195204 158856
rect 194508 158840 194560 158846
rect 194508 158782 194560 158788
rect 194692 158840 194744 158846
rect 194692 158782 194744 158788
rect 193220 157616 193272 157622
rect 193220 157558 193272 157564
rect 193232 157334 193260 157558
rect 193232 157306 193720 157334
rect 193128 152108 193180 152114
rect 193128 152050 193180 152056
rect 193692 150226 193720 157306
rect 194324 155032 194376 155038
rect 194324 154974 194376 154980
rect 193692 150198 193766 150226
rect 191760 150062 191834 150090
rect 192404 150062 192478 150090
rect 193048 150062 193122 150090
rect 191806 149940 191834 150062
rect 192450 149940 192478 150062
rect 193094 149940 193122 150062
rect 193738 149940 193766 150198
rect 194336 150090 194364 154974
rect 194520 153474 194548 158782
rect 194968 155100 195020 155106
rect 194968 155042 195020 155048
rect 194508 153468 194560 153474
rect 194508 153410 194560 153416
rect 194980 150090 195008 155042
rect 195164 152182 195192 158850
rect 195532 157826 195560 163200
rect 195520 157820 195572 157826
rect 195520 157762 195572 157768
rect 196256 156324 196308 156330
rect 196256 156266 196308 156272
rect 195612 152244 195664 152250
rect 195612 152186 195664 152192
rect 195152 152176 195204 152182
rect 195152 152118 195204 152124
rect 195624 150090 195652 152186
rect 195888 152108 195940 152114
rect 195888 152050 195940 152056
rect 195900 151910 195928 152050
rect 195888 151904 195940 151910
rect 195888 151846 195940 151852
rect 196268 150226 196296 156266
rect 196360 155106 196388 163200
rect 196992 159316 197044 159322
rect 196992 159258 197044 159264
rect 196348 155100 196400 155106
rect 196348 155042 196400 155048
rect 197004 153542 197032 159258
rect 197188 158982 197216 163200
rect 198016 160002 198044 163200
rect 198004 159996 198056 160002
rect 198004 159938 198056 159944
rect 197176 158976 197228 158982
rect 197176 158918 197228 158924
rect 197360 158772 197412 158778
rect 197360 158714 197412 158720
rect 197372 157622 197400 158714
rect 198738 158536 198794 158545
rect 198738 158471 198794 158480
rect 197360 157616 197412 157622
rect 197360 157558 197412 157564
rect 197544 153604 197596 153610
rect 197544 153546 197596 153552
rect 196900 153536 196952 153542
rect 196900 153478 196952 153484
rect 196992 153536 197044 153542
rect 196992 153478 197044 153484
rect 196912 150226 196940 153478
rect 197556 150226 197584 153546
rect 198188 153128 198240 153134
rect 198188 153070 198240 153076
rect 198200 150226 198228 153070
rect 198752 151814 198780 158471
rect 198844 156534 198872 163200
rect 198924 160064 198976 160070
rect 198924 160006 198976 160012
rect 198832 156528 198884 156534
rect 198832 156470 198884 156476
rect 198936 153610 198964 160006
rect 199672 155038 199700 163200
rect 200592 161474 200620 163200
rect 200592 161446 200712 161474
rect 200684 159050 200712 161446
rect 201420 159322 201448 163200
rect 201408 159316 201460 159322
rect 201408 159258 201460 159264
rect 200672 159044 200724 159050
rect 200672 158986 200724 158992
rect 200396 158908 200448 158914
rect 200396 158850 200448 158856
rect 200304 156256 200356 156262
rect 200304 156198 200356 156204
rect 199660 155032 199712 155038
rect 199660 154974 199712 154980
rect 200120 154488 200172 154494
rect 200120 154430 200172 154436
rect 198924 153604 198976 153610
rect 198924 153546 198976 153552
rect 199384 153536 199436 153542
rect 199436 153484 199608 153490
rect 199384 153478 199608 153484
rect 199396 153462 199608 153478
rect 199580 153406 199608 153462
rect 199476 153400 199528 153406
rect 199476 153342 199528 153348
rect 199568 153400 199620 153406
rect 199568 153342 199620 153348
rect 198752 151786 198872 151814
rect 198844 150226 198872 151786
rect 199488 150226 199516 153342
rect 200132 150226 200160 154430
rect 196268 150198 196342 150226
rect 196912 150198 196986 150226
rect 197556 150198 197630 150226
rect 198200 150198 198274 150226
rect 198844 150198 198918 150226
rect 199488 150198 199562 150226
rect 200132 150198 200206 150226
rect 200316 150210 200344 156198
rect 200408 153542 200436 158850
rect 201316 156664 201368 156670
rect 201316 156606 201368 156612
rect 201328 156466 201356 156606
rect 201316 156460 201368 156466
rect 201316 156402 201368 156408
rect 202248 156398 202276 163200
rect 202236 156392 202288 156398
rect 202236 156334 202288 156340
rect 203076 156262 203104 163200
rect 203904 159118 203932 163200
rect 204732 159361 204760 163200
rect 204718 159352 204774 159361
rect 204718 159287 204774 159296
rect 203800 159112 203852 159118
rect 203800 159054 203852 159060
rect 203892 159112 203944 159118
rect 203892 159054 203944 159060
rect 203812 158914 203840 159054
rect 203800 158908 203852 158914
rect 203800 158850 203852 158856
rect 204904 158908 204956 158914
rect 204904 158850 204956 158856
rect 203708 158840 203760 158846
rect 203708 158782 203760 158788
rect 203432 157548 203484 157554
rect 203432 157490 203484 157496
rect 203064 156256 203116 156262
rect 203064 156198 203116 156204
rect 202696 154420 202748 154426
rect 202696 154362 202748 154368
rect 202052 154352 202104 154358
rect 202052 154294 202104 154300
rect 200396 153536 200448 153542
rect 200396 153478 200448 153484
rect 200764 151972 200816 151978
rect 200764 151914 200816 151920
rect 200776 150226 200804 151914
rect 202064 150226 202092 154294
rect 202708 150226 202736 154362
rect 203340 152040 203392 152046
rect 203340 151982 203392 151988
rect 203352 150226 203380 151982
rect 203444 151814 203472 157490
rect 203720 152998 203748 158782
rect 204916 157554 204944 158850
rect 204904 157548 204956 157554
rect 204904 157490 204956 157496
rect 204904 157344 204956 157350
rect 204258 157312 204314 157321
rect 204904 157286 204956 157292
rect 204996 157344 205048 157350
rect 204996 157286 205048 157292
rect 204258 157247 204314 157256
rect 203708 152992 203760 152998
rect 203708 152934 203760 152940
rect 203444 151786 204024 151814
rect 203996 150226 204024 151786
rect 194336 150062 194410 150090
rect 194980 150062 195054 150090
rect 195624 150062 195698 150090
rect 194382 149940 194410 150062
rect 195026 149940 195054 150062
rect 195670 149940 195698 150062
rect 196314 149940 196342 150198
rect 196958 149940 196986 150198
rect 197602 149940 197630 150198
rect 198246 149940 198274 150198
rect 198890 149940 198918 150198
rect 199534 149940 199562 150198
rect 200178 149940 200206 150198
rect 200304 150204 200356 150210
rect 200776 150198 200850 150226
rect 200304 150146 200356 150152
rect 200822 149940 200850 150198
rect 201454 150204 201506 150210
rect 202064 150198 202138 150226
rect 202708 150198 202782 150226
rect 203352 150198 203426 150226
rect 203996 150198 204070 150226
rect 204272 150210 204300 157247
rect 204916 156534 204944 157286
rect 204904 156528 204956 156534
rect 204904 156470 204956 156476
rect 205008 156398 205036 157286
rect 204996 156392 205048 156398
rect 204996 156334 205048 156340
rect 204628 155848 204680 155854
rect 204628 155790 204680 155796
rect 204640 150226 204668 155790
rect 205560 154358 205588 163200
rect 206480 155854 206508 163200
rect 207308 158778 207336 163200
rect 208136 158846 208164 163200
rect 208124 158840 208176 158846
rect 208124 158782 208176 158788
rect 207296 158772 207348 158778
rect 207296 158714 207348 158720
rect 206560 157480 206612 157486
rect 206560 157422 206612 157428
rect 206468 155848 206520 155854
rect 206468 155790 206520 155796
rect 205548 154352 205600 154358
rect 205548 154294 205600 154300
rect 205916 153196 205968 153202
rect 205916 153138 205968 153144
rect 205928 150226 205956 153138
rect 206572 150226 206600 157422
rect 208964 154426 208992 163200
rect 209792 156398 209820 163200
rect 210620 159118 210648 163200
rect 211448 160070 211476 163200
rect 211436 160064 211488 160070
rect 211436 160006 211488 160012
rect 210516 159112 210568 159118
rect 210516 159054 210568 159060
rect 210608 159112 210660 159118
rect 210608 159054 210660 159060
rect 210528 158914 210556 159054
rect 210516 158908 210568 158914
rect 210516 158850 210568 158856
rect 211988 158840 212040 158846
rect 211988 158782 212040 158788
rect 211620 156460 211672 156466
rect 211620 156402 211672 156408
rect 209780 156392 209832 156398
rect 209780 156334 209832 156340
rect 209136 156188 209188 156194
rect 209136 156130 209188 156136
rect 208952 154420 209004 154426
rect 208952 154362 209004 154368
rect 207204 153332 207256 153338
rect 207204 153274 207256 153280
rect 207216 150226 207244 153274
rect 207848 153264 207900 153270
rect 207848 153206 207900 153212
rect 207860 150226 207888 153206
rect 208492 152108 208544 152114
rect 208492 152050 208544 152056
rect 208504 150226 208532 152050
rect 209148 150226 209176 156130
rect 211252 155372 211304 155378
rect 211252 155314 211304 155320
rect 209780 153944 209832 153950
rect 209780 153886 209832 153892
rect 209792 150226 209820 153886
rect 210424 153740 210476 153746
rect 210424 153682 210476 153688
rect 210436 150226 210464 153682
rect 211068 152516 211120 152522
rect 211068 152458 211120 152464
rect 211080 150226 211108 152458
rect 201454 150146 201506 150152
rect 201466 149940 201494 150146
rect 202110 149940 202138 150198
rect 202754 149940 202782 150198
rect 203398 149940 203426 150198
rect 204042 149940 204070 150198
rect 204260 150204 204312 150210
rect 204640 150198 204714 150226
rect 204260 150146 204312 150152
rect 204686 149940 204714 150198
rect 205318 150204 205370 150210
rect 205928 150198 206002 150226
rect 206572 150198 206646 150226
rect 207216 150198 207290 150226
rect 207860 150198 207934 150226
rect 208504 150198 208578 150226
rect 209148 150198 209222 150226
rect 209792 150198 209866 150226
rect 210436 150198 210510 150226
rect 211080 150198 211154 150226
rect 211264 150210 211292 155314
rect 211632 150226 211660 156402
rect 212000 152522 212028 158782
rect 212368 153785 212396 163200
rect 212632 159316 212684 159322
rect 212632 159258 212684 159264
rect 212354 153776 212410 153785
rect 212354 153711 212410 153720
rect 211988 152516 212040 152522
rect 211988 152458 212040 152464
rect 212644 152046 212672 159258
rect 213196 156194 213224 163200
rect 214024 159322 214052 163200
rect 214012 159316 214064 159322
rect 214012 159258 214064 159264
rect 213736 158908 213788 158914
rect 214748 158908 214800 158914
rect 213736 158850 213788 158856
rect 214576 158868 214748 158896
rect 213184 156188 213236 156194
rect 213184 156130 213236 156136
rect 212908 153808 212960 153814
rect 212908 153750 212960 153756
rect 212632 152040 212684 152046
rect 212632 151982 212684 151988
rect 212920 150226 212948 153750
rect 213748 152182 213776 158850
rect 214576 158778 214604 158868
rect 214748 158850 214800 158856
rect 214852 158846 214880 163200
rect 215300 159112 215352 159118
rect 215300 159054 215352 159060
rect 214840 158840 214892 158846
rect 214840 158782 214892 158788
rect 214564 158772 214616 158778
rect 214564 158714 214616 158720
rect 213828 156936 213880 156942
rect 213828 156878 213880 156884
rect 213920 156936 213972 156942
rect 213920 156878 213972 156884
rect 213840 155378 213868 156878
rect 213932 156534 213960 156878
rect 213920 156528 213972 156534
rect 213920 156470 213972 156476
rect 214564 156528 214616 156534
rect 214564 156470 214616 156476
rect 214576 156262 214604 156470
rect 214564 156256 214616 156262
rect 214564 156198 214616 156204
rect 213920 156120 213972 156126
rect 213920 156062 213972 156068
rect 213828 155372 213880 155378
rect 213828 155314 213880 155320
rect 213552 152176 213604 152182
rect 213552 152118 213604 152124
rect 213736 152176 213788 152182
rect 213736 152118 213788 152124
rect 213564 150226 213592 152118
rect 213932 151814 213960 156062
rect 214840 155304 214892 155310
rect 214840 155246 214892 155252
rect 213932 151786 214236 151814
rect 214208 150226 214236 151786
rect 214852 150226 214880 155246
rect 215312 153134 215340 159054
rect 215680 153950 215708 163200
rect 216508 156398 216536 163200
rect 216680 159248 216732 159254
rect 216680 159190 216732 159196
rect 216496 156392 216548 156398
rect 216496 156334 216548 156340
rect 216692 155378 216720 159190
rect 217336 158982 217364 163200
rect 218256 159254 218284 163200
rect 219084 163146 219112 163200
rect 219176 163146 219204 163254
rect 219084 163118 219204 163146
rect 218244 159248 218296 159254
rect 218244 159190 218296 159196
rect 217324 158976 217376 158982
rect 217324 158918 217376 158924
rect 218244 158024 218296 158030
rect 218244 157966 218296 157972
rect 216772 156800 216824 156806
rect 216772 156742 216824 156748
rect 216680 155372 216732 155378
rect 216680 155314 216732 155320
rect 215668 153944 215720 153950
rect 215668 153886 215720 153892
rect 215484 153672 215536 153678
rect 215484 153614 215536 153620
rect 215300 153128 215352 153134
rect 215300 153070 215352 153076
rect 205318 150146 205370 150152
rect 205330 149940 205358 150146
rect 205974 149940 206002 150198
rect 206618 149940 206646 150198
rect 207262 149940 207290 150198
rect 207906 149940 207934 150198
rect 208550 149940 208578 150198
rect 209194 149940 209222 150198
rect 209838 149940 209866 150198
rect 210482 149940 210510 150198
rect 211126 149940 211154 150198
rect 211252 150204 211304 150210
rect 211632 150198 211706 150226
rect 211252 150146 211304 150152
rect 211678 149940 211706 150198
rect 212310 150204 212362 150210
rect 212920 150198 212994 150226
rect 213564 150198 213638 150226
rect 214208 150198 214282 150226
rect 214852 150198 214926 150226
rect 212310 150146 212362 150152
rect 212322 149940 212350 150146
rect 212966 149940 212994 150198
rect 213610 149940 213638 150198
rect 214254 149940 214282 150198
rect 214898 149940 214926 150198
rect 215496 150090 215524 153614
rect 216128 152652 216180 152658
rect 216128 152594 216180 152600
rect 216140 150090 216168 152594
rect 216784 150090 216812 156742
rect 217416 155236 217468 155242
rect 217416 155178 217468 155184
rect 217428 150090 217456 155178
rect 218060 153876 218112 153882
rect 218060 153818 218112 153824
rect 218072 150090 218100 153818
rect 218256 150210 218284 157966
rect 219360 153882 219388 163254
rect 219898 163200 219954 164400
rect 220726 163200 220782 164400
rect 221554 163200 221610 164400
rect 222382 163200 222438 164400
rect 223210 163200 223266 164400
rect 224130 163200 224186 164400
rect 224958 163200 225014 164400
rect 225786 163200 225842 164400
rect 226614 163200 226670 164400
rect 227442 163200 227498 164400
rect 228270 163200 228326 164400
rect 229098 163200 229154 164400
rect 230018 163200 230074 164400
rect 230846 163200 230902 164400
rect 231674 163200 231730 164400
rect 232502 163200 232558 164400
rect 233330 163200 233386 164400
rect 234158 163200 234214 164400
rect 234264 163254 234476 163282
rect 219912 156806 219940 163200
rect 220636 159180 220688 159186
rect 220636 159122 220688 159128
rect 220452 158976 220504 158982
rect 220452 158918 220504 158924
rect 219900 156800 219952 156806
rect 219900 156742 219952 156748
rect 219992 156732 220044 156738
rect 219992 156674 220044 156680
rect 219900 156664 219952 156670
rect 219900 156606 219952 156612
rect 219912 156126 219940 156606
rect 219900 156120 219952 156126
rect 219900 156062 219952 156068
rect 219348 153876 219400 153882
rect 219348 153818 219400 153824
rect 218704 152244 218756 152250
rect 218704 152186 218756 152192
rect 218244 150204 218296 150210
rect 218244 150146 218296 150152
rect 218716 150090 218744 152186
rect 219394 150204 219446 150210
rect 219394 150146 219446 150152
rect 215496 150062 215570 150090
rect 216140 150062 216214 150090
rect 216784 150062 216858 150090
rect 217428 150062 217502 150090
rect 218072 150062 218146 150090
rect 218716 150062 218790 150090
rect 215542 149940 215570 150062
rect 216186 149940 216214 150062
rect 216830 149940 216858 150062
rect 217474 149940 217502 150062
rect 218118 149940 218146 150062
rect 218762 149940 218790 150062
rect 219406 149940 219434 150146
rect 220004 150090 220032 156674
rect 220084 156664 220136 156670
rect 220084 156606 220136 156612
rect 220096 156194 220124 156606
rect 220084 156188 220136 156194
rect 220084 156130 220136 156136
rect 220464 152658 220492 158918
rect 220648 156194 220676 159122
rect 220740 159118 220768 163200
rect 220728 159112 220780 159118
rect 220728 159054 220780 159060
rect 221568 158846 221596 163200
rect 221464 158840 221516 158846
rect 221464 158782 221516 158788
rect 221556 158840 221608 158846
rect 221556 158782 221608 158788
rect 220636 156188 220688 156194
rect 220636 156130 220688 156136
rect 220544 156120 220596 156126
rect 220544 156062 220596 156068
rect 220452 152652 220504 152658
rect 220452 152594 220504 152600
rect 220556 150226 220584 156062
rect 221280 152720 221332 152726
rect 221280 152662 221332 152668
rect 220556 150198 220722 150226
rect 220004 150062 220078 150090
rect 220050 149940 220078 150062
rect 220694 149940 220722 150198
rect 221292 150090 221320 152662
rect 221476 152250 221504 158782
rect 222108 158772 222160 158778
rect 222108 158714 222160 158720
rect 222120 156262 222148 158714
rect 222108 156256 222160 156262
rect 222108 156198 222160 156204
rect 221924 155304 221976 155310
rect 221924 155246 221976 155252
rect 221464 152244 221516 152250
rect 221464 152186 221516 152192
rect 221936 150090 221964 155246
rect 222396 153814 222424 163200
rect 223120 156936 223172 156942
rect 223120 156878 223172 156884
rect 222568 156868 222620 156874
rect 222568 156810 222620 156816
rect 222384 153808 222436 153814
rect 222384 153750 222436 153756
rect 222580 150090 222608 156810
rect 223132 150226 223160 156878
rect 223224 156738 223252 163200
rect 223580 159384 223632 159390
rect 223580 159326 223632 159332
rect 223592 157334 223620 159326
rect 224144 159186 224172 163200
rect 224972 159390 225000 163200
rect 225800 161474 225828 163200
rect 225800 161446 225920 161474
rect 225052 159520 225104 159526
rect 225052 159462 225104 159468
rect 224960 159384 225012 159390
rect 224960 159326 225012 159332
rect 224132 159180 224184 159186
rect 224132 159122 224184 159128
rect 224776 158840 224828 158846
rect 224776 158782 224828 158788
rect 223592 157306 223896 157334
rect 223212 156732 223264 156738
rect 223212 156674 223264 156680
rect 223868 150226 223896 157306
rect 224500 156052 224552 156058
rect 224500 155994 224552 156000
rect 224512 150226 224540 155994
rect 224788 152726 224816 158782
rect 225064 153202 225092 159462
rect 225144 157004 225196 157010
rect 225144 156946 225196 156952
rect 225052 153196 225104 153202
rect 225052 153138 225104 153144
rect 224776 152720 224828 152726
rect 224776 152662 224828 152668
rect 225156 150226 225184 156946
rect 225788 154556 225840 154562
rect 225788 154498 225840 154504
rect 225800 150226 225828 154498
rect 225892 154494 225920 161446
rect 226628 156942 226656 163200
rect 227076 157412 227128 157418
rect 227076 157354 227128 157360
rect 226616 156936 226668 156942
rect 226616 156878 226668 156884
rect 225880 154488 225932 154494
rect 225880 154430 225932 154436
rect 226432 152584 226484 152590
rect 226432 152526 226484 152532
rect 226444 150226 226472 152526
rect 227088 150226 227116 157354
rect 227456 152425 227484 163200
rect 227720 159044 227772 159050
rect 227720 158986 227772 158992
rect 227732 156126 227760 158986
rect 227720 156120 227772 156126
rect 227720 156062 227772 156068
rect 227720 155440 227772 155446
rect 227720 155382 227772 155388
rect 227442 152416 227498 152425
rect 227442 152351 227498 152360
rect 227732 150226 227760 155382
rect 228284 152590 228312 163200
rect 228364 155984 228416 155990
rect 228364 155926 228416 155932
rect 228272 152584 228324 152590
rect 228272 152526 228324 152532
rect 228376 150226 228404 155926
rect 229112 153746 229140 163200
rect 229652 157072 229704 157078
rect 229652 157014 229704 157020
rect 229192 154896 229244 154902
rect 229192 154838 229244 154844
rect 229100 153740 229152 153746
rect 229100 153682 229152 153688
rect 229008 153196 229060 153202
rect 229008 153138 229060 153144
rect 229020 150226 229048 153138
rect 223132 150198 223298 150226
rect 223868 150198 223942 150226
rect 224512 150198 224586 150226
rect 225156 150198 225230 150226
rect 225800 150198 225874 150226
rect 226444 150198 226518 150226
rect 227088 150198 227162 150226
rect 227732 150198 227806 150226
rect 228376 150198 228450 150226
rect 229020 150198 229094 150226
rect 229204 150210 229232 154838
rect 229664 150226 229692 157014
rect 230032 156874 230060 163200
rect 230860 159050 230888 163200
rect 231688 159526 231716 163200
rect 231676 159520 231728 159526
rect 231676 159462 231728 159468
rect 230848 159044 230900 159050
rect 230848 158986 230900 158992
rect 231308 158840 231360 158846
rect 231308 158782 231360 158788
rect 230020 156868 230072 156874
rect 230020 156810 230072 156816
rect 230940 156324 230992 156330
rect 230940 156266 230992 156272
rect 230952 150226 230980 156266
rect 231320 154902 231348 158782
rect 231860 158092 231912 158098
rect 231860 158034 231912 158040
rect 231308 154896 231360 154902
rect 231308 154838 231360 154844
rect 231584 152448 231636 152454
rect 231584 152390 231636 152396
rect 231596 150226 231624 152390
rect 231872 151814 231900 158034
rect 232516 154562 232544 163200
rect 233344 158098 233372 163200
rect 234172 163146 234200 163200
rect 234264 163146 234292 163254
rect 234172 163118 234292 163146
rect 234160 159452 234212 159458
rect 234160 159394 234212 159400
rect 233332 158092 233384 158098
rect 233332 158034 233384 158040
rect 232872 154828 232924 154834
rect 232872 154770 232924 154776
rect 232504 154556 232556 154562
rect 232504 154498 232556 154504
rect 231872 151786 232268 151814
rect 232240 150226 232268 151786
rect 232884 150226 232912 154770
rect 233516 154012 233568 154018
rect 233516 153954 233568 153960
rect 233528 150226 233556 153954
rect 234172 150226 234200 159394
rect 234448 153202 234476 163254
rect 234986 163200 235042 164400
rect 235906 163200 235962 164400
rect 236734 163200 236790 164400
rect 237562 163200 237618 164400
rect 238390 163200 238446 164400
rect 239218 163200 239274 164400
rect 240046 163200 240102 164400
rect 240874 163200 240930 164400
rect 241794 163200 241850 164400
rect 242622 163200 242678 164400
rect 243450 163200 243506 164400
rect 244278 163200 244334 164400
rect 245106 163200 245162 164400
rect 245934 163200 245990 164400
rect 246762 163200 246818 164400
rect 247682 163200 247738 164400
rect 248510 163200 248566 164400
rect 249338 163200 249394 164400
rect 249444 163254 249748 163282
rect 235000 159458 235028 163200
rect 234988 159452 235040 159458
rect 234988 159394 235040 159400
rect 234804 157140 234856 157146
rect 234804 157082 234856 157088
rect 234436 153196 234488 153202
rect 234436 153138 234488 153144
rect 234816 150226 234844 157082
rect 235448 154080 235500 154086
rect 235448 154022 235500 154028
rect 235460 150226 235488 154022
rect 235920 154018 235948 163200
rect 236092 157684 236144 157690
rect 236092 157626 236144 157632
rect 235908 154012 235960 154018
rect 235908 153954 235960 153960
rect 236104 150226 236132 157626
rect 236748 155242 236776 163200
rect 237576 158846 237604 163200
rect 238404 158982 238432 163200
rect 238392 158976 238444 158982
rect 238392 158918 238444 158924
rect 237564 158840 237616 158846
rect 237564 158782 237616 158788
rect 238852 158228 238904 158234
rect 238852 158170 238904 158176
rect 237380 158160 237432 158166
rect 237380 158102 237432 158108
rect 236736 155236 236788 155242
rect 236736 155178 236788 155184
rect 236736 152788 236788 152794
rect 236736 152730 236788 152736
rect 236748 150226 236776 152730
rect 237392 150226 237420 158102
rect 238024 154760 238076 154766
rect 238024 154702 238076 154708
rect 238036 150226 238064 154702
rect 238668 153468 238720 153474
rect 238668 153410 238720 153416
rect 238680 150226 238708 153410
rect 221292 150062 221366 150090
rect 221936 150062 222010 150090
rect 222580 150062 222654 150090
rect 221338 149940 221366 150062
rect 221982 149940 222010 150062
rect 222626 149940 222654 150062
rect 223270 149940 223298 150198
rect 223914 149940 223942 150198
rect 224558 149940 224586 150198
rect 225202 149940 225230 150198
rect 225846 149940 225874 150198
rect 226490 149940 226518 150198
rect 227134 149940 227162 150198
rect 227778 149940 227806 150198
rect 228422 149940 228450 150198
rect 229066 149940 229094 150198
rect 229192 150204 229244 150210
rect 229664 150198 229738 150226
rect 229192 150146 229244 150152
rect 229710 149940 229738 150198
rect 230342 150204 230394 150210
rect 230952 150198 231026 150226
rect 231596 150198 231670 150226
rect 232240 150198 232314 150226
rect 232884 150198 232958 150226
rect 233528 150198 233602 150226
rect 234172 150198 234246 150226
rect 234816 150198 234890 150226
rect 235460 150198 235534 150226
rect 236104 150198 236178 150226
rect 236748 150198 236822 150226
rect 237392 150198 237466 150226
rect 238036 150198 238110 150226
rect 238680 150198 238754 150226
rect 238864 150210 238892 158170
rect 239232 153678 239260 163200
rect 239312 159588 239364 159594
rect 239312 159530 239364 159536
rect 239220 153672 239272 153678
rect 239220 153614 239272 153620
rect 239324 150226 239352 159530
rect 240060 158030 240088 163200
rect 240324 159656 240376 159662
rect 240324 159598 240376 159604
rect 240048 158024 240100 158030
rect 240048 157966 240100 157972
rect 240140 154624 240192 154630
rect 240140 154566 240192 154572
rect 240152 151814 240180 154566
rect 240336 152794 240364 159598
rect 240888 158778 240916 163200
rect 241808 159662 241836 163200
rect 241796 159656 241848 159662
rect 241796 159598 241848 159604
rect 242440 158976 242492 158982
rect 242440 158918 242492 158924
rect 240876 158772 240928 158778
rect 240876 158714 240928 158720
rect 242072 158296 242124 158302
rect 242072 158238 242124 158244
rect 240692 154964 240744 154970
rect 240692 154906 240744 154912
rect 240324 152788 240376 152794
rect 240324 152730 240376 152736
rect 240704 151814 240732 154906
rect 241888 152788 241940 152794
rect 241888 152730 241940 152736
rect 240152 151786 240640 151814
rect 240704 151786 241284 151814
rect 240612 150226 240640 151786
rect 241256 150226 241284 151786
rect 241900 150226 241928 152730
rect 242084 151814 242112 158238
rect 242452 152046 242480 158918
rect 242636 154086 242664 163200
rect 243360 158772 243412 158778
rect 243360 158714 243412 158720
rect 243084 154692 243136 154698
rect 243084 154634 243136 154640
rect 242624 154080 242676 154086
rect 242624 154022 242676 154028
rect 242440 152040 242492 152046
rect 242440 151982 242492 151988
rect 242084 151786 242480 151814
rect 242452 150226 242480 151786
rect 243096 150226 243124 154634
rect 243372 151978 243400 158714
rect 243464 155310 243492 163200
rect 244292 158846 244320 163200
rect 244280 158840 244332 158846
rect 244280 158782 244332 158788
rect 245016 158364 245068 158370
rect 245016 158306 245068 158312
rect 243452 155304 243504 155310
rect 243452 155246 243504 155252
rect 243728 153400 243780 153406
rect 243728 153342 243780 153348
rect 243360 151972 243412 151978
rect 243360 151914 243412 151920
rect 243740 150226 243768 153342
rect 244372 152380 244424 152386
rect 244372 152322 244424 152328
rect 244384 150226 244412 152322
rect 245028 150226 245056 158306
rect 245120 152454 245148 163200
rect 245844 159724 245896 159730
rect 245844 159666 245896 159672
rect 245660 154148 245712 154154
rect 245660 154090 245712 154096
rect 245108 152448 245160 152454
rect 245108 152390 245160 152396
rect 245672 150226 245700 154090
rect 230342 150146 230394 150152
rect 230354 149940 230382 150146
rect 230998 149940 231026 150198
rect 231642 149940 231670 150198
rect 232286 149940 232314 150198
rect 232930 149940 232958 150198
rect 233574 149940 233602 150198
rect 234218 149940 234246 150198
rect 234862 149940 234890 150198
rect 235506 149940 235534 150198
rect 236150 149940 236178 150198
rect 236794 149940 236822 150198
rect 237438 149940 237466 150198
rect 238082 149940 238110 150198
rect 238726 149940 238754 150198
rect 238852 150204 238904 150210
rect 239324 150198 239398 150226
rect 238852 150146 238904 150152
rect 239370 149940 239398 150198
rect 240002 150204 240054 150210
rect 240612 150198 240686 150226
rect 241256 150198 241330 150226
rect 241900 150198 241974 150226
rect 242452 150198 242526 150226
rect 243096 150198 243170 150226
rect 243740 150198 243814 150226
rect 244384 150198 244458 150226
rect 245028 150198 245102 150226
rect 245672 150198 245746 150226
rect 245856 150210 245884 159666
rect 245948 154154 245976 163200
rect 246776 158166 246804 163200
rect 247592 158432 247644 158438
rect 247592 158374 247644 158380
rect 246764 158160 246816 158166
rect 246764 158102 246816 158108
rect 246304 157208 246356 157214
rect 246304 157150 246356 157156
rect 245936 154148 245988 154154
rect 245936 154090 245988 154096
rect 246316 150226 246344 157150
rect 247132 155508 247184 155514
rect 247132 155450 247184 155456
rect 240002 150146 240054 150152
rect 240014 149940 240042 150146
rect 240658 149940 240686 150198
rect 241302 149940 241330 150198
rect 241946 149940 241974 150198
rect 242498 149940 242526 150198
rect 243142 149940 243170 150198
rect 243786 149940 243814 150198
rect 244430 149940 244458 150198
rect 245074 149940 245102 150198
rect 245718 149940 245746 150198
rect 245844 150204 245896 150210
rect 246316 150198 246390 150226
rect 247144 150210 247172 155450
rect 247604 150226 247632 158374
rect 247696 152794 247724 163200
rect 248524 159730 248552 163200
rect 249352 163146 249380 163200
rect 249444 163146 249472 163254
rect 249352 163118 249472 163146
rect 248512 159724 248564 159730
rect 248512 159666 248564 159672
rect 249720 153610 249748 163254
rect 250166 163200 250222 164400
rect 250994 163200 251050 164400
rect 251822 163200 251878 164400
rect 251928 163254 252232 163282
rect 250076 158636 250128 158642
rect 250076 158578 250128 158584
rect 248880 153604 248932 153610
rect 248880 153546 248932 153552
rect 249708 153604 249760 153610
rect 249708 153546 249760 153552
rect 247684 152788 247736 152794
rect 247684 152730 247736 152736
rect 248892 150226 248920 153546
rect 249524 152312 249576 152318
rect 249524 152254 249576 152260
rect 249536 150226 249564 152254
rect 250088 151814 250116 158578
rect 250180 155446 250208 163200
rect 251008 159594 251036 163200
rect 251836 163146 251864 163200
rect 251928 163146 251956 163254
rect 251836 163118 251956 163146
rect 250996 159588 251048 159594
rect 250996 159530 251048 159536
rect 251456 157616 251508 157622
rect 251456 157558 251508 157564
rect 250168 155440 250220 155446
rect 250168 155382 250220 155388
rect 250812 154216 250864 154222
rect 250812 154158 250864 154164
rect 250088 151786 250208 151814
rect 250180 150226 250208 151786
rect 250824 150226 250852 154158
rect 251468 150226 251496 157558
rect 252204 152862 252232 163254
rect 252650 163200 252706 164400
rect 253570 163200 253626 164400
rect 254398 163200 254454 164400
rect 255226 163200 255282 164400
rect 256054 163200 256110 164400
rect 256882 163200 256938 164400
rect 257710 163200 257766 164400
rect 258538 163200 258594 164400
rect 259458 163200 259514 164400
rect 260286 163200 260342 164400
rect 261114 163200 261170 164400
rect 261942 163200 261998 164400
rect 262770 163200 262826 164400
rect 263598 163200 263654 164400
rect 264426 163200 264482 164400
rect 265346 163200 265402 164400
rect 266174 163200 266230 164400
rect 267002 163200 267058 164400
rect 267830 163200 267886 164400
rect 268658 163200 268714 164400
rect 269486 163200 269542 164400
rect 270314 163200 270370 164400
rect 271234 163200 271290 164400
rect 272062 163200 272118 164400
rect 272168 163254 272656 163282
rect 252560 158500 252612 158506
rect 252560 158442 252612 158448
rect 252100 152856 252152 152862
rect 252100 152798 252152 152804
rect 252192 152856 252244 152862
rect 252192 152798 252244 152804
rect 252112 150226 252140 152798
rect 252572 151814 252600 158442
rect 252664 154222 252692 163200
rect 253388 155644 253440 155650
rect 253388 155586 253440 155592
rect 252652 154216 252704 154222
rect 252652 154158 252704 154164
rect 252572 151786 252784 151814
rect 252756 150226 252784 151786
rect 253400 150226 253428 155586
rect 253584 154970 253612 163200
rect 253940 159792 253992 159798
rect 253940 159734 253992 159740
rect 253572 154964 253624 154970
rect 253572 154906 253624 154912
rect 245844 150146 245896 150152
rect 246362 149940 246390 150198
rect 246994 150204 247046 150210
rect 246994 150146 247046 150152
rect 247132 150204 247184 150210
rect 247604 150198 247678 150226
rect 247132 150146 247184 150152
rect 247006 149940 247034 150146
rect 247650 149940 247678 150198
rect 248282 150204 248334 150210
rect 248892 150198 248966 150226
rect 249536 150198 249610 150226
rect 250180 150198 250254 150226
rect 250824 150198 250898 150226
rect 251468 150198 251542 150226
rect 252112 150198 252186 150226
rect 252756 150198 252830 150226
rect 253400 150198 253474 150226
rect 253952 150210 253980 159734
rect 254412 158778 254440 163200
rect 255240 159798 255268 163200
rect 255228 159792 255280 159798
rect 255228 159734 255280 159740
rect 254400 158772 254452 158778
rect 254400 158714 254452 158720
rect 255412 158772 255464 158778
rect 255412 158714 255464 158720
rect 255320 158568 255372 158574
rect 255320 158510 255372 158516
rect 254032 155712 254084 155718
rect 254032 155654 254084 155660
rect 254044 150226 254072 155654
rect 255332 150226 255360 158510
rect 255424 152386 255452 158714
rect 255872 155576 255924 155582
rect 255872 155518 255924 155524
rect 255412 152380 255464 152386
rect 255412 152322 255464 152328
rect 255884 151814 255912 155518
rect 256068 153406 256096 163200
rect 256792 158704 256844 158710
rect 256792 158646 256844 158652
rect 256516 153536 256568 153542
rect 256516 153478 256568 153484
rect 256056 153400 256108 153406
rect 256056 153342 256108 153348
rect 256528 151814 256556 153478
rect 255884 151786 256004 151814
rect 256528 151786 256648 151814
rect 255976 150226 256004 151786
rect 256620 150226 256648 151786
rect 248282 150146 248334 150152
rect 248294 149940 248322 150146
rect 248938 149940 248966 150198
rect 249582 149940 249610 150198
rect 250226 149940 250254 150198
rect 250870 149940 250898 150198
rect 251514 149940 251542 150198
rect 252158 149940 252186 150198
rect 252802 149940 252830 150198
rect 253446 149940 253474 150198
rect 253940 150204 253992 150210
rect 254044 150198 254118 150226
rect 253940 150146 253992 150152
rect 254090 149940 254118 150198
rect 254722 150204 254774 150210
rect 255332 150198 255406 150226
rect 255976 150198 256050 150226
rect 256620 150198 256694 150226
rect 256804 150210 256832 158646
rect 256896 158234 256924 163200
rect 256884 158228 256936 158234
rect 256884 158170 256936 158176
rect 257724 153066 257752 163200
rect 258552 158778 258580 163200
rect 259472 161474 259500 163200
rect 259472 161446 259592 161474
rect 258540 158772 258592 158778
rect 258540 158714 258592 158720
rect 259460 157956 259512 157962
rect 259460 157898 259512 157904
rect 258080 157548 258132 157554
rect 258080 157490 258132 157496
rect 257252 153060 257304 153066
rect 257252 153002 257304 153008
rect 257712 153060 257764 153066
rect 257712 153002 257764 153008
rect 257264 150226 257292 153002
rect 254722 150146 254774 150152
rect 254734 149940 254762 150146
rect 255378 149940 255406 150198
rect 256022 149940 256050 150198
rect 256666 149940 256694 150198
rect 256792 150204 256844 150210
rect 257264 150198 257338 150226
rect 258092 150210 258120 157490
rect 258540 154284 258592 154290
rect 258540 154226 258592 154232
rect 258552 150226 258580 154226
rect 256792 150146 256844 150152
rect 257310 149940 257338 150198
rect 257942 150204 257994 150210
rect 257942 150146 257994 150152
rect 258080 150204 258132 150210
rect 258552 150198 258626 150226
rect 259472 150210 259500 157898
rect 259564 153406 259592 161446
rect 259828 159860 259880 159866
rect 259828 159802 259880 159808
rect 259552 153400 259604 153406
rect 259552 153342 259604 153348
rect 259840 150226 259868 159802
rect 260300 155514 260328 163200
rect 261128 158846 261156 163200
rect 261956 159866 261984 163200
rect 261944 159860 261996 159866
rect 261944 159802 261996 159808
rect 261116 158840 261168 158846
rect 261116 158782 261168 158788
rect 261024 158772 261076 158778
rect 261024 158714 261076 158720
rect 260840 155780 260892 155786
rect 260840 155722 260892 155728
rect 260288 155508 260340 155514
rect 260288 155450 260340 155456
rect 260852 151814 260880 155722
rect 261036 151842 261064 158714
rect 261392 155372 261444 155378
rect 261392 155314 261444 155320
rect 261024 151836 261076 151842
rect 260852 151786 260972 151814
rect 260944 150226 260972 151786
rect 261404 151814 261432 155314
rect 262784 153474 262812 163200
rect 263048 157888 263100 157894
rect 263048 157830 263100 157836
rect 262772 153468 262824 153474
rect 262772 153410 262824 153416
rect 262404 152924 262456 152930
rect 262404 152866 262456 152872
rect 261404 151786 261800 151814
rect 261024 151778 261076 151784
rect 261772 150226 261800 151786
rect 262416 150226 262444 152866
rect 263060 150226 263088 157830
rect 263612 155582 263640 163200
rect 264440 158778 264468 163200
rect 264888 159928 264940 159934
rect 264888 159870 264940 159876
rect 264428 158772 264480 158778
rect 264428 158714 264480 158720
rect 263784 157752 263836 157758
rect 263784 157694 263836 157700
rect 263692 155916 263744 155922
rect 263692 155858 263744 155864
rect 263600 155576 263652 155582
rect 263600 155518 263652 155524
rect 263600 155372 263652 155378
rect 263600 155314 263652 155320
rect 258080 150146 258132 150152
rect 257954 149940 257982 150146
rect 258598 149940 258626 150198
rect 259230 150204 259282 150210
rect 259230 150146 259282 150152
rect 259460 150204 259512 150210
rect 259840 150198 259914 150226
rect 259460 150146 259512 150152
rect 259242 149940 259270 150146
rect 259886 149940 259914 150198
rect 260518 150204 260570 150210
rect 260944 150198 261202 150226
rect 261772 150198 261846 150226
rect 262416 150198 262490 150226
rect 263060 150198 263134 150226
rect 263612 150210 263640 155314
rect 263704 150226 263732 155858
rect 263796 155378 263824 157694
rect 263784 155372 263836 155378
rect 263784 155314 263836 155320
rect 264900 151814 264928 159870
rect 265164 157276 265216 157282
rect 265164 157218 265216 157224
rect 265176 151814 265204 157218
rect 265360 152318 265388 163200
rect 266084 155168 266136 155174
rect 266084 155110 266136 155116
rect 265348 152312 265400 152318
rect 265348 152254 265400 152260
rect 266096 151814 266124 155110
rect 266188 154290 266216 163200
rect 266912 156188 266964 156194
rect 266912 156130 266964 156136
rect 266176 154284 266228 154290
rect 266176 154226 266228 154232
rect 264900 151786 265020 151814
rect 265176 151786 265664 151814
rect 266096 151786 266308 151814
rect 264992 150226 265020 151786
rect 265636 150226 265664 151786
rect 266280 150226 266308 151786
rect 266924 150226 266952 156130
rect 267016 155650 267044 163200
rect 267844 158778 267872 163200
rect 268672 159934 268700 163200
rect 268660 159928 268712 159934
rect 268660 159870 268712 159876
rect 267648 158772 267700 158778
rect 267648 158714 267700 158720
rect 267832 158772 267884 158778
rect 267832 158714 267884 158720
rect 267004 155644 267056 155650
rect 267004 155586 267056 155592
rect 267660 152998 267688 158714
rect 267740 157820 267792 157826
rect 267740 157762 267792 157768
rect 267556 152992 267608 152998
rect 267556 152934 267608 152940
rect 267648 152992 267700 152998
rect 267648 152934 267700 152940
rect 267568 150226 267596 152934
rect 267752 151814 267780 157762
rect 269212 156256 269264 156262
rect 269212 156198 269264 156204
rect 268844 155100 268896 155106
rect 268844 155042 268896 155048
rect 267752 151786 268240 151814
rect 268212 150226 268240 151786
rect 268856 150226 268884 155042
rect 269224 151814 269252 156198
rect 269500 153270 269528 163200
rect 270132 159996 270184 160002
rect 270132 159938 270184 159944
rect 269488 153264 269540 153270
rect 269488 153206 269540 153212
rect 269224 151786 269528 151814
rect 269500 150226 269528 151786
rect 270144 150226 270172 159938
rect 270328 157010 270356 163200
rect 271248 160002 271276 163200
rect 272076 163146 272104 163200
rect 272168 163146 272196 163254
rect 272076 163118 272196 163146
rect 271236 159996 271288 160002
rect 271236 159938 271288 159944
rect 270316 157004 270368 157010
rect 270316 156946 270368 156952
rect 270500 156596 270552 156602
rect 270500 156538 270552 156544
rect 270512 151814 270540 156538
rect 272064 156120 272116 156126
rect 272064 156062 272116 156068
rect 271420 155032 271472 155038
rect 271420 154974 271472 154980
rect 270868 152924 270920 152930
rect 270868 152866 270920 152872
rect 270880 152318 270908 152866
rect 270868 152312 270920 152318
rect 270868 152254 270920 152260
rect 270512 151786 270816 151814
rect 270788 150226 270816 151786
rect 271432 150226 271460 154974
rect 272076 150226 272104 156062
rect 272524 152312 272576 152318
rect 272524 152254 272576 152260
rect 272536 151842 272564 152254
rect 272628 151910 272656 163254
rect 272890 163200 272946 164400
rect 273718 163200 273774 164400
rect 274546 163200 274602 164400
rect 275374 163200 275430 164400
rect 276202 163200 276258 164400
rect 277122 163200 277178 164400
rect 277950 163200 278006 164400
rect 278778 163200 278834 164400
rect 279606 163200 279662 164400
rect 279712 163254 280016 163282
rect 272800 159996 272852 160002
rect 272800 159938 272852 159944
rect 272812 152114 272840 159938
rect 272904 153338 272932 163200
rect 273260 157344 273312 157350
rect 273260 157286 273312 157292
rect 272892 153332 272944 153338
rect 272892 153274 272944 153280
rect 272708 152108 272760 152114
rect 272708 152050 272760 152056
rect 272800 152108 272852 152114
rect 272800 152050 272852 152056
rect 272616 151904 272668 151910
rect 272616 151846 272668 151852
rect 272524 151836 272576 151842
rect 272524 151778 272576 151784
rect 272720 150226 272748 152050
rect 273272 150226 273300 157286
rect 273732 157146 273760 163200
rect 274560 159497 274588 163200
rect 275388 160002 275416 163200
rect 275376 159996 275428 160002
rect 275376 159938 275428 159944
rect 274546 159488 274602 159497
rect 274546 159423 274602 159432
rect 275190 159352 275246 159361
rect 275190 159287 275246 159296
rect 273720 157140 273772 157146
rect 273720 157082 273772 157088
rect 273904 156528 273956 156534
rect 273904 156470 273956 156476
rect 273916 150226 273944 156470
rect 274548 152176 274600 152182
rect 274548 152118 274600 152124
rect 274560 150226 274588 152118
rect 275204 150226 275232 159287
rect 276020 155848 276072 155854
rect 276020 155790 276072 155796
rect 275836 154352 275888 154358
rect 275836 154294 275888 154300
rect 275848 150226 275876 154294
rect 276032 151814 276060 155790
rect 276216 154358 276244 163200
rect 277136 157078 277164 163200
rect 277124 157072 277176 157078
rect 277124 157014 277176 157020
rect 277124 154896 277176 154902
rect 277124 154838 277176 154844
rect 276204 154352 276256 154358
rect 276204 154294 276256 154300
rect 276032 151786 276520 151814
rect 276492 150226 276520 151786
rect 277136 150226 277164 154838
rect 277768 152516 277820 152522
rect 277768 152458 277820 152464
rect 277780 150226 277808 152458
rect 277964 152182 277992 163200
rect 278792 159118 278820 163200
rect 279620 163146 279648 163200
rect 279712 163146 279740 163254
rect 279620 163118 279740 163146
rect 278688 159112 278740 159118
rect 278686 159080 278688 159089
rect 278780 159112 278832 159118
rect 278740 159080 278742 159089
rect 278780 159054 278832 159060
rect 279884 159112 279936 159118
rect 279884 159054 279936 159060
rect 278686 159015 278742 159024
rect 279056 156460 279108 156466
rect 279056 156402 279108 156408
rect 278412 154420 278464 154426
rect 278412 154362 278464 154368
rect 277952 152176 278004 152182
rect 277952 152118 278004 152124
rect 278424 150226 278452 154362
rect 279068 150226 279096 156402
rect 279896 153134 279924 159054
rect 279988 154426 280016 163254
rect 280434 163200 280490 164400
rect 281262 163200 281318 164400
rect 282090 163200 282146 164400
rect 283010 163200 283066 164400
rect 283838 163200 283894 164400
rect 284666 163200 284722 164400
rect 285494 163200 285550 164400
rect 286322 163200 286378 164400
rect 287150 163200 287206 164400
rect 287978 163200 288034 164400
rect 288898 163200 288954 164400
rect 289726 163200 289782 164400
rect 290554 163200 290610 164400
rect 291382 163200 291438 164400
rect 292210 163200 292266 164400
rect 292316 163254 292528 163282
rect 280344 160064 280396 160070
rect 280344 160006 280396 160012
rect 280068 159112 280120 159118
rect 280066 159080 280068 159089
rect 280120 159080 280122 159089
rect 280066 159015 280122 159024
rect 279976 154420 280028 154426
rect 279976 154362 280028 154368
rect 279700 153128 279752 153134
rect 279700 153070 279752 153076
rect 279884 153128 279936 153134
rect 279884 153070 279936 153076
rect 279712 150226 279740 153070
rect 280356 150226 280384 160006
rect 280448 157214 280476 163200
rect 281276 160070 281304 163200
rect 281264 160064 281316 160070
rect 281264 160006 281316 160012
rect 282104 159322 282132 163200
rect 281540 159316 281592 159322
rect 281540 159258 281592 159264
rect 282092 159316 282144 159322
rect 282092 159258 282144 159264
rect 280436 157208 280488 157214
rect 280436 157150 280488 157156
rect 280986 153776 281042 153785
rect 280986 153711 281042 153720
rect 281000 150226 281028 153711
rect 260518 150146 260570 150152
rect 260530 149940 260558 150146
rect 261174 149940 261202 150198
rect 261818 149940 261846 150198
rect 262462 149940 262490 150198
rect 263106 149940 263134 150198
rect 263600 150204 263652 150210
rect 263704 150198 263778 150226
rect 263600 150146 263652 150152
rect 263750 149940 263778 150198
rect 264382 150204 264434 150210
rect 264992 150198 265066 150226
rect 265636 150198 265710 150226
rect 266280 150198 266354 150226
rect 266924 150198 266998 150226
rect 267568 150198 267642 150226
rect 268212 150198 268286 150226
rect 268856 150198 268930 150226
rect 269500 150198 269574 150226
rect 270144 150198 270218 150226
rect 270788 150198 270862 150226
rect 271432 150198 271506 150226
rect 272076 150198 272150 150226
rect 272720 150198 272794 150226
rect 273272 150198 273346 150226
rect 273916 150198 273990 150226
rect 274560 150198 274634 150226
rect 275204 150198 275278 150226
rect 275848 150198 275922 150226
rect 276492 150198 276566 150226
rect 277136 150198 277210 150226
rect 277780 150198 277854 150226
rect 278424 150198 278498 150226
rect 279068 150198 279142 150226
rect 279712 150198 279786 150226
rect 280356 150198 280430 150226
rect 281000 150198 281074 150226
rect 281552 150210 281580 159258
rect 283024 159118 283052 163200
rect 282920 159112 282972 159118
rect 282920 159054 282972 159060
rect 283012 159112 283064 159118
rect 283012 159054 283064 159060
rect 282932 158930 282960 159054
rect 282932 158902 283052 158930
rect 281632 156664 281684 156670
rect 281632 156606 281684 156612
rect 281644 150226 281672 156606
rect 282920 152244 282972 152250
rect 282920 152186 282972 152192
rect 282932 150226 282960 152186
rect 283024 151842 283052 158902
rect 283852 156670 283880 163200
rect 284680 159118 284708 163200
rect 285404 159248 285456 159254
rect 285404 159190 285456 159196
rect 284208 159112 284260 159118
rect 284208 159054 284260 159060
rect 284668 159112 284720 159118
rect 284668 159054 284720 159060
rect 283840 156664 283892 156670
rect 283840 156606 283892 156612
rect 283104 156392 283156 156398
rect 283104 156334 283156 156340
rect 283012 151836 283064 151842
rect 283012 151778 283064 151784
rect 264382 150146 264434 150152
rect 264394 149940 264422 150146
rect 265038 149940 265066 150198
rect 265682 149940 265710 150198
rect 266326 149940 266354 150198
rect 266970 149940 266998 150198
rect 267614 149940 267642 150198
rect 268258 149940 268286 150198
rect 268902 149940 268930 150198
rect 269546 149940 269574 150198
rect 270190 149940 270218 150198
rect 270834 149940 270862 150198
rect 271478 149940 271506 150198
rect 272122 149940 272150 150198
rect 272766 149940 272794 150198
rect 273318 149940 273346 150198
rect 273962 149940 273990 150198
rect 274606 149940 274634 150198
rect 275250 149940 275278 150198
rect 275894 149940 275922 150198
rect 276538 149940 276566 150198
rect 277182 149940 277210 150198
rect 277826 149940 277854 150198
rect 278470 149940 278498 150198
rect 279114 149940 279142 150198
rect 279758 149940 279786 150198
rect 280402 149940 280430 150198
rect 281046 149940 281074 150198
rect 281540 150204 281592 150210
rect 281644 150198 281718 150226
rect 281540 150146 281592 150152
rect 281690 149940 281718 150198
rect 282322 150204 282374 150210
rect 282932 150198 283006 150226
rect 283116 150210 283144 156334
rect 284220 153950 284248 159054
rect 283656 153944 283708 153950
rect 283656 153886 283708 153892
rect 284208 153944 284260 153950
rect 284208 153886 284260 153892
rect 283668 150226 283696 153886
rect 284852 152652 284904 152658
rect 284852 152594 284904 152600
rect 282322 150146 282374 150152
rect 282334 149940 282362 150146
rect 282978 149940 283006 150198
rect 283104 150204 283156 150210
rect 283104 150146 283156 150152
rect 283622 150198 283696 150226
rect 284864 150226 284892 152594
rect 285416 151814 285444 159190
rect 285508 152250 285536 163200
rect 285864 159112 285916 159118
rect 285864 159054 285916 159060
rect 285680 156800 285732 156806
rect 285680 156742 285732 156748
rect 285496 152244 285548 152250
rect 285496 152186 285548 152192
rect 285416 151786 285536 151814
rect 285508 150226 285536 151786
rect 284254 150204 284306 150210
rect 283622 149940 283650 150198
rect 284864 150198 284938 150226
rect 285508 150198 285582 150226
rect 285692 150210 285720 156742
rect 285876 152522 285904 159054
rect 286336 153882 286364 163200
rect 287164 156806 287192 163200
rect 287992 159254 288020 163200
rect 287980 159248 288032 159254
rect 287980 159190 288032 159196
rect 288912 159186 288940 163200
rect 288348 159180 288400 159186
rect 288348 159122 288400 159128
rect 288900 159180 288952 159186
rect 288900 159122 288952 159128
rect 287152 156800 287204 156806
rect 287152 156742 287204 156748
rect 286140 153876 286192 153882
rect 286140 153818 286192 153824
rect 286324 153876 286376 153882
rect 286324 153818 286376 153824
rect 285864 152516 285916 152522
rect 285864 152458 285916 152464
rect 286152 150226 286180 153818
rect 288360 152726 288388 159122
rect 289360 156732 289412 156738
rect 289360 156674 289412 156680
rect 288716 153808 288768 153814
rect 288716 153750 288768 153756
rect 288072 152720 288124 152726
rect 288072 152662 288124 152668
rect 288348 152720 288400 152726
rect 288348 152662 288400 152668
rect 287428 151836 287480 151842
rect 287428 151778 287480 151784
rect 287440 150226 287468 151778
rect 288084 150226 288112 152662
rect 288728 150226 288756 153750
rect 289372 150226 289400 156674
rect 289740 155718 289768 163200
rect 290568 157282 290596 163200
rect 290648 159384 290700 159390
rect 290648 159326 290700 159332
rect 290556 157276 290608 157282
rect 290556 157218 290608 157224
rect 289728 155712 289780 155718
rect 289728 155654 289780 155660
rect 290004 152720 290056 152726
rect 290004 152662 290056 152668
rect 290016 150226 290044 152662
rect 290660 150226 290688 159326
rect 291292 154488 291344 154494
rect 291292 154430 291344 154436
rect 291304 150226 291332 154430
rect 291396 152726 291424 163200
rect 292224 163146 292252 163200
rect 292316 163146 292344 163254
rect 292224 163118 292344 163146
rect 291936 156936 291988 156942
rect 291936 156878 291988 156884
rect 291384 152720 291436 152726
rect 291384 152662 291436 152668
rect 291844 152516 291896 152522
rect 291844 152458 291896 152464
rect 291856 152250 291884 152458
rect 291844 152244 291896 152250
rect 291844 152186 291896 152192
rect 291948 150226 291976 156878
rect 292500 152250 292528 163254
rect 293038 163200 293094 164400
rect 293866 163200 293922 164400
rect 294786 163200 294842 164400
rect 295614 163200 295670 164400
rect 296442 163200 296498 164400
rect 297270 163200 297326 164400
rect 298098 163200 298154 164400
rect 298926 163200 298982 164400
rect 299032 163254 299428 163282
rect 293052 155854 293080 163200
rect 293880 156738 293908 163200
rect 294800 159390 294828 163200
rect 295628 159526 295656 163200
rect 295524 159520 295576 159526
rect 295524 159462 295576 159468
rect 295616 159520 295668 159526
rect 295616 159462 295668 159468
rect 294788 159384 294840 159390
rect 294788 159326 294840 159332
rect 295156 159044 295208 159050
rect 295156 158986 295208 158992
rect 294052 156868 294104 156874
rect 294052 156810 294104 156816
rect 293868 156732 293920 156738
rect 293868 156674 293920 156680
rect 293040 155848 293092 155854
rect 293040 155790 293092 155796
rect 293868 153740 293920 153746
rect 293868 153682 293920 153688
rect 293224 152652 293276 152658
rect 293224 152594 293276 152600
rect 292578 152416 292634 152425
rect 292578 152351 292634 152360
rect 292488 152244 292540 152250
rect 292488 152186 292540 152192
rect 292592 150226 292620 152351
rect 293236 150226 293264 152594
rect 293880 150226 293908 153682
rect 294064 151814 294092 156810
rect 294064 151786 294552 151814
rect 294524 150226 294552 151786
rect 295168 150226 295196 158986
rect 295536 151814 295564 159462
rect 296456 155786 296484 163200
rect 297088 158092 297140 158098
rect 297088 158034 297140 158040
rect 296444 155780 296496 155786
rect 296444 155722 296496 155728
rect 296444 154556 296496 154562
rect 296444 154498 296496 154504
rect 295536 151786 295840 151814
rect 295812 150226 295840 151786
rect 296456 150226 296484 154498
rect 297100 150226 297128 158034
rect 297284 156874 297312 163200
rect 298008 159452 298060 159458
rect 298008 159394 298060 159400
rect 297272 156868 297324 156874
rect 297272 156810 297324 156816
rect 297732 153196 297784 153202
rect 297732 153138 297784 153144
rect 297744 150226 297772 153138
rect 298020 151814 298048 159394
rect 298112 158914 298140 163200
rect 298940 163146 298968 163200
rect 299032 163146 299060 163254
rect 298940 163118 299060 163146
rect 298100 158908 298152 158914
rect 298100 158850 298152 158856
rect 299020 154012 299072 154018
rect 299020 153954 299072 153960
rect 298020 151786 298416 151814
rect 298388 150226 298416 151786
rect 299032 150226 299060 153954
rect 299400 152590 299428 163254
rect 299754 163200 299810 164400
rect 300674 163200 300730 164400
rect 301502 163200 301558 164400
rect 302330 163200 302386 164400
rect 303158 163200 303214 164400
rect 303986 163200 304042 164400
rect 304814 163200 304870 164400
rect 305642 163200 305698 164400
rect 306562 163200 306618 164400
rect 307390 163200 307446 164400
rect 308218 163200 308274 164400
rect 309046 163200 309102 164400
rect 309874 163200 309930 164400
rect 310702 163200 310758 164400
rect 311530 163200 311586 164400
rect 311636 163254 311848 163282
rect 299480 159044 299532 159050
rect 299480 158986 299532 158992
rect 299388 152584 299440 152590
rect 299388 152526 299440 152532
rect 284254 150146 284306 150152
rect 284266 149940 284294 150146
rect 284910 149940 284938 150198
rect 285554 149940 285582 150198
rect 285680 150204 285732 150210
rect 286152 150198 286226 150226
rect 285680 150146 285732 150152
rect 286198 149940 286226 150198
rect 286830 150204 286882 150210
rect 287440 150198 287514 150226
rect 288084 150198 288158 150226
rect 288728 150198 288802 150226
rect 289372 150198 289446 150226
rect 290016 150198 290090 150226
rect 290660 150198 290734 150226
rect 291304 150198 291378 150226
rect 291948 150198 292022 150226
rect 292592 150198 292666 150226
rect 293236 150198 293310 150226
rect 293880 150198 293954 150226
rect 294524 150198 294598 150226
rect 295168 150198 295242 150226
rect 295812 150198 295886 150226
rect 296456 150198 296530 150226
rect 297100 150198 297174 150226
rect 297744 150198 297818 150226
rect 298388 150198 298462 150226
rect 299032 150198 299106 150226
rect 299492 150210 299520 158986
rect 299768 155242 299796 163200
rect 300308 158908 300360 158914
rect 300308 158850 300360 158856
rect 299664 155236 299716 155242
rect 299664 155178 299716 155184
rect 299756 155236 299808 155242
rect 299756 155178 299808 155184
rect 299676 150226 299704 155178
rect 300320 153202 300348 158850
rect 300688 158098 300716 163200
rect 301516 159458 301544 163200
rect 301504 159452 301556 159458
rect 301504 159394 301556 159400
rect 302344 159118 302372 163200
rect 302424 159656 302476 159662
rect 302424 159598 302476 159604
rect 302332 159112 302384 159118
rect 302332 159054 302384 159060
rect 300676 158092 300728 158098
rect 300676 158034 300728 158040
rect 302240 158024 302292 158030
rect 302240 157966 302292 157972
rect 301596 153672 301648 153678
rect 301596 153614 301648 153620
rect 300308 153196 300360 153202
rect 300308 153138 300360 153144
rect 300952 152040 301004 152046
rect 300952 151982 301004 151988
rect 300964 150226 300992 151982
rect 301608 150226 301636 153614
rect 302252 150226 302280 157966
rect 286830 150146 286882 150152
rect 286842 149940 286870 150146
rect 287486 149940 287514 150198
rect 288130 149940 288158 150198
rect 288774 149940 288802 150198
rect 289418 149940 289446 150198
rect 290062 149940 290090 150198
rect 290706 149940 290734 150198
rect 291350 149940 291378 150198
rect 291994 149940 292022 150198
rect 292638 149940 292666 150198
rect 293282 149940 293310 150198
rect 293926 149940 293954 150198
rect 294570 149940 294598 150198
rect 295214 149940 295242 150198
rect 295858 149940 295886 150198
rect 296502 149940 296530 150198
rect 297146 149940 297174 150198
rect 297790 149940 297818 150198
rect 298434 149940 298462 150198
rect 299078 149940 299106 150198
rect 299480 150204 299532 150210
rect 299676 150198 299750 150226
rect 299480 150146 299532 150152
rect 299722 149940 299750 150198
rect 300354 150204 300406 150210
rect 300964 150198 301038 150226
rect 301608 150198 301682 150226
rect 302252 150198 302326 150226
rect 302436 150210 302464 159598
rect 303172 155922 303200 163200
rect 303160 155916 303212 155922
rect 303160 155858 303212 155864
rect 302884 151972 302936 151978
rect 302884 151914 302936 151920
rect 302896 150226 302924 151914
rect 304000 151842 304028 163200
rect 304724 155304 304776 155310
rect 304724 155246 304776 155252
rect 304080 154080 304132 154086
rect 304080 154022 304132 154028
rect 303988 151836 304040 151842
rect 303988 151778 304040 151784
rect 304092 150226 304120 154022
rect 304736 150226 304764 155246
rect 304828 152046 304856 163200
rect 305368 158976 305420 158982
rect 305368 158918 305420 158924
rect 304816 152040 304868 152046
rect 304816 151982 304868 151988
rect 305380 150226 305408 158918
rect 305656 158914 305684 163200
rect 305644 158908 305696 158914
rect 305644 158850 305696 158856
rect 306576 155174 306604 163200
rect 307404 159050 307432 163200
rect 308232 159730 308260 163200
rect 308220 159724 308272 159730
rect 308220 159666 308272 159672
rect 309060 159662 309088 163200
rect 309888 161474 309916 163200
rect 309888 161446 310008 161474
rect 308588 159656 308640 159662
rect 308588 159598 308640 159604
rect 309048 159656 309100 159662
rect 309048 159598 309100 159604
rect 307392 159044 307444 159050
rect 307392 158986 307444 158992
rect 307300 158908 307352 158914
rect 307300 158850 307352 158856
rect 306932 158160 306984 158166
rect 306932 158102 306984 158108
rect 306564 155168 306616 155174
rect 306564 155110 306616 155116
rect 306656 154148 306708 154154
rect 306656 154090 306708 154096
rect 306012 152448 306064 152454
rect 306012 152390 306064 152396
rect 306024 150226 306052 152390
rect 306668 150226 306696 154090
rect 306944 151814 306972 158102
rect 307312 152454 307340 158850
rect 307944 152788 307996 152794
rect 307944 152730 307996 152736
rect 307300 152448 307352 152454
rect 307300 152390 307352 152396
rect 306944 151786 307340 151814
rect 307312 150226 307340 151786
rect 307956 150226 307984 152730
rect 308600 150226 308628 159598
rect 309876 155440 309928 155446
rect 309876 155382 309928 155388
rect 309232 153604 309284 153610
rect 309232 153546 309284 153552
rect 309244 150226 309272 153546
rect 309888 150226 309916 155382
rect 309980 155310 310008 161446
rect 310612 159588 310664 159594
rect 310612 159530 310664 159536
rect 309968 155304 310020 155310
rect 309968 155246 310020 155252
rect 310624 150226 310652 159530
rect 310716 158982 310744 163200
rect 311544 163146 311572 163200
rect 311636 163146 311664 163254
rect 311544 163118 311664 163146
rect 310704 158976 310756 158982
rect 310704 158918 310756 158924
rect 311716 154216 311768 154222
rect 311716 154158 311768 154164
rect 311164 152856 311216 152862
rect 311164 152798 311216 152804
rect 300354 150146 300406 150152
rect 300366 149940 300394 150146
rect 301010 149940 301038 150198
rect 301654 149940 301682 150198
rect 302298 149940 302326 150198
rect 302424 150204 302476 150210
rect 302896 150198 302970 150226
rect 302424 150146 302476 150152
rect 302942 149940 302970 150198
rect 303574 150204 303626 150210
rect 304092 150198 304166 150226
rect 304736 150198 304810 150226
rect 305380 150198 305454 150226
rect 306024 150198 306098 150226
rect 306668 150198 306742 150226
rect 307312 150198 307386 150226
rect 307956 150198 308030 150226
rect 308600 150198 308674 150226
rect 309244 150198 309318 150226
rect 309888 150198 309962 150226
rect 303574 150146 303626 150152
rect 303586 149940 303614 150146
rect 304138 149940 304166 150198
rect 304782 149940 304810 150198
rect 305426 149940 305454 150198
rect 306070 149940 306098 150198
rect 306714 149940 306742 150198
rect 307358 149940 307386 150198
rect 308002 149940 308030 150198
rect 308646 149940 308674 150198
rect 309290 149940 309318 150198
rect 309934 149940 309962 150198
rect 310578 150198 310652 150226
rect 311176 150226 311204 152798
rect 311728 151814 311756 154158
rect 311820 152794 311848 163254
rect 312450 163200 312506 164400
rect 313278 163200 313334 164400
rect 314106 163200 314162 164400
rect 314934 163200 314990 164400
rect 315762 163200 315818 164400
rect 316590 163200 316646 164400
rect 317418 163200 317474 164400
rect 318338 163200 318394 164400
rect 318444 163254 318748 163282
rect 312464 158914 312492 163200
rect 313188 158976 313240 158982
rect 313188 158918 313240 158924
rect 312452 158908 312504 158914
rect 312452 158850 312504 158856
rect 312452 154964 312504 154970
rect 312452 154906 312504 154912
rect 311808 152788 311860 152794
rect 311808 152730 311860 152736
rect 311728 151786 311848 151814
rect 311820 150226 311848 151786
rect 312464 150226 312492 154906
rect 313200 152386 313228 158918
rect 313292 154018 313320 163200
rect 314120 159798 314148 163200
rect 313740 159792 313792 159798
rect 313740 159734 313792 159740
rect 314108 159792 314160 159798
rect 314108 159734 314160 159740
rect 313464 158908 313516 158914
rect 313464 158850 313516 158856
rect 313280 154012 313332 154018
rect 313280 153954 313332 153960
rect 313476 152425 313504 158850
rect 313462 152416 313518 152425
rect 313096 152380 313148 152386
rect 313096 152322 313148 152328
rect 313188 152380 313240 152386
rect 313462 152351 313518 152360
rect 313188 152322 313240 152328
rect 313108 150226 313136 152322
rect 313752 150226 313780 159734
rect 314948 158982 314976 163200
rect 315776 159594 315804 163200
rect 315764 159588 315816 159594
rect 315764 159530 315816 159536
rect 314936 158976 314988 158982
rect 314936 158918 314988 158924
rect 315028 158228 315080 158234
rect 315028 158170 315080 158176
rect 314384 153536 314436 153542
rect 314384 153478 314436 153484
rect 314396 150226 314424 153478
rect 315040 150226 315068 158170
rect 316604 155378 316632 163200
rect 317432 158846 317460 163200
rect 318352 163146 318380 163200
rect 318444 163146 318472 163254
rect 318352 163118 318472 163146
rect 317144 158840 317196 158846
rect 317144 158782 317196 158788
rect 317420 158840 317472 158846
rect 317420 158782 317472 158788
rect 318432 158840 318484 158846
rect 318432 158782 318484 158788
rect 316592 155372 316644 155378
rect 316592 155314 316644 155320
rect 316960 153400 317012 153406
rect 316960 153342 317012 153348
rect 315672 153060 315724 153066
rect 315672 153002 315724 153008
rect 315684 150226 315712 153002
rect 316316 152312 316368 152318
rect 316316 152254 316368 152260
rect 316328 150226 316356 152254
rect 316972 150226 317000 153342
rect 317156 153066 317184 158782
rect 317604 155508 317656 155514
rect 317604 155450 317656 155456
rect 317144 153060 317196 153066
rect 317144 153002 317196 153008
rect 317616 150226 317644 155450
rect 318444 153066 318472 158782
rect 318248 153060 318300 153066
rect 318248 153002 318300 153008
rect 318432 153060 318484 153066
rect 318432 153002 318484 153008
rect 318260 150226 318288 153002
rect 318720 152862 318748 163254
rect 319166 163200 319222 164400
rect 319994 163200 320050 164400
rect 320822 163200 320878 164400
rect 321650 163200 321706 164400
rect 322478 163200 322534 164400
rect 323306 163200 323362 164400
rect 324226 163200 324282 164400
rect 325054 163200 325110 164400
rect 325882 163200 325938 164400
rect 326710 163200 326766 164400
rect 327538 163200 327594 164400
rect 328366 163200 328422 164400
rect 329194 163200 329250 164400
rect 330114 163200 330170 164400
rect 330942 163200 330998 164400
rect 331770 163200 331826 164400
rect 332598 163200 332654 164400
rect 333426 163200 333482 164400
rect 334254 163200 334310 164400
rect 335082 163200 335138 164400
rect 336002 163200 336058 164400
rect 336108 163254 336320 163282
rect 318984 159860 319036 159866
rect 318984 159802 319036 159808
rect 318708 152856 318760 152862
rect 318708 152798 318760 152804
rect 318996 150226 319024 159802
rect 319180 158846 319208 163200
rect 319168 158840 319220 158846
rect 319168 158782 319220 158788
rect 320008 154086 320036 163200
rect 320836 159866 320864 163200
rect 320824 159860 320876 159866
rect 320824 159802 320876 159808
rect 321560 158840 321612 158846
rect 321560 158782 321612 158788
rect 320272 158772 320324 158778
rect 320272 158714 320324 158720
rect 320180 155576 320232 155582
rect 320180 155518 320232 155524
rect 319996 154080 320048 154086
rect 319996 154022 320048 154028
rect 319536 153468 319588 153474
rect 319536 153410 319588 153416
rect 311176 150198 311250 150226
rect 311820 150198 311894 150226
rect 312464 150198 312538 150226
rect 313108 150198 313182 150226
rect 313752 150198 313826 150226
rect 314396 150198 314470 150226
rect 315040 150198 315114 150226
rect 315684 150198 315758 150226
rect 316328 150198 316402 150226
rect 316972 150198 317046 150226
rect 317616 150198 317690 150226
rect 318260 150198 318334 150226
rect 310578 149940 310606 150198
rect 311222 149940 311250 150198
rect 311866 149940 311894 150198
rect 312510 149940 312538 150198
rect 313154 149940 313182 150198
rect 313798 149940 313826 150198
rect 314442 149940 314470 150198
rect 315086 149940 315114 150198
rect 315730 149940 315758 150198
rect 316374 149940 316402 150198
rect 317018 149940 317046 150198
rect 317662 149940 317690 150198
rect 318306 149940 318334 150198
rect 318950 150198 319024 150226
rect 319548 150226 319576 153410
rect 320192 150226 320220 155518
rect 320284 152318 320312 158714
rect 320916 152992 320968 152998
rect 320916 152934 320968 152940
rect 320272 152312 320324 152318
rect 320272 152254 320324 152260
rect 320928 150226 320956 152934
rect 321572 152930 321600 158782
rect 321664 158778 321692 163200
rect 322492 158846 322520 163200
rect 322480 158840 322532 158846
rect 322480 158782 322532 158788
rect 321652 158772 321704 158778
rect 321652 158714 321704 158720
rect 322112 155644 322164 155650
rect 322112 155586 322164 155592
rect 322020 154284 322072 154290
rect 322020 154226 322072 154232
rect 321468 152924 321520 152930
rect 321468 152866 321520 152872
rect 321560 152924 321612 152930
rect 321560 152866 321612 152872
rect 319548 150198 319622 150226
rect 320192 150198 320266 150226
rect 318950 149940 318978 150198
rect 319594 149940 319622 150198
rect 320238 149940 320266 150198
rect 320882 150198 320956 150226
rect 321480 150226 321508 152866
rect 322032 150498 322060 154226
rect 322124 151814 322152 155586
rect 323320 154154 323348 163200
rect 324044 159928 324096 159934
rect 324044 159870 324096 159876
rect 323308 154148 323360 154154
rect 323308 154090 323360 154096
rect 323492 152924 323544 152930
rect 323492 152866 323544 152872
rect 323504 152318 323532 152866
rect 323400 152312 323452 152318
rect 323400 152254 323452 152260
rect 323492 152312 323544 152318
rect 323492 152254 323544 152260
rect 322124 151786 322796 151814
rect 322032 150470 322152 150498
rect 322124 150226 322152 150470
rect 322768 150226 322796 151786
rect 323412 150226 323440 152254
rect 324056 150226 324084 159870
rect 324240 152930 324268 163200
rect 324688 153264 324740 153270
rect 324688 153206 324740 153212
rect 324228 152924 324280 152930
rect 324228 152866 324280 152872
rect 324700 150226 324728 153206
rect 325068 151910 325096 163200
rect 325332 157004 325384 157010
rect 325332 156946 325384 156952
rect 325056 151904 325108 151910
rect 325056 151846 325108 151852
rect 325344 150226 325372 156946
rect 325896 152998 325924 163200
rect 326724 154222 326752 163200
rect 327448 160064 327500 160070
rect 327448 160006 327500 160012
rect 327460 159322 327488 160006
rect 327552 159322 327580 163200
rect 328380 159934 328408 163200
rect 329208 160002 329236 163200
rect 329104 159996 329156 160002
rect 329104 159938 329156 159944
rect 329196 159996 329248 160002
rect 329196 159938 329248 159944
rect 328368 159928 328420 159934
rect 328368 159870 328420 159876
rect 328550 159488 328606 159497
rect 328550 159423 328606 159432
rect 327448 159316 327500 159322
rect 327448 159258 327500 159264
rect 327540 159316 327592 159322
rect 327540 159258 327592 159264
rect 327908 157140 327960 157146
rect 327908 157082 327960 157088
rect 326712 154216 326764 154222
rect 326712 154158 326764 154164
rect 327264 153332 327316 153338
rect 327264 153274 327316 153280
rect 325884 152992 325936 152998
rect 325884 152934 325936 152940
rect 325976 152108 326028 152114
rect 325976 152050 326028 152056
rect 325988 150226 326016 152050
rect 326620 151972 326672 151978
rect 326620 151914 326672 151920
rect 326632 150226 326660 151914
rect 327276 150226 327304 153274
rect 327920 150226 327948 157082
rect 328564 150226 328592 159423
rect 329116 151814 329144 159938
rect 330128 155446 330156 163200
rect 330668 160132 330720 160138
rect 330668 160074 330720 160080
rect 330680 159322 330708 160074
rect 330576 159316 330628 159322
rect 330576 159258 330628 159264
rect 330668 159316 330720 159322
rect 330668 159258 330720 159264
rect 330588 158778 330616 159258
rect 330576 158772 330628 158778
rect 330576 158714 330628 158720
rect 330484 157072 330536 157078
rect 330484 157014 330536 157020
rect 330116 155440 330168 155446
rect 330116 155382 330168 155388
rect 329840 154352 329892 154358
rect 329840 154294 329892 154300
rect 329116 151786 329236 151814
rect 329208 150226 329236 151786
rect 329852 150226 329880 154294
rect 330392 152312 330444 152318
rect 330392 152254 330444 152260
rect 330404 152114 330432 152254
rect 330392 152108 330444 152114
rect 330392 152050 330444 152056
rect 330496 150226 330524 157014
rect 330956 152318 330984 163200
rect 331784 161474 331812 163200
rect 331784 161446 331904 161474
rect 331772 153128 331824 153134
rect 331772 153070 331824 153076
rect 330944 152312 330996 152318
rect 330944 152254 330996 152260
rect 331128 152176 331180 152182
rect 331128 152118 331180 152124
rect 331140 150226 331168 152118
rect 331784 150226 331812 153070
rect 331876 152182 331904 161446
rect 332416 154420 332468 154426
rect 332416 154362 332468 154368
rect 331864 152176 331916 152182
rect 331864 152118 331916 152124
rect 332428 150226 332456 154362
rect 332612 153134 332640 163200
rect 332692 157208 332744 157214
rect 332692 157150 332744 157156
rect 332600 153128 332652 153134
rect 332600 153070 332652 153076
rect 332704 151814 332732 157150
rect 333440 155514 333468 163200
rect 334268 160070 334296 163200
rect 335096 160070 335124 163200
rect 336016 163146 336044 163200
rect 336108 163146 336136 163254
rect 336016 163118 336136 163146
rect 335360 160132 335412 160138
rect 335360 160074 335412 160080
rect 334164 160064 334216 160070
rect 334164 160006 334216 160012
rect 334256 160064 334308 160070
rect 334256 160006 334308 160012
rect 335084 160064 335136 160070
rect 335084 160006 335136 160012
rect 333704 159316 333756 159322
rect 333704 159258 333756 159264
rect 333428 155508 333480 155514
rect 333428 155450 333480 155456
rect 332704 151786 333100 151814
rect 333072 150226 333100 151786
rect 333716 150226 333744 159258
rect 334176 151814 334204 160006
rect 335372 159322 335400 160074
rect 335360 159316 335412 159322
rect 335360 159258 335412 159264
rect 335544 156664 335596 156670
rect 335544 156606 335596 156612
rect 334900 153944 334952 153950
rect 334900 153886 334952 153892
rect 334176 151786 334388 151814
rect 334360 150226 334388 151786
rect 334912 150226 334940 153886
rect 335556 150226 335584 156606
rect 336292 152658 336320 163254
rect 336830 163200 336886 164400
rect 337658 163200 337714 164400
rect 338486 163200 338542 164400
rect 339314 163200 339370 164400
rect 340142 163200 340198 164400
rect 340970 163200 341026 164400
rect 341890 163200 341946 164400
rect 342718 163200 342774 164400
rect 343546 163200 343602 164400
rect 344374 163200 344430 164400
rect 345202 163200 345258 164400
rect 346030 163200 346086 164400
rect 346858 163200 346914 164400
rect 347778 163200 347834 164400
rect 348606 163200 348662 164400
rect 348712 163254 349108 163282
rect 336844 153950 336872 163200
rect 337672 156670 337700 163200
rect 338500 161474 338528 163200
rect 338500 161446 338712 161474
rect 338684 159390 338712 161446
rect 339328 159526 339356 163200
rect 339224 159520 339276 159526
rect 339224 159462 339276 159468
rect 339316 159520 339368 159526
rect 339316 159462 339368 159468
rect 338672 159384 338724 159390
rect 338316 159322 338620 159338
rect 338672 159326 338724 159332
rect 339236 159338 339264 159462
rect 339420 159446 339632 159474
rect 339420 159338 339448 159446
rect 339604 159390 339632 159446
rect 338304 159316 338632 159322
rect 338356 159310 338580 159316
rect 338304 159258 338356 159264
rect 339236 159310 339448 159338
rect 339500 159384 339552 159390
rect 339500 159326 339552 159332
rect 339592 159384 339644 159390
rect 339592 159326 339644 159332
rect 338580 159258 338632 159264
rect 338396 159248 338448 159254
rect 338396 159190 338448 159196
rect 338120 156800 338172 156806
rect 338120 156742 338172 156748
rect 337660 156664 337712 156670
rect 337660 156606 337712 156612
rect 336832 153944 336884 153950
rect 336832 153886 336884 153892
rect 337476 153876 337528 153882
rect 337476 153818 337528 153824
rect 336188 152652 336240 152658
rect 336188 152594 336240 152600
rect 336280 152652 336332 152658
rect 336280 152594 336332 152600
rect 336200 150226 336228 152594
rect 336832 152516 336884 152522
rect 336832 152458 336884 152464
rect 336844 150226 336872 152458
rect 337488 150226 337516 153818
rect 338132 150226 338160 156742
rect 338408 151814 338436 159190
rect 339408 159180 339460 159186
rect 339408 159122 339460 159128
rect 338408 151786 338804 151814
rect 338776 150226 338804 151786
rect 339420 150226 339448 159122
rect 339512 152522 339540 159326
rect 339960 157276 340012 157282
rect 339960 157218 340012 157224
rect 339592 155712 339644 155718
rect 339592 155654 339644 155660
rect 339500 152516 339552 152522
rect 339500 152458 339552 152464
rect 339604 151814 339632 155654
rect 339972 151814 340000 157218
rect 340156 153950 340184 163200
rect 340984 155582 341012 163200
rect 341904 159186 341932 163200
rect 342444 159384 342496 159390
rect 342444 159326 342496 159332
rect 342352 159248 342404 159254
rect 342352 159190 342404 159196
rect 341892 159180 341944 159186
rect 341892 159122 341944 159128
rect 340972 155576 341024 155582
rect 340972 155518 341024 155524
rect 340144 153944 340196 153950
rect 340144 153886 340196 153892
rect 342364 153202 342392 159190
rect 342260 153196 342312 153202
rect 342260 153138 342312 153144
rect 342352 153196 342404 153202
rect 342352 153138 342404 153144
rect 341340 152720 341392 152726
rect 341340 152662 341392 152668
rect 339604 151786 339908 151814
rect 339972 151786 340736 151814
rect 339880 150498 339908 151786
rect 339880 150470 340092 150498
rect 340064 150226 340092 150470
rect 340708 150226 340736 151786
rect 321480 150198 321554 150226
rect 322124 150198 322198 150226
rect 322768 150198 322842 150226
rect 323412 150198 323486 150226
rect 324056 150198 324130 150226
rect 324700 150198 324774 150226
rect 325344 150198 325418 150226
rect 325988 150198 326062 150226
rect 326632 150198 326706 150226
rect 327276 150198 327350 150226
rect 327920 150198 327994 150226
rect 328564 150198 328638 150226
rect 329208 150198 329282 150226
rect 329852 150198 329926 150226
rect 330496 150198 330570 150226
rect 331140 150198 331214 150226
rect 331784 150198 331858 150226
rect 332428 150198 332502 150226
rect 333072 150198 333146 150226
rect 333716 150198 333790 150226
rect 334360 150198 334434 150226
rect 334912 150198 334986 150226
rect 335556 150198 335630 150226
rect 336200 150198 336274 150226
rect 336844 150198 336918 150226
rect 337488 150198 337562 150226
rect 338132 150198 338206 150226
rect 338776 150198 338850 150226
rect 339420 150198 339494 150226
rect 340064 150198 340138 150226
rect 340708 150198 340782 150226
rect 320882 149940 320910 150198
rect 321526 149940 321554 150198
rect 322170 149940 322198 150198
rect 322814 149940 322842 150198
rect 323458 149940 323486 150198
rect 324102 149940 324130 150198
rect 324746 149940 324774 150198
rect 325390 149940 325418 150198
rect 326034 149940 326062 150198
rect 326678 149940 326706 150198
rect 327322 149940 327350 150198
rect 327966 149940 327994 150198
rect 328610 149940 328638 150198
rect 329254 149940 329282 150198
rect 329898 149940 329926 150198
rect 330542 149940 330570 150198
rect 331186 149940 331214 150198
rect 331830 149940 331858 150198
rect 332474 149940 332502 150198
rect 333118 149940 333146 150198
rect 333762 149940 333790 150198
rect 334406 149940 334434 150198
rect 334958 149940 334986 150198
rect 335602 149940 335630 150198
rect 336246 149940 336274 150198
rect 336890 149940 336918 150198
rect 337534 149940 337562 150198
rect 338178 149940 338206 150198
rect 338822 149940 338850 150198
rect 339466 149940 339494 150198
rect 340110 149940 340138 150198
rect 340754 149940 340782 150198
rect 341352 150090 341380 152662
rect 342272 152250 342300 153138
rect 342456 152726 342484 159326
rect 342732 159254 342760 163200
rect 342720 159248 342772 159254
rect 342720 159190 342772 159196
rect 343272 156732 343324 156738
rect 343272 156674 343324 156680
rect 342628 155848 342680 155854
rect 342628 155790 342680 155796
rect 342444 152720 342496 152726
rect 342444 152662 342496 152668
rect 341984 152244 342036 152250
rect 341984 152186 342036 152192
rect 342260 152244 342312 152250
rect 342260 152186 342312 152192
rect 341996 150090 342024 152186
rect 342640 150090 342668 155790
rect 343284 150090 343312 156674
rect 343560 154290 343588 163200
rect 343824 159248 343876 159254
rect 343824 159190 343876 159196
rect 343548 154284 343600 154290
rect 343548 154226 343600 154232
rect 343836 151910 343864 159190
rect 344388 156738 344416 163200
rect 345216 161474 345244 163200
rect 345216 161446 345336 161474
rect 344376 156732 344428 156738
rect 344376 156674 344428 156680
rect 345204 155780 345256 155786
rect 345204 155722 345256 155728
rect 343916 153196 343968 153202
rect 343916 153138 343968 153144
rect 343824 151904 343876 151910
rect 343824 151846 343876 151852
rect 343928 150090 343956 153138
rect 344560 152720 344612 152726
rect 344560 152662 344612 152668
rect 344572 150090 344600 152662
rect 345216 150090 345244 155722
rect 345308 153202 345336 161446
rect 346044 159390 346072 163200
rect 346032 159384 346084 159390
rect 346032 159326 346084 159332
rect 345848 156868 345900 156874
rect 345848 156810 345900 156816
rect 345296 153196 345348 153202
rect 345296 153138 345348 153144
rect 345756 153196 345808 153202
rect 345756 153138 345808 153144
rect 345400 152658 345612 152674
rect 345388 152652 345624 152658
rect 345440 152646 345572 152652
rect 345388 152594 345440 152600
rect 345572 152594 345624 152600
rect 345664 152584 345716 152590
rect 345664 152526 345716 152532
rect 345676 152454 345704 152526
rect 345768 152454 345796 153138
rect 345664 152448 345716 152454
rect 345664 152390 345716 152396
rect 345756 152448 345808 152454
rect 345756 152390 345808 152396
rect 345860 150090 345888 156810
rect 346872 154358 346900 163200
rect 347792 159730 347820 163200
rect 348620 163146 348648 163200
rect 348712 163146 348740 163254
rect 348620 163118 348740 163146
rect 347688 159724 347740 159730
rect 347688 159666 347740 159672
rect 347780 159724 347832 159730
rect 347780 159666 347832 159672
rect 347700 159610 347728 159666
rect 347700 159582 348096 159610
rect 348068 159458 348096 159582
rect 347964 159452 348016 159458
rect 347964 159394 348016 159400
rect 348056 159452 348108 159458
rect 348056 159394 348108 159400
rect 347780 155236 347832 155242
rect 347780 155178 347832 155184
rect 346860 154352 346912 154358
rect 346860 154294 346912 154300
rect 347136 152720 347188 152726
rect 347136 152662 347188 152668
rect 346676 152448 346728 152454
rect 346676 152390 346728 152396
rect 346492 152244 346544 152250
rect 346492 152186 346544 152192
rect 346584 152244 346636 152250
rect 346584 152186 346636 152192
rect 346504 150090 346532 152186
rect 346596 151910 346624 152186
rect 346688 151910 346716 152390
rect 346584 151904 346636 151910
rect 346584 151846 346636 151852
rect 346676 151904 346728 151910
rect 346676 151846 346728 151852
rect 347148 150090 347176 152662
rect 347792 150090 347820 155178
rect 347976 150210 348004 159394
rect 348424 158092 348476 158098
rect 348424 158034 348476 158040
rect 348436 150226 348464 158034
rect 349080 152726 349108 163254
rect 349434 163200 349490 164400
rect 350262 163200 350318 164400
rect 351090 163200 351146 164400
rect 351918 163200 351974 164400
rect 352746 163200 352802 164400
rect 353666 163200 353722 164400
rect 354494 163200 354550 164400
rect 355322 163200 355378 164400
rect 356150 163200 356206 164400
rect 356978 163200 357034 164400
rect 357084 163254 357388 163282
rect 349448 153202 349476 163200
rect 349804 159520 349856 159526
rect 349804 159462 349856 159468
rect 349816 159254 349844 159462
rect 349804 159248 349856 159254
rect 349804 159190 349856 159196
rect 349712 159112 349764 159118
rect 349712 159054 349764 159060
rect 349436 153196 349488 153202
rect 349436 153138 349488 153144
rect 349068 152720 349120 152726
rect 349068 152662 349120 152668
rect 349724 150226 349752 159054
rect 350276 154426 350304 163200
rect 351104 159458 351132 163200
rect 351092 159452 351144 159458
rect 351092 159394 351144 159400
rect 351932 159118 351960 163200
rect 351920 159112 351972 159118
rect 351920 159054 351972 159060
rect 350356 155916 350408 155922
rect 350356 155858 350408 155864
rect 350264 154420 350316 154426
rect 350264 154362 350316 154368
rect 347964 150204 348016 150210
rect 348436 150198 348510 150226
rect 347964 150146 348016 150152
rect 341352 150062 341426 150090
rect 341996 150062 342070 150090
rect 342640 150062 342714 150090
rect 343284 150062 343358 150090
rect 343928 150062 344002 150090
rect 344572 150062 344646 150090
rect 345216 150062 345290 150090
rect 345860 150062 345934 150090
rect 346504 150062 346578 150090
rect 347148 150062 347222 150090
rect 347792 150062 347866 150090
rect 341398 149940 341426 150062
rect 342042 149940 342070 150062
rect 342686 149940 342714 150062
rect 343330 149940 343358 150062
rect 343974 149940 344002 150062
rect 344618 149940 344646 150062
rect 345262 149940 345290 150062
rect 345906 149940 345934 150062
rect 346550 149940 346578 150062
rect 347194 149940 347222 150062
rect 347838 149940 347866 150062
rect 348482 149940 348510 150198
rect 349114 150204 349166 150210
rect 349724 150198 349798 150226
rect 349114 150146 349166 150152
rect 349126 149940 349154 150146
rect 349770 149940 349798 150198
rect 350368 150090 350396 155858
rect 352380 152720 352432 152726
rect 352380 152662 352432 152668
rect 352472 152720 352524 152726
rect 352472 152662 352524 152668
rect 352392 152590 352420 152662
rect 352288 152584 352340 152590
rect 352288 152526 352340 152532
rect 352380 152584 352432 152590
rect 352380 152526 352432 152532
rect 351644 152040 351696 152046
rect 351644 151982 351696 151988
rect 351000 151836 351052 151842
rect 351000 151778 351052 151784
rect 351012 150226 351040 151778
rect 351656 150226 351684 151982
rect 352300 150226 352328 152526
rect 352484 151910 352512 152662
rect 352760 152046 352788 163200
rect 353208 159044 353260 159050
rect 353208 158986 353260 158992
rect 352932 155168 352984 155174
rect 352932 155110 352984 155116
rect 352748 152040 352800 152046
rect 352748 151982 352800 151988
rect 352472 151904 352524 151910
rect 352472 151846 352524 151852
rect 352944 150226 352972 155110
rect 353220 151814 353248 158986
rect 353680 154494 353708 163200
rect 354220 159520 354272 159526
rect 354220 159462 354272 159468
rect 353668 154488 353720 154494
rect 353668 154430 353720 154436
rect 353220 151786 353616 151814
rect 353588 150226 353616 151786
rect 354232 150226 354260 159462
rect 354508 152386 354536 163200
rect 354864 159656 354916 159662
rect 354864 159598 354916 159604
rect 355232 159656 355284 159662
rect 355232 159598 355284 159604
rect 354680 155304 354732 155310
rect 354680 155246 354732 155252
rect 354496 152380 354548 152386
rect 354496 152322 354548 152328
rect 351012 150198 351086 150226
rect 351656 150198 351730 150226
rect 352300 150198 352374 150226
rect 352944 150198 353018 150226
rect 353588 150198 353662 150226
rect 354232 150198 354306 150226
rect 354692 150210 354720 155246
rect 354876 150226 354904 159598
rect 355244 158846 355272 159598
rect 355232 158840 355284 158846
rect 355232 158782 355284 158788
rect 355336 151910 355364 163200
rect 356164 159458 356192 163200
rect 356992 163146 357020 163200
rect 357084 163146 357112 163254
rect 356992 163118 357112 163146
rect 355600 159452 355652 159458
rect 355600 159394 355652 159400
rect 356152 159452 356204 159458
rect 356152 159394 356204 159400
rect 355612 159050 355640 159394
rect 355600 159044 355652 159050
rect 355600 158986 355652 158992
rect 357360 154562 357388 163254
rect 357806 163200 357862 164400
rect 358634 163200 358690 164400
rect 359554 163200 359610 164400
rect 360382 163200 360438 164400
rect 361210 163200 361266 164400
rect 362038 163200 362094 164400
rect 362866 163200 362922 164400
rect 363694 163200 363750 164400
rect 364522 163200 364578 164400
rect 365442 163200 365498 164400
rect 366270 163200 366326 164400
rect 367098 163200 367154 164400
rect 367926 163200 367982 164400
rect 368754 163200 368810 164400
rect 369582 163200 369638 164400
rect 370410 163200 370466 164400
rect 371330 163200 371386 164400
rect 372158 163200 372214 164400
rect 372986 163200 373042 164400
rect 373814 163200 373870 164400
rect 374642 163200 374698 164400
rect 375470 163200 375526 164400
rect 376298 163200 376354 164400
rect 377218 163200 377274 164400
rect 378046 163200 378102 164400
rect 378874 163200 378930 164400
rect 379702 163200 379758 164400
rect 380530 163200 380586 164400
rect 380636 163254 380848 163282
rect 357532 159860 357584 159866
rect 357532 159802 357584 159808
rect 357544 158982 357572 159802
rect 357820 159798 357848 163200
rect 357992 159860 358044 159866
rect 357992 159802 358044 159808
rect 357808 159792 357860 159798
rect 357808 159734 357860 159740
rect 357440 158976 357492 158982
rect 357440 158918 357492 158924
rect 357532 158976 357584 158982
rect 357532 158918 357584 158924
rect 357348 154556 357400 154562
rect 357348 154498 357400 154504
rect 357452 152794 357480 158918
rect 357900 154012 357952 154018
rect 357900 153954 357952 153960
rect 356796 152788 356848 152794
rect 356796 152730 356848 152736
rect 357440 152788 357492 152794
rect 357440 152730 357492 152736
rect 356152 152448 356204 152454
rect 356152 152390 356204 152396
rect 355324 151904 355376 151910
rect 355324 151846 355376 151852
rect 356164 150226 356192 152390
rect 356808 150226 356836 152730
rect 357438 152416 357494 152425
rect 357438 152351 357494 152360
rect 357452 150226 357480 152351
rect 357912 150498 357940 153954
rect 358004 151814 358032 159802
rect 358648 159526 358676 163200
rect 358912 159588 358964 159594
rect 358912 159530 358964 159536
rect 358636 159520 358688 159526
rect 358636 159462 358688 159468
rect 358004 151786 358768 151814
rect 357912 150470 358124 150498
rect 358096 150226 358124 150470
rect 358740 150226 358768 151786
rect 350368 150062 350442 150090
rect 350414 149940 350442 150062
rect 351058 149940 351086 150198
rect 351702 149940 351730 150198
rect 352346 149940 352374 150198
rect 352990 149940 353018 150198
rect 353634 149940 353662 150198
rect 354278 149940 354306 150198
rect 354680 150204 354732 150210
rect 354876 150198 354950 150226
rect 354680 150146 354732 150152
rect 354922 149940 354950 150198
rect 355554 150204 355606 150210
rect 356164 150198 356238 150226
rect 356808 150198 356882 150226
rect 357452 150198 357526 150226
rect 358096 150198 358170 150226
rect 358740 150198 358814 150226
rect 358924 150210 358952 159530
rect 359568 152794 359596 163200
rect 360396 153814 360424 163200
rect 361224 161474 361252 163200
rect 361224 161446 361344 161474
rect 361316 158846 361344 161446
rect 361304 158840 361356 158846
rect 361304 158782 361356 158788
rect 360660 155372 360712 155378
rect 360660 155314 360712 155320
rect 360384 153808 360436 153814
rect 360384 153750 360436 153756
rect 359372 152788 359424 152794
rect 359372 152730 359424 152736
rect 359556 152788 359608 152794
rect 359556 152730 359608 152736
rect 359384 150226 359412 152730
rect 360672 150226 360700 155314
rect 361304 153060 361356 153066
rect 361304 153002 361356 153008
rect 361316 150226 361344 153002
rect 362052 152862 362080 163200
rect 362880 159594 362908 163200
rect 362960 159656 363012 159662
rect 362960 159598 363012 159604
rect 362868 159588 362920 159594
rect 362868 159530 362920 159536
rect 361948 152856 362000 152862
rect 361948 152798 362000 152804
rect 362040 152856 362092 152862
rect 362040 152798 362092 152804
rect 361960 150226 361988 152798
rect 362592 152108 362644 152114
rect 362592 152050 362644 152056
rect 362604 150226 362632 152050
rect 362972 151978 363000 159598
rect 363512 158976 363564 158982
rect 363512 158918 363564 158924
rect 363236 154080 363288 154086
rect 363236 154022 363288 154028
rect 362960 151972 363012 151978
rect 362960 151914 363012 151920
rect 363248 150226 363276 154022
rect 363524 151814 363552 158918
rect 363708 154018 363736 163200
rect 363696 154012 363748 154018
rect 363696 153954 363748 153960
rect 364536 152386 364564 163200
rect 365456 159798 365484 163200
rect 366284 161474 366312 163200
rect 366284 161446 366496 161474
rect 365352 159792 365404 159798
rect 365352 159734 365404 159740
rect 365444 159792 365496 159798
rect 365444 159734 365496 159740
rect 365364 158982 365392 159734
rect 365168 158976 365220 158982
rect 365168 158918 365220 158924
rect 365352 158976 365404 158982
rect 365352 158918 365404 158924
rect 364524 152380 364576 152386
rect 364524 152322 364576 152328
rect 364524 151972 364576 151978
rect 364524 151914 364576 151920
rect 363524 151786 363920 151814
rect 363892 150226 363920 151786
rect 364536 150226 364564 151914
rect 365180 150226 365208 158918
rect 365720 154148 365772 154154
rect 365720 154090 365772 154096
rect 365732 150226 365760 154090
rect 366468 152930 366496 161446
rect 367112 155242 367140 163200
rect 367940 158778 367968 163200
rect 367192 158772 367244 158778
rect 367192 158714 367244 158720
rect 367928 158772 367980 158778
rect 367928 158714 367980 158720
rect 367100 155236 367152 155242
rect 367100 155178 367152 155184
rect 367204 153066 367232 158714
rect 368296 154216 368348 154222
rect 368296 154158 368348 154164
rect 367192 153060 367244 153066
rect 367192 153002 367244 153008
rect 367652 152992 367704 152998
rect 367652 152934 367704 152940
rect 366364 152924 366416 152930
rect 366364 152866 366416 152872
rect 366456 152924 366508 152930
rect 366456 152866 366508 152872
rect 366376 150226 366404 152866
rect 367008 151836 367060 151842
rect 367008 151778 367060 151784
rect 367020 150226 367048 151778
rect 367664 150226 367692 152934
rect 368308 150226 368336 154158
rect 368768 152998 368796 163200
rect 369492 159928 369544 159934
rect 369492 159870 369544 159876
rect 368940 153060 368992 153066
rect 368940 153002 368992 153008
rect 369032 153060 369084 153066
rect 369032 153002 369084 153008
rect 368756 152992 368808 152998
rect 368756 152934 368808 152940
rect 368952 150226 368980 153002
rect 369044 152386 369072 153002
rect 369032 152380 369084 152386
rect 369032 152322 369084 152328
rect 369504 151814 369532 159870
rect 369596 159662 369624 163200
rect 370228 159996 370280 160002
rect 370228 159938 370280 159944
rect 369584 159656 369636 159662
rect 369584 159598 369636 159604
rect 369860 155440 369912 155446
rect 369860 155382 369912 155388
rect 369504 151786 369624 151814
rect 369596 150226 369624 151786
rect 355554 150146 355606 150152
rect 355566 149940 355594 150146
rect 356210 149940 356238 150198
rect 356854 149940 356882 150198
rect 357498 149940 357526 150198
rect 358142 149940 358170 150198
rect 358786 149940 358814 150198
rect 358912 150204 358964 150210
rect 359384 150198 359458 150226
rect 358912 150146 358964 150152
rect 359430 149940 359458 150198
rect 360062 150204 360114 150210
rect 360672 150198 360746 150226
rect 361316 150198 361390 150226
rect 361960 150198 362034 150226
rect 362604 150198 362678 150226
rect 363248 150198 363322 150226
rect 363892 150198 363966 150226
rect 364536 150198 364610 150226
rect 365180 150198 365254 150226
rect 365732 150198 365806 150226
rect 366376 150198 366450 150226
rect 367020 150198 367094 150226
rect 367664 150198 367738 150226
rect 368308 150198 368382 150226
rect 368952 150198 369026 150226
rect 369596 150198 369670 150226
rect 369872 150210 369900 155382
rect 370240 150226 370268 159938
rect 370424 154086 370452 163200
rect 370412 154080 370464 154086
rect 370412 154022 370464 154028
rect 371344 152386 371372 163200
rect 372172 159934 372200 163200
rect 372160 159928 372212 159934
rect 372160 159870 372212 159876
rect 373000 153134 373028 163200
rect 373448 155508 373500 155514
rect 373448 155450 373500 155456
rect 372804 153128 372856 153134
rect 372804 153070 372856 153076
rect 372988 153128 373040 153134
rect 372988 153070 373040 153076
rect 371332 152380 371384 152386
rect 371332 152322 371384 152328
rect 371516 152312 371568 152318
rect 371516 152254 371568 152260
rect 371528 150226 371556 152254
rect 372160 152176 372212 152182
rect 372160 152118 372212 152124
rect 372172 150226 372200 152118
rect 372816 150226 372844 153070
rect 373460 150226 373488 155450
rect 373828 155310 373856 163200
rect 374656 160002 374684 163200
rect 374736 160064 374788 160070
rect 374736 160006 374788 160012
rect 374644 159996 374696 160002
rect 374644 159938 374696 159944
rect 374092 159316 374144 159322
rect 374092 159258 374144 159264
rect 373816 155304 373868 155310
rect 373816 155246 373868 155252
rect 374104 150226 374132 159258
rect 374748 150226 374776 160006
rect 375484 152658 375512 163200
rect 376312 159866 376340 163200
rect 376300 159860 376352 159866
rect 376300 159802 376352 159808
rect 375564 156664 375616 156670
rect 375564 156606 375616 156612
rect 375380 152652 375432 152658
rect 375380 152594 375432 152600
rect 375472 152652 375524 152658
rect 375472 152594 375524 152600
rect 375392 150226 375420 152594
rect 360062 150146 360114 150152
rect 360074 149940 360102 150146
rect 360718 149940 360746 150198
rect 361362 149940 361390 150198
rect 362006 149940 362034 150198
rect 362650 149940 362678 150198
rect 363294 149940 363322 150198
rect 363938 149940 363966 150198
rect 364582 149940 364610 150198
rect 365226 149940 365254 150198
rect 365778 149940 365806 150198
rect 366422 149940 366450 150198
rect 367066 149940 367094 150198
rect 367710 149940 367738 150198
rect 368354 149940 368382 150198
rect 368998 149940 369026 150198
rect 369642 149940 369670 150198
rect 369860 150204 369912 150210
rect 370240 150198 370314 150226
rect 369860 150146 369912 150152
rect 370286 149940 370314 150198
rect 370918 150204 370970 150210
rect 371528 150198 371602 150226
rect 372172 150198 372246 150226
rect 372816 150198 372890 150226
rect 373460 150198 373534 150226
rect 374104 150198 374178 150226
rect 374748 150198 374822 150226
rect 375392 150198 375466 150226
rect 375576 150210 375604 156606
rect 377232 153882 377260 163200
rect 378060 159322 378088 163200
rect 378888 160070 378916 163200
rect 378876 160064 378928 160070
rect 378876 160006 378928 160012
rect 379716 159730 379744 163200
rect 380544 163146 380572 163200
rect 380636 163146 380664 163254
rect 380544 163118 380664 163146
rect 378784 159724 378836 159730
rect 378784 159666 378836 159672
rect 379704 159724 379756 159730
rect 379704 159666 379756 159672
rect 378048 159316 378100 159322
rect 378048 159258 378100 159264
rect 377956 159248 378008 159254
rect 377956 159190 378008 159196
rect 376024 153876 376076 153882
rect 376024 153818 376076 153824
rect 377220 153876 377272 153882
rect 377220 153818 377272 153824
rect 376036 150226 376064 153818
rect 377312 152516 377364 152522
rect 377312 152458 377364 152464
rect 377324 150226 377352 152458
rect 377968 150226 377996 159190
rect 378232 159180 378284 159186
rect 378232 159122 378284 159128
rect 378140 155576 378192 155582
rect 378140 155518 378192 155524
rect 370918 150146 370970 150152
rect 370930 149940 370958 150146
rect 371574 149940 371602 150198
rect 372218 149940 372246 150198
rect 372862 149940 372890 150198
rect 373506 149940 373534 150198
rect 374150 149940 374178 150198
rect 374794 149940 374822 150198
rect 375438 149940 375466 150198
rect 375564 150204 375616 150210
rect 376036 150198 376110 150226
rect 375564 150146 375616 150152
rect 376082 149940 376110 150198
rect 376714 150204 376766 150210
rect 377324 150198 377398 150226
rect 377968 150198 378042 150226
rect 378152 150210 378180 155518
rect 378244 152522 378272 159122
rect 378692 158976 378744 158982
rect 378692 158918 378744 158924
rect 378704 158778 378732 158918
rect 378692 158772 378744 158778
rect 378692 158714 378744 158720
rect 378600 153944 378652 153950
rect 378600 153886 378652 153892
rect 378232 152516 378284 152522
rect 378232 152458 378284 152464
rect 378612 150226 378640 153886
rect 378796 151842 378824 159666
rect 380820 153950 380848 163254
rect 381358 163200 381414 164400
rect 382186 163200 382242 164400
rect 383106 163200 383162 164400
rect 383934 163200 383990 164400
rect 384762 163200 384818 164400
rect 385590 163200 385646 164400
rect 386418 163200 386474 164400
rect 387246 163200 387302 164400
rect 387352 163254 387656 163282
rect 381176 154284 381228 154290
rect 381176 154226 381228 154232
rect 380808 153944 380860 153950
rect 380808 153886 380860 153892
rect 379888 152516 379940 152522
rect 379888 152458 379940 152464
rect 378784 151836 378836 151842
rect 378784 151778 378836 151784
rect 379900 150226 379928 152458
rect 380532 152244 380584 152250
rect 380532 152186 380584 152192
rect 380544 150226 380572 152186
rect 381188 150226 381216 154226
rect 381372 152318 381400 163200
rect 381820 156732 381872 156738
rect 381820 156674 381872 156680
rect 381360 152312 381412 152318
rect 381360 152254 381412 152260
rect 381832 150226 381860 156674
rect 382200 152522 382228 163200
rect 382832 159384 382884 159390
rect 382832 159326 382884 159332
rect 382556 159044 382608 159050
rect 382556 158986 382608 158992
rect 382568 152726 382596 158986
rect 382464 152720 382516 152726
rect 382464 152662 382516 152668
rect 382556 152720 382608 152726
rect 382556 152662 382608 152668
rect 382188 152516 382240 152522
rect 382188 152458 382240 152464
rect 382476 150226 382504 152662
rect 382844 151814 382872 159326
rect 383120 159050 383148 163200
rect 383108 159044 383160 159050
rect 383108 158986 383160 158992
rect 383752 154352 383804 154358
rect 383752 154294 383804 154300
rect 382844 151786 383148 151814
rect 383120 150226 383148 151786
rect 383764 150226 383792 154294
rect 383948 154154 383976 163200
rect 384776 158914 384804 163200
rect 385604 159254 385632 163200
rect 385592 159248 385644 159254
rect 385592 159190 385644 159196
rect 386432 159118 386460 163200
rect 387260 163146 387288 163200
rect 387352 163146 387380 163254
rect 387260 163118 387380 163146
rect 385500 159112 385552 159118
rect 385500 159054 385552 159060
rect 386420 159112 386472 159118
rect 386420 159054 386472 159060
rect 384764 158908 384816 158914
rect 384764 158850 384816 158856
rect 384948 158840 385000 158846
rect 384948 158782 385000 158788
rect 383936 154148 383988 154154
rect 383936 154090 383988 154096
rect 384960 152250 384988 158782
rect 385316 158772 385368 158778
rect 385316 158714 385368 158720
rect 385040 152584 385092 152590
rect 385040 152526 385092 152532
rect 384948 152244 385000 152250
rect 384948 152186 385000 152192
rect 384396 151836 384448 151842
rect 384396 151778 384448 151784
rect 384408 150226 384436 151778
rect 385052 150226 385080 152526
rect 385328 151842 385356 158714
rect 385512 152590 385540 159054
rect 386236 158976 386288 158982
rect 386236 158918 386288 158924
rect 385592 153196 385644 153202
rect 385592 153138 385644 153144
rect 385500 152584 385552 152590
rect 385500 152526 385552 152532
rect 385316 151836 385368 151842
rect 385604 151814 385632 153138
rect 386248 151978 386276 158918
rect 386328 154420 386380 154426
rect 386328 154362 386380 154368
rect 386236 151972 386288 151978
rect 386236 151914 386288 151920
rect 385604 151786 385724 151814
rect 385316 151778 385368 151784
rect 385696 150226 385724 151786
rect 386340 150226 386368 154362
rect 387628 154222 387656 163254
rect 388074 163200 388130 164400
rect 388994 163200 389050 164400
rect 389822 163200 389878 164400
rect 390650 163200 390706 164400
rect 391478 163200 391534 164400
rect 392306 163200 392362 164400
rect 393134 163200 393190 164400
rect 393962 163200 394018 164400
rect 394882 163200 394938 164400
rect 395710 163200 395766 164400
rect 396538 163200 396594 164400
rect 397366 163200 397422 164400
rect 398194 163200 398250 164400
rect 399022 163200 399078 164400
rect 399850 163200 399906 164400
rect 399956 163254 400168 163282
rect 387708 159112 387760 159118
rect 387708 159054 387760 159060
rect 387616 154216 387668 154222
rect 387616 154158 387668 154164
rect 387720 152726 387748 159054
rect 388088 158778 388116 163200
rect 388444 159996 388496 160002
rect 388444 159938 388496 159944
rect 388352 159316 388404 159322
rect 388352 159258 388404 159264
rect 388076 158772 388128 158778
rect 388076 158714 388128 158720
rect 386972 152720 387024 152726
rect 386972 152662 387024 152668
rect 387708 152720 387760 152726
rect 387708 152662 387760 152668
rect 386984 150226 387012 152662
rect 387616 152584 387668 152590
rect 387616 152526 387668 152532
rect 387628 150226 387656 152526
rect 388364 152182 388392 159258
rect 388352 152176 388404 152182
rect 388352 152118 388404 152124
rect 388456 152114 388484 159938
rect 389008 159322 389036 163200
rect 389836 160002 389864 163200
rect 389824 159996 389876 160002
rect 389824 159938 389876 159944
rect 388996 159316 389048 159322
rect 388996 159258 389048 159264
rect 389640 158908 389692 158914
rect 389640 158850 389692 158856
rect 388904 154488 388956 154494
rect 388904 154430 388956 154436
rect 388444 152108 388496 152114
rect 388444 152050 388496 152056
rect 388260 152040 388312 152046
rect 388260 151982 388312 151988
rect 388272 150226 388300 151982
rect 388916 150226 388944 154430
rect 389652 152454 389680 158850
rect 390376 158772 390428 158778
rect 390376 158714 390428 158720
rect 390388 153202 390416 158714
rect 390664 154358 390692 163200
rect 390836 159452 390888 159458
rect 390836 159394 390888 159400
rect 390652 154352 390704 154358
rect 390652 154294 390704 154300
rect 390376 153196 390428 153202
rect 390376 153138 390428 153144
rect 389548 152448 389600 152454
rect 389548 152390 389600 152396
rect 389640 152448 389692 152454
rect 389640 152390 389692 152396
rect 389560 150226 389588 152390
rect 390192 151904 390244 151910
rect 390192 151846 390244 151852
rect 390204 150226 390232 151846
rect 390848 150226 390876 159394
rect 391492 158982 391520 163200
rect 392320 159390 392348 163200
rect 392768 159520 392820 159526
rect 392768 159462 392820 159468
rect 392308 159384 392360 159390
rect 392308 159326 392360 159332
rect 391480 158976 391532 158982
rect 391480 158918 391532 158924
rect 391480 154556 391532 154562
rect 391480 154498 391532 154504
rect 391492 150226 391520 154498
rect 392124 152244 392176 152250
rect 392124 152186 392176 152192
rect 392136 150226 392164 152186
rect 392780 150226 392808 159462
rect 393148 152590 393176 163200
rect 393976 154290 394004 163200
rect 394792 159588 394844 159594
rect 394792 159530 394844 159536
rect 394332 158976 394384 158982
rect 394332 158918 394384 158924
rect 393964 154284 394016 154290
rect 393964 154226 394016 154232
rect 394056 153808 394108 153814
rect 394056 153750 394108 153756
rect 393412 152788 393464 152794
rect 393412 152730 393464 152736
rect 393136 152584 393188 152590
rect 393136 152526 393188 152532
rect 393424 150226 393452 152730
rect 394068 150226 394096 153750
rect 394344 152250 394372 158918
rect 394332 152244 394384 152250
rect 394332 152186 394384 152192
rect 394700 151836 394752 151842
rect 394804 151814 394832 159530
rect 394896 152794 394924 163200
rect 395528 159792 395580 159798
rect 395528 159734 395580 159740
rect 395540 152862 395568 159734
rect 395724 159186 395752 163200
rect 396172 159928 396224 159934
rect 396172 159870 396224 159876
rect 395712 159180 395764 159186
rect 395712 159122 395764 159128
rect 395436 152856 395488 152862
rect 395436 152798 395488 152804
rect 395528 152856 395580 152862
rect 395528 152798 395580 152804
rect 394884 152788 394936 152794
rect 394884 152730 394936 152736
rect 394804 151786 394924 151814
rect 394700 151778 394752 151784
rect 394712 150226 394740 151778
rect 376714 150146 376766 150152
rect 376726 149940 376754 150146
rect 377370 149940 377398 150198
rect 378014 149940 378042 150198
rect 378140 150204 378192 150210
rect 378612 150198 378686 150226
rect 378140 150146 378192 150152
rect 378658 149940 378686 150198
rect 379290 150204 379342 150210
rect 379900 150198 379974 150226
rect 380544 150198 380618 150226
rect 381188 150198 381262 150226
rect 381832 150198 381906 150226
rect 382476 150198 382550 150226
rect 383120 150198 383194 150226
rect 383764 150198 383838 150226
rect 384408 150198 384482 150226
rect 385052 150198 385126 150226
rect 385696 150198 385770 150226
rect 386340 150198 386414 150226
rect 386984 150198 387058 150226
rect 387628 150198 387702 150226
rect 388272 150198 388346 150226
rect 388916 150198 388990 150226
rect 389560 150198 389634 150226
rect 390204 150198 390278 150226
rect 390848 150198 390922 150226
rect 391492 150198 391566 150226
rect 392136 150198 392210 150226
rect 392780 150198 392854 150226
rect 393424 150198 393498 150226
rect 394068 150198 394142 150226
rect 394712 150198 394786 150226
rect 394896 150210 394924 151786
rect 395448 150226 395476 152798
rect 396184 151842 396212 159870
rect 396552 159798 396580 163200
rect 396540 159792 396592 159798
rect 396540 159734 396592 159740
rect 397380 154018 397408 163200
rect 398104 160064 398156 160070
rect 398104 160006 398156 160012
rect 396540 154012 396592 154018
rect 396540 153954 396592 153960
rect 397368 154012 397420 154018
rect 397368 153954 397420 153960
rect 396172 151836 396224 151842
rect 396172 151778 396224 151784
rect 379290 150146 379342 150152
rect 379302 149940 379330 150146
rect 379946 149940 379974 150198
rect 380590 149940 380618 150198
rect 381234 149940 381262 150198
rect 381878 149940 381906 150198
rect 382522 149940 382550 150198
rect 383166 149940 383194 150198
rect 383810 149940 383838 150198
rect 384454 149940 384482 150198
rect 385098 149940 385126 150198
rect 385742 149940 385770 150198
rect 386386 149940 386414 150198
rect 387030 149940 387058 150198
rect 387674 149940 387702 150198
rect 388318 149940 388346 150198
rect 388962 149940 388990 150198
rect 389606 149940 389634 150198
rect 390250 149940 390278 150198
rect 390894 149940 390922 150198
rect 391538 149940 391566 150198
rect 392182 149940 392210 150198
rect 392826 149940 392854 150198
rect 393470 149940 393498 150198
rect 394114 149940 394142 150198
rect 394758 149940 394786 150198
rect 394884 150204 394936 150210
rect 394884 150146 394936 150152
rect 395402 150198 395476 150226
rect 396552 150226 396580 153954
rect 398116 153066 398144 160006
rect 398208 154426 398236 163200
rect 399036 159594 399064 163200
rect 399864 163146 399892 163200
rect 399956 163146 399984 163254
rect 399864 163118 399984 163146
rect 399024 159588 399076 159594
rect 399024 159530 399076 159536
rect 399852 159248 399904 159254
rect 399852 159190 399904 159196
rect 399116 155236 399168 155242
rect 399116 155178 399168 155184
rect 398196 154420 398248 154426
rect 398196 154362 398248 154368
rect 397184 153060 397236 153066
rect 397184 153002 397236 153008
rect 398104 153060 398156 153066
rect 398104 153002 398156 153008
rect 397196 150226 397224 153002
rect 398472 152924 398524 152930
rect 398472 152866 398524 152872
rect 397828 152856 397880 152862
rect 397828 152798 397880 152804
rect 397840 150226 397868 152798
rect 398484 150226 398512 152866
rect 399128 150226 399156 155178
rect 399864 151978 399892 159190
rect 400140 152862 400168 163254
rect 400770 163200 400826 164400
rect 401598 163200 401654 164400
rect 402426 163200 402482 164400
rect 403254 163200 403310 164400
rect 404082 163200 404138 164400
rect 404910 163200 404966 164400
rect 405738 163200 405794 164400
rect 406658 163200 406714 164400
rect 406764 163254 407068 163282
rect 400784 154494 400812 163200
rect 401048 159656 401100 159662
rect 401048 159598 401100 159604
rect 400772 154488 400824 154494
rect 400772 154430 400824 154436
rect 400404 152992 400456 152998
rect 400404 152934 400456 152940
rect 400128 152856 400180 152862
rect 400128 152798 400180 152804
rect 399760 151972 399812 151978
rect 399760 151914 399812 151920
rect 399852 151972 399904 151978
rect 399852 151914 399904 151920
rect 399772 150226 399800 151914
rect 400416 150226 400444 152934
rect 401060 150226 401088 159598
rect 401612 155242 401640 163200
rect 401600 155236 401652 155242
rect 401600 155178 401652 155184
rect 401692 154080 401744 154086
rect 401692 154022 401744 154028
rect 401704 150226 401732 154022
rect 402440 152930 402468 163200
rect 403268 159934 403296 163200
rect 404096 160070 404124 163200
rect 404084 160064 404136 160070
rect 404084 160006 404136 160012
rect 403256 159928 403308 159934
rect 403256 159870 403308 159876
rect 403440 159384 403492 159390
rect 403440 159326 403492 159332
rect 403164 155304 403216 155310
rect 403164 155246 403216 155252
rect 402428 152924 402480 152930
rect 402428 152866 402480 152872
rect 402336 152380 402388 152386
rect 402336 152322 402388 152328
rect 402348 150226 402376 152322
rect 402980 151836 403032 151842
rect 402980 151778 403032 151784
rect 402992 150226 403020 151778
rect 396034 150204 396086 150210
rect 395402 149940 395430 150198
rect 396552 150198 396626 150226
rect 397196 150198 397270 150226
rect 397840 150198 397914 150226
rect 398484 150198 398558 150226
rect 399128 150198 399202 150226
rect 399772 150198 399846 150226
rect 400416 150198 400490 150226
rect 401060 150198 401134 150226
rect 401704 150198 401778 150226
rect 402348 150198 402422 150226
rect 402992 150198 403066 150226
rect 403176 150210 403204 155246
rect 403452 152046 403480 159326
rect 403900 159316 403952 159322
rect 403900 159258 403952 159264
rect 403624 153128 403676 153134
rect 403624 153070 403676 153076
rect 403440 152040 403492 152046
rect 403440 151982 403492 151988
rect 403636 150226 403664 153070
rect 403912 151910 403940 159258
rect 404924 158846 404952 163200
rect 405372 159180 405424 159186
rect 405372 159122 405424 159128
rect 404912 158840 404964 158846
rect 404912 158782 404964 158788
rect 405384 152114 405412 159122
rect 405648 158840 405700 158846
rect 405648 158782 405700 158788
rect 405660 152658 405688 158782
rect 405752 158778 405780 163200
rect 406672 163146 406700 163200
rect 406764 163146 406792 163254
rect 406672 163118 406792 163146
rect 406200 159860 406252 159866
rect 406200 159802 406252 159808
rect 405832 159724 405884 159730
rect 405832 159666 405884 159672
rect 405740 158772 405792 158778
rect 405740 158714 405792 158720
rect 405556 152652 405608 152658
rect 405556 152594 405608 152600
rect 405648 152652 405700 152658
rect 405648 152594 405700 152600
rect 404912 152108 404964 152114
rect 404912 152050 404964 152056
rect 405372 152108 405424 152114
rect 405372 152050 405424 152056
rect 403900 151904 403952 151910
rect 403900 151846 403952 151852
rect 404924 150226 404952 152050
rect 405568 150226 405596 152594
rect 405844 152386 405872 159666
rect 405832 152380 405884 152386
rect 405832 152322 405884 152328
rect 406212 150226 406240 159802
rect 406844 153876 406896 153882
rect 406844 153818 406896 153824
rect 406856 150226 406884 153818
rect 407040 152998 407068 163254
rect 407486 163200 407542 164400
rect 408314 163200 408370 164400
rect 409142 163200 409198 164400
rect 409970 163200 410026 164400
rect 410798 163200 410854 164400
rect 411626 163200 411682 164400
rect 412546 163200 412602 164400
rect 413374 163200 413430 164400
rect 414202 163200 414258 164400
rect 415030 163200 415086 164400
rect 415136 163254 415348 163282
rect 407500 159526 407528 163200
rect 407488 159520 407540 159526
rect 407488 159462 407540 159468
rect 408132 153060 408184 153066
rect 408132 153002 408184 153008
rect 407028 152992 407080 152998
rect 407028 152934 407080 152940
rect 407488 152176 407540 152182
rect 407488 152118 407540 152124
rect 407500 150226 407528 152118
rect 408144 150226 408172 153002
rect 408328 152425 408356 163200
rect 408500 159588 408552 159594
rect 408500 159530 408552 159536
rect 408512 153134 408540 159530
rect 409156 158982 409184 163200
rect 409984 159730 410012 163200
rect 409972 159724 410024 159730
rect 409972 159666 410024 159672
rect 410812 159594 410840 163200
rect 410800 159588 410852 159594
rect 410800 159530 410852 159536
rect 411444 159044 411496 159050
rect 411444 158986 411496 158992
rect 409144 158976 409196 158982
rect 409144 158918 409196 158924
rect 410892 158976 410944 158982
rect 410892 158918 410944 158924
rect 409144 158772 409196 158778
rect 409144 158714 409196 158720
rect 408500 153128 408552 153134
rect 408500 153070 408552 153076
rect 408314 152416 408370 152425
rect 409156 152386 409184 158714
rect 409420 153944 409472 153950
rect 409420 153886 409472 153892
rect 408314 152351 408370 152360
rect 408776 152380 408828 152386
rect 408776 152322 408828 152328
rect 409144 152380 409196 152386
rect 409144 152322 409196 152328
rect 408788 150226 408816 152322
rect 409432 150226 409460 153886
rect 410708 152516 410760 152522
rect 410708 152458 410760 152464
rect 410064 152312 410116 152318
rect 410064 152254 410116 152260
rect 410076 150226 410104 152254
rect 410720 150226 410748 152458
rect 410904 152386 410932 158918
rect 410892 152380 410944 152386
rect 410892 152322 410944 152328
rect 411456 150226 411484 158986
rect 411640 153066 411668 163200
rect 412560 159118 412588 163200
rect 412548 159112 412600 159118
rect 412548 159054 412600 159060
rect 413388 158778 413416 163200
rect 413836 159996 413888 160002
rect 413836 159938 413888 159944
rect 413652 159792 413704 159798
rect 413652 159734 413704 159740
rect 413376 158772 413428 158778
rect 413376 158714 413428 158720
rect 411996 154148 412048 154154
rect 411996 154090 412048 154096
rect 411628 153060 411680 153066
rect 411628 153002 411680 153008
rect 396034 150146 396086 150152
rect 396046 149940 396074 150146
rect 396598 149940 396626 150198
rect 397242 149940 397270 150198
rect 397886 149940 397914 150198
rect 398530 149940 398558 150198
rect 399174 149940 399202 150198
rect 399818 149940 399846 150198
rect 400462 149940 400490 150198
rect 401106 149940 401134 150198
rect 401750 149940 401778 150198
rect 402394 149940 402422 150198
rect 403038 149940 403066 150198
rect 403164 150204 403216 150210
rect 403636 150198 403710 150226
rect 403164 150146 403216 150152
rect 403682 149940 403710 150198
rect 404314 150204 404366 150210
rect 404924 150198 404998 150226
rect 405568 150198 405642 150226
rect 406212 150198 406286 150226
rect 406856 150198 406930 150226
rect 407500 150198 407574 150226
rect 408144 150198 408218 150226
rect 408788 150198 408862 150226
rect 409432 150198 409506 150226
rect 410076 150198 410150 150226
rect 410720 150198 410794 150226
rect 404314 150146 404366 150152
rect 404326 149940 404354 150146
rect 404970 149940 404998 150198
rect 405614 149940 405642 150198
rect 406258 149940 406286 150198
rect 406902 149940 406930 150198
rect 407546 149940 407574 150198
rect 408190 149940 408218 150198
rect 408834 149940 408862 150198
rect 409478 149940 409506 150198
rect 410122 149940 410150 150198
rect 410766 149940 410794 150198
rect 411410 150198 411484 150226
rect 412008 150226 412036 154090
rect 412640 152448 412692 152454
rect 412640 152390 412692 152396
rect 412652 150226 412680 152390
rect 413664 151842 413692 159734
rect 413848 151978 413876 159938
rect 414216 159662 414244 163200
rect 415044 163146 415072 163200
rect 415136 163146 415164 163254
rect 415044 163118 415164 163146
rect 414204 159656 414256 159662
rect 414204 159598 414256 159604
rect 413928 159112 413980 159118
rect 413928 159054 413980 159060
rect 413940 152810 413968 159054
rect 414572 154216 414624 154222
rect 414572 154158 414624 154164
rect 413940 152782 414060 152810
rect 414032 152726 414060 152782
rect 413928 152720 413980 152726
rect 413928 152662 413980 152668
rect 414020 152720 414072 152726
rect 414020 152662 414072 152668
rect 413836 151972 413888 151978
rect 413836 151914 413888 151920
rect 413284 151836 413336 151842
rect 413284 151778 413336 151784
rect 413652 151836 413704 151842
rect 413652 151778 413704 151784
rect 413296 150226 413324 151778
rect 413940 150226 413968 152662
rect 414584 150226 414612 154158
rect 415216 153196 415268 153202
rect 415216 153138 415268 153144
rect 415124 153128 415176 153134
rect 415124 153070 415176 153076
rect 415136 152182 415164 153070
rect 415124 152176 415176 152182
rect 415124 152118 415176 152124
rect 415228 150226 415256 153138
rect 415320 153134 415348 163254
rect 415858 163200 415914 164400
rect 416686 163200 416742 164400
rect 417514 163200 417570 164400
rect 418434 163200 418490 164400
rect 419262 163200 419318 164400
rect 420090 163200 420146 164400
rect 420918 163200 420974 164400
rect 421746 163200 421802 164400
rect 422574 163200 422630 164400
rect 423402 163200 423458 164400
rect 424322 163200 424378 164400
rect 425150 163200 425206 164400
rect 425978 163200 426034 164400
rect 426084 163254 426388 163282
rect 415872 153202 415900 163200
rect 416596 159928 416648 159934
rect 416596 159870 416648 159876
rect 415860 153196 415912 153202
rect 415860 153138 415912 153144
rect 415308 153128 415360 153134
rect 415308 153070 415360 153076
rect 416608 151978 416636 159870
rect 416700 158982 416728 163200
rect 417528 159390 417556 163200
rect 417884 159724 417936 159730
rect 417884 159666 417936 159672
rect 417516 159384 417568 159390
rect 417516 159326 417568 159332
rect 416688 158976 416740 158982
rect 416688 158918 416740 158924
rect 417148 154352 417200 154358
rect 417148 154294 417200 154300
rect 416504 151972 416556 151978
rect 416504 151914 416556 151920
rect 416596 151972 416648 151978
rect 416596 151914 416648 151920
rect 415860 151904 415912 151910
rect 415860 151846 415912 151852
rect 415872 150226 415900 151846
rect 416516 150226 416544 151914
rect 417160 150226 417188 154294
rect 417896 152250 417924 159666
rect 418448 152454 418476 163200
rect 419276 152590 419304 163200
rect 420104 158982 420132 163200
rect 420932 159730 420960 163200
rect 420920 159724 420972 159730
rect 420920 159666 420972 159672
rect 419540 158976 419592 158982
rect 419540 158918 419592 158924
rect 420092 158976 420144 158982
rect 420092 158918 420144 158924
rect 419080 152584 419132 152590
rect 419080 152526 419132 152532
rect 419264 152584 419316 152590
rect 419264 152526 419316 152532
rect 418436 152448 418488 152454
rect 418436 152390 418488 152396
rect 417792 152244 417844 152250
rect 417792 152186 417844 152192
rect 417884 152244 417936 152250
rect 417884 152186 417936 152192
rect 417804 150226 417832 152186
rect 418436 152040 418488 152046
rect 418436 151982 418488 151988
rect 418448 150226 418476 151982
rect 419092 150226 419120 152526
rect 419552 151978 419580 158918
rect 419632 158772 419684 158778
rect 419632 158714 419684 158720
rect 419540 151972 419592 151978
rect 419540 151914 419592 151920
rect 419644 151842 419672 158714
rect 419724 154284 419776 154290
rect 419724 154226 419776 154232
rect 419632 151836 419684 151842
rect 419632 151778 419684 151784
rect 419736 150226 419764 154226
rect 421760 152794 421788 163200
rect 422300 154012 422352 154018
rect 422300 153954 422352 153960
rect 420368 152788 420420 152794
rect 420368 152730 420420 152736
rect 421748 152788 421800 152794
rect 421748 152730 421800 152736
rect 420380 150226 420408 152730
rect 421748 152244 421800 152250
rect 421748 152186 421800 152192
rect 421012 152108 421064 152114
rect 421012 152050 421064 152056
rect 421024 150226 421052 152050
rect 421760 151910 421788 152186
rect 421656 151904 421708 151910
rect 421656 151846 421708 151852
rect 421748 151904 421800 151910
rect 421748 151846 421800 151852
rect 421668 150226 421696 151846
rect 422312 150226 422340 153954
rect 422588 152046 422616 163200
rect 423036 154420 423088 154426
rect 423036 154362 423088 154368
rect 422576 152040 422628 152046
rect 422576 151982 422628 151988
rect 423048 150226 423076 154362
rect 423416 152250 423444 163200
rect 424336 159798 424364 163200
rect 424324 159792 424376 159798
rect 424324 159734 424376 159740
rect 423588 158976 423640 158982
rect 423588 158918 423640 158924
rect 423600 152318 423628 158918
rect 424876 154488 424928 154494
rect 424876 154430 424928 154436
rect 424232 152856 424284 152862
rect 424232 152798 424284 152804
rect 423588 152312 423640 152318
rect 423588 152254 423640 152260
rect 423404 152244 423456 152250
rect 423404 152186 423456 152192
rect 423588 152176 423640 152182
rect 423588 152118 423640 152124
rect 412008 150198 412082 150226
rect 412652 150198 412726 150226
rect 413296 150198 413370 150226
rect 413940 150198 414014 150226
rect 414584 150198 414658 150226
rect 415228 150198 415302 150226
rect 415872 150198 415946 150226
rect 416516 150198 416590 150226
rect 417160 150198 417234 150226
rect 417804 150198 417878 150226
rect 418448 150198 418522 150226
rect 419092 150198 419166 150226
rect 419736 150198 419810 150226
rect 420380 150198 420454 150226
rect 421024 150198 421098 150226
rect 421668 150198 421742 150226
rect 422312 150198 422386 150226
rect 411410 149940 411438 150198
rect 412054 149940 412082 150198
rect 412698 149940 412726 150198
rect 413342 149940 413370 150198
rect 413986 149940 414014 150198
rect 414630 149940 414658 150198
rect 415274 149940 415302 150198
rect 415918 149940 415946 150198
rect 416562 149940 416590 150198
rect 417206 149940 417234 150198
rect 417850 149940 417878 150198
rect 418494 149940 418522 150198
rect 419138 149940 419166 150198
rect 419782 149940 419810 150198
rect 420426 149940 420454 150198
rect 421070 149940 421098 150198
rect 421714 149940 421742 150198
rect 422358 149940 422386 150198
rect 423002 150198 423076 150226
rect 423600 150226 423628 152118
rect 424244 150226 424272 152798
rect 424888 150226 424916 154430
rect 425164 152862 425192 163200
rect 425992 163146 426020 163200
rect 426084 163146 426112 163254
rect 425992 163118 426112 163146
rect 425520 155236 425572 155242
rect 425520 155178 425572 155184
rect 425152 152856 425204 152862
rect 425152 152798 425204 152804
rect 425532 150226 425560 155178
rect 426164 152924 426216 152930
rect 426164 152866 426216 152872
rect 426256 152924 426308 152930
rect 426256 152866 426308 152872
rect 426176 150226 426204 152866
rect 426268 152318 426296 152866
rect 426360 152318 426388 163254
rect 426806 163200 426862 164400
rect 427634 163200 427690 164400
rect 428462 163200 428518 164400
rect 429290 163200 429346 164400
rect 430210 163200 430266 164400
rect 430316 163254 430528 163282
rect 426820 161474 426848 163200
rect 426820 161446 426940 161474
rect 426256 152312 426308 152318
rect 426256 152254 426308 152260
rect 426348 152312 426400 152318
rect 426348 152254 426400 152260
rect 426912 152114 426940 161446
rect 427360 160064 427412 160070
rect 427360 160006 427412 160012
rect 427176 152924 427228 152930
rect 427176 152866 427228 152872
rect 427188 152726 427216 152866
rect 427084 152720 427136 152726
rect 427084 152662 427136 152668
rect 427176 152720 427228 152726
rect 427176 152662 427228 152668
rect 427096 152182 427124 152662
rect 427084 152176 427136 152182
rect 427084 152118 427136 152124
rect 426808 152108 426860 152114
rect 426808 152050 426860 152056
rect 426900 152108 426952 152114
rect 426900 152050 426952 152056
rect 426820 150226 426848 152050
rect 427372 150226 427400 160006
rect 427648 159458 427676 163200
rect 427636 159452 427688 159458
rect 427636 159394 427688 159400
rect 428476 152658 428504 163200
rect 429304 152998 429332 163200
rect 430224 163146 430252 163200
rect 430316 163146 430344 163254
rect 430224 163118 430344 163146
rect 429936 159520 429988 159526
rect 429936 159462 429988 159468
rect 429200 152992 429252 152998
rect 429200 152934 429252 152940
rect 429292 152992 429344 152998
rect 429292 152934 429344 152940
rect 428004 152652 428056 152658
rect 428004 152594 428056 152600
rect 428464 152652 428516 152658
rect 428464 152594 428516 152600
rect 428016 150226 428044 152594
rect 428648 152380 428700 152386
rect 428648 152322 428700 152328
rect 428660 150226 428688 152322
rect 429212 151814 429240 152934
rect 429212 151786 429332 151814
rect 429304 150226 429332 151786
rect 429948 150226 429976 159462
rect 430500 152930 430528 163254
rect 431038 163200 431094 164400
rect 431866 163200 431922 164400
rect 432694 163200 432750 164400
rect 433522 163200 433578 164400
rect 434350 163200 434406 164400
rect 434456 163254 434668 163282
rect 430488 152924 430540 152930
rect 430488 152866 430540 152872
rect 430578 152416 430634 152425
rect 431052 152386 431080 163200
rect 431592 152720 431644 152726
rect 431592 152662 431644 152668
rect 431224 152516 431276 152522
rect 431224 152458 431276 152464
rect 431316 152516 431368 152522
rect 431316 152458 431368 152464
rect 430578 152351 430634 152360
rect 431040 152380 431092 152386
rect 430592 150226 430620 152351
rect 431040 152322 431092 152328
rect 431236 150226 431264 152458
rect 431328 152318 431356 152458
rect 431316 152312 431368 152318
rect 431316 152254 431368 152260
rect 431500 152244 431552 152250
rect 431500 152186 431552 152192
rect 431512 152046 431540 152186
rect 431604 152046 431632 152662
rect 431880 152425 431908 163200
rect 432512 159588 432564 159594
rect 432512 159530 432564 159536
rect 431866 152416 431922 152425
rect 431866 152351 431922 152360
rect 431500 152040 431552 152046
rect 431500 151982 431552 151988
rect 431592 152040 431644 152046
rect 431592 151982 431644 151988
rect 431868 151904 431920 151910
rect 431868 151846 431920 151852
rect 431880 150226 431908 151846
rect 432524 150226 432552 159530
rect 432708 153066 432736 163200
rect 433064 153264 433116 153270
rect 433116 153212 433288 153218
rect 433064 153206 433288 153212
rect 433076 153190 433288 153206
rect 433260 153134 433288 153190
rect 433156 153128 433208 153134
rect 433156 153070 433208 153076
rect 433248 153128 433300 153134
rect 433248 153070 433300 153076
rect 432696 153060 432748 153066
rect 432696 153002 432748 153008
rect 433168 150226 433196 153070
rect 433340 152788 433392 152794
rect 433340 152730 433392 152736
rect 433432 152788 433484 152794
rect 433432 152730 433484 152736
rect 433352 151910 433380 152730
rect 433444 152590 433472 152730
rect 433536 152590 433564 163200
rect 434364 163146 434392 163200
rect 434456 163146 434484 163254
rect 434364 163118 434484 163146
rect 434640 152726 434668 163254
rect 435178 163200 435234 164400
rect 436098 163200 436154 164400
rect 436926 163200 436982 164400
rect 437032 163254 437336 163282
rect 435088 159656 435140 159662
rect 435088 159598 435140 159604
rect 434628 152720 434680 152726
rect 434628 152662 434680 152668
rect 433432 152584 433484 152590
rect 433432 152526 433484 152532
rect 433524 152584 433576 152590
rect 433524 152526 433576 152532
rect 433800 152176 433852 152182
rect 433800 152118 433852 152124
rect 433340 151904 433392 151910
rect 433340 151846 433392 151852
rect 433812 150226 433840 152118
rect 434444 151836 434496 151842
rect 434444 151778 434496 151784
rect 434456 150226 434484 151778
rect 435100 150226 435128 159598
rect 435192 158778 435220 163200
rect 435180 158772 435232 158778
rect 435180 158714 435232 158720
rect 435824 158772 435876 158778
rect 435824 158714 435876 158720
rect 435836 153202 435864 158714
rect 435732 153196 435784 153202
rect 435732 153138 435784 153144
rect 435824 153196 435876 153202
rect 435824 153138 435876 153144
rect 435744 150226 435772 153138
rect 436112 151910 436140 163200
rect 436940 163146 436968 163200
rect 437032 163146 437060 163254
rect 436940 163118 437060 163146
rect 437308 153202 437336 163254
rect 437754 163200 437810 164400
rect 438582 163200 438638 164400
rect 439410 163200 439466 164400
rect 440238 163200 440294 164400
rect 441066 163200 441122 164400
rect 441172 163254 441476 163282
rect 437664 159384 437716 159390
rect 437664 159326 437716 159332
rect 437296 153196 437348 153202
rect 437296 153138 437348 153144
rect 436376 153128 436428 153134
rect 436376 153070 436428 153076
rect 436100 151904 436152 151910
rect 436100 151846 436152 151852
rect 436388 150226 436416 153070
rect 436744 152516 436796 152522
rect 436744 152458 436796 152464
rect 436756 152182 436784 152458
rect 436744 152176 436796 152182
rect 436744 152118 436796 152124
rect 437020 151972 437072 151978
rect 437020 151914 437072 151920
rect 437032 150226 437060 151914
rect 437676 150226 437704 159326
rect 437768 152454 437796 163200
rect 438596 153134 438624 163200
rect 438492 153128 438544 153134
rect 438492 153070 438544 153076
rect 438584 153128 438636 153134
rect 438584 153070 438636 153076
rect 438504 152590 438532 153070
rect 438952 152788 439004 152794
rect 438952 152730 439004 152736
rect 438492 152584 438544 152590
rect 438492 152526 438544 152532
rect 438308 152516 438360 152522
rect 438308 152458 438360 152464
rect 437756 152448 437808 152454
rect 437756 152390 437808 152396
rect 438320 150226 438348 152458
rect 438964 150226 438992 152730
rect 439424 151978 439452 163200
rect 439596 152040 439648 152046
rect 439596 151982 439648 151988
rect 439412 151972 439464 151978
rect 439412 151914 439464 151920
rect 439608 150226 439636 151982
rect 440252 151842 440280 163200
rect 441080 163146 441108 163200
rect 441172 163146 441200 163254
rect 441080 163118 441200 163146
rect 440332 159724 440384 159730
rect 440332 159666 440384 159672
rect 440240 151836 440292 151842
rect 440240 151778 440292 151784
rect 440344 150226 440372 159666
rect 441448 152590 441476 163254
rect 441986 163200 442042 164400
rect 442814 163200 442870 164400
rect 443642 163200 443698 164400
rect 444470 163200 444526 164400
rect 445298 163200 445354 164400
rect 445404 163254 445708 163282
rect 440976 152584 441028 152590
rect 440976 152526 441028 152532
rect 441436 152584 441488 152590
rect 441436 152526 441488 152532
rect 440988 151910 441016 152526
rect 442000 152250 442028 163200
rect 442724 159792 442776 159798
rect 442724 159734 442776 159740
rect 442172 152312 442224 152318
rect 442172 152254 442224 152260
rect 441528 152244 441580 152250
rect 441528 152186 441580 152192
rect 441988 152244 442040 152250
rect 441988 152186 442040 152192
rect 440884 151904 440936 151910
rect 440884 151846 440936 151852
rect 440976 151904 441028 151910
rect 440976 151846 441028 151852
rect 423600 150198 423674 150226
rect 424244 150198 424318 150226
rect 424888 150198 424962 150226
rect 425532 150198 425606 150226
rect 426176 150198 426250 150226
rect 426820 150198 426894 150226
rect 427372 150198 427446 150226
rect 428016 150198 428090 150226
rect 428660 150198 428734 150226
rect 429304 150198 429378 150226
rect 429948 150198 430022 150226
rect 430592 150198 430666 150226
rect 431236 150198 431310 150226
rect 431880 150198 431954 150226
rect 432524 150198 432598 150226
rect 433168 150198 433242 150226
rect 433812 150198 433886 150226
rect 434456 150198 434530 150226
rect 435100 150198 435174 150226
rect 435744 150198 435818 150226
rect 436388 150198 436462 150226
rect 437032 150198 437106 150226
rect 437676 150198 437750 150226
rect 438320 150198 438394 150226
rect 438964 150198 439038 150226
rect 439608 150198 439682 150226
rect 423002 149940 423030 150198
rect 423646 149940 423674 150198
rect 424290 149940 424318 150198
rect 424934 149940 424962 150198
rect 425578 149940 425606 150198
rect 426222 149940 426250 150198
rect 426866 149940 426894 150198
rect 427418 149940 427446 150198
rect 428062 149940 428090 150198
rect 428706 149940 428734 150198
rect 429350 149940 429378 150198
rect 429994 149940 430022 150198
rect 430638 149940 430666 150198
rect 431282 149940 431310 150198
rect 431926 149940 431954 150198
rect 432570 149940 432598 150198
rect 433214 149940 433242 150198
rect 433858 149940 433886 150198
rect 434502 149940 434530 150198
rect 435146 149940 435174 150198
rect 435790 149940 435818 150198
rect 436434 149940 436462 150198
rect 437078 149940 437106 150198
rect 437722 149940 437750 150198
rect 438366 149940 438394 150198
rect 439010 149940 439038 150198
rect 439654 149940 439682 150198
rect 440298 150198 440372 150226
rect 440896 150226 440924 151846
rect 441540 150226 441568 152186
rect 442184 150226 442212 152254
rect 442736 151814 442764 159734
rect 442828 152794 442856 163200
rect 443460 152856 443512 152862
rect 443460 152798 443512 152804
rect 442816 152788 442868 152794
rect 442816 152730 442868 152736
rect 442736 151786 442856 151814
rect 442828 150226 442856 151786
rect 443472 150226 443500 152798
rect 443656 152250 443684 163200
rect 444484 152862 444512 163200
rect 445312 163146 445340 163200
rect 445404 163146 445432 163254
rect 445312 163118 445432 163146
rect 445392 159452 445444 159458
rect 445392 159394 445444 159400
rect 444472 152856 444524 152862
rect 444472 152798 444524 152804
rect 443644 152244 443696 152250
rect 443644 152186 443696 152192
rect 444104 152176 444156 152182
rect 444104 152118 444156 152124
rect 444116 150226 444144 152118
rect 444748 152108 444800 152114
rect 444748 152050 444800 152056
rect 444760 150226 444788 152050
rect 445404 150226 445432 159394
rect 445680 152182 445708 163254
rect 446126 163200 446182 164400
rect 446954 163200 447010 164400
rect 447874 163200 447930 164400
rect 448702 163200 448758 164400
rect 449530 163200 449586 164400
rect 450358 163200 450414 164400
rect 451186 163200 451242 164400
rect 452014 163200 452070 164400
rect 452842 163200 452898 164400
rect 453762 163200 453818 164400
rect 454590 163200 454646 164400
rect 455418 163200 455474 164400
rect 456246 163200 456302 164400
rect 457074 163200 457130 164400
rect 457902 163200 457958 164400
rect 458730 163200 458786 164400
rect 459650 163200 459706 164400
rect 460478 163200 460534 164400
rect 461306 163200 461362 164400
rect 462134 163200 462190 164400
rect 462962 163200 463018 164400
rect 463790 163200 463846 164400
rect 464618 163200 464674 164400
rect 465538 163200 465594 164400
rect 466366 163200 466422 164400
rect 467194 163200 467250 164400
rect 468022 163200 468078 164400
rect 468850 163200 468906 164400
rect 469678 163200 469734 164400
rect 470506 163200 470562 164400
rect 471426 163200 471482 164400
rect 472254 163200 472310 164400
rect 473082 163200 473138 164400
rect 473910 163200 473966 164400
rect 474738 163200 474794 164400
rect 475566 163200 475622 164400
rect 476394 163200 476450 164400
rect 477314 163200 477370 164400
rect 478142 163200 478198 164400
rect 478970 163200 479026 164400
rect 479798 163200 479854 164400
rect 480626 163200 480682 164400
rect 481454 163200 481510 164400
rect 482282 163200 482338 164400
rect 483202 163200 483258 164400
rect 484030 163200 484086 164400
rect 484858 163200 484914 164400
rect 485686 163200 485742 164400
rect 486514 163200 486570 164400
rect 487342 163200 487398 164400
rect 488170 163200 488226 164400
rect 488276 163254 488488 163282
rect 446140 158914 446168 163200
rect 446128 158908 446180 158914
rect 446128 158850 446180 158856
rect 446680 152992 446732 152998
rect 446680 152934 446732 152940
rect 446036 152652 446088 152658
rect 446036 152594 446088 152600
rect 445668 152176 445720 152182
rect 445668 152118 445720 152124
rect 446048 150226 446076 152594
rect 446692 150226 446720 152934
rect 446968 152658 446996 163200
rect 447888 159390 447916 163200
rect 448716 159594 448744 163200
rect 448704 159588 448756 159594
rect 448704 159530 448756 159536
rect 449544 159526 449572 163200
rect 450372 159934 450400 163200
rect 450360 159928 450412 159934
rect 450360 159870 450412 159876
rect 449532 159520 449584 159526
rect 449532 159462 449584 159468
rect 451200 159458 451228 163200
rect 451188 159452 451240 159458
rect 451188 159394 451240 159400
rect 447876 159384 447928 159390
rect 447876 159326 447928 159332
rect 452028 158846 452056 163200
rect 452016 158840 452068 158846
rect 452016 158782 452068 158788
rect 452856 158778 452884 163200
rect 453776 159390 453804 163200
rect 453764 159384 453816 159390
rect 453764 159326 453816 159332
rect 454604 158982 454632 163200
rect 455432 159050 455460 163200
rect 456064 159588 456116 159594
rect 456064 159530 456116 159536
rect 455788 159520 455840 159526
rect 455788 159462 455840 159468
rect 455420 159044 455472 159050
rect 455420 158986 455472 158992
rect 454592 158976 454644 158982
rect 454592 158918 454644 158924
rect 453948 158908 454000 158914
rect 453948 158850 454000 158856
rect 452844 158772 452896 158778
rect 452844 158714 452896 158720
rect 453960 153202 453988 158850
rect 452476 153196 452528 153202
rect 452476 153138 452528 153144
rect 453948 153196 454000 153202
rect 453948 153138 454000 153144
rect 449256 153060 449308 153066
rect 449256 153002 449308 153008
rect 447324 152924 447376 152930
rect 447324 152866 447376 152872
rect 446956 152652 447008 152658
rect 446956 152594 447008 152600
rect 447336 150226 447364 152866
rect 448610 152416 448666 152425
rect 447968 152380 448020 152386
rect 448610 152351 448666 152360
rect 447968 152322 448020 152328
rect 447980 150226 448008 152322
rect 448624 150226 448652 152351
rect 449268 150226 449296 153002
rect 450544 152720 450596 152726
rect 450544 152662 450596 152668
rect 449900 152516 449952 152522
rect 449900 152458 449952 152464
rect 449912 150226 449940 152458
rect 450556 150226 450584 152662
rect 451832 151972 451884 151978
rect 451832 151914 451884 151920
rect 451188 151904 451240 151910
rect 451188 151846 451240 151852
rect 451200 150226 451228 151846
rect 451844 150226 451872 151914
rect 452488 150226 452516 153138
rect 453764 153128 453816 153134
rect 453764 153070 453816 153076
rect 453120 152448 453172 152454
rect 453120 152390 453172 152396
rect 453132 150226 453160 152390
rect 453776 150226 453804 153070
rect 455696 152584 455748 152590
rect 455696 152526 455748 152532
rect 454408 152040 454460 152046
rect 454408 151982 454460 151988
rect 454420 150226 454448 151982
rect 455052 151836 455104 151842
rect 455052 151778 455104 151784
rect 455064 150226 455092 151778
rect 455708 150226 455736 152526
rect 455800 151842 455828 159462
rect 456076 151978 456104 159530
rect 456260 158914 456288 163200
rect 457088 159526 457116 163200
rect 457168 159928 457220 159934
rect 457168 159870 457220 159876
rect 457076 159520 457128 159526
rect 457076 159462 457128 159468
rect 456800 159452 456852 159458
rect 456800 159394 456852 159400
rect 456248 158908 456300 158914
rect 456248 158850 456300 158856
rect 456340 152312 456392 152318
rect 456340 152254 456392 152260
rect 456064 151972 456116 151978
rect 456064 151914 456116 151920
rect 455788 151836 455840 151842
rect 455788 151778 455840 151784
rect 456352 150226 456380 152254
rect 456812 152046 456840 159394
rect 456892 159316 456944 159322
rect 456892 159258 456944 159264
rect 456904 153134 456932 159258
rect 456892 153128 456944 153134
rect 456892 153070 456944 153076
rect 456984 152788 457036 152794
rect 456984 152730 457036 152736
rect 456800 152040 456852 152046
rect 456800 151982 456852 151988
rect 456996 150226 457024 152730
rect 457180 151910 457208 159870
rect 457916 159322 457944 163200
rect 458744 159934 458772 163200
rect 458732 159928 458784 159934
rect 458732 159870 458784 159876
rect 459664 159662 459692 163200
rect 459652 159656 459704 159662
rect 459652 159598 459704 159604
rect 460492 159594 460520 163200
rect 460480 159588 460532 159594
rect 460480 159530 460532 159536
rect 459652 159384 459704 159390
rect 459652 159326 459704 159332
rect 457904 159316 457956 159322
rect 457904 159258 457956 159264
rect 458180 158840 458232 158846
rect 458180 158782 458232 158788
rect 458192 152726 458220 158782
rect 459560 158772 459612 158778
rect 459560 158714 459612 158720
rect 459468 153196 459520 153202
rect 459468 153138 459520 153144
rect 458272 152856 458324 152862
rect 458272 152798 458324 152804
rect 458180 152720 458232 152726
rect 458180 152662 458232 152668
rect 457628 152244 457680 152250
rect 457628 152186 457680 152192
rect 457168 151904 457220 151910
rect 457168 151846 457220 151852
rect 457640 150226 457668 152186
rect 458284 150226 458312 152798
rect 458824 152176 458876 152182
rect 458824 152118 458876 152124
rect 440896 150198 440970 150226
rect 441540 150198 441614 150226
rect 442184 150198 442258 150226
rect 442828 150198 442902 150226
rect 443472 150198 443546 150226
rect 444116 150198 444190 150226
rect 444760 150198 444834 150226
rect 445404 150198 445478 150226
rect 446048 150198 446122 150226
rect 446692 150198 446766 150226
rect 447336 150198 447410 150226
rect 447980 150198 448054 150226
rect 448624 150198 448698 150226
rect 449268 150198 449342 150226
rect 449912 150198 449986 150226
rect 450556 150198 450630 150226
rect 451200 150198 451274 150226
rect 451844 150198 451918 150226
rect 452488 150198 452562 150226
rect 453132 150198 453206 150226
rect 453776 150198 453850 150226
rect 454420 150198 454494 150226
rect 455064 150198 455138 150226
rect 455708 150198 455782 150226
rect 456352 150198 456426 150226
rect 456996 150198 457070 150226
rect 457640 150198 457714 150226
rect 440298 149940 440326 150198
rect 440942 149940 440970 150198
rect 441586 149940 441614 150198
rect 442230 149940 442258 150198
rect 442874 149940 442902 150198
rect 443518 149940 443546 150198
rect 444162 149940 444190 150198
rect 444806 149940 444834 150198
rect 445450 149940 445478 150198
rect 446094 149940 446122 150198
rect 446738 149940 446766 150198
rect 447382 149940 447410 150198
rect 448026 149940 448054 150198
rect 448670 149940 448698 150198
rect 449314 149940 449342 150198
rect 449958 149940 449986 150198
rect 450602 149940 450630 150198
rect 451246 149940 451274 150198
rect 451890 149940 451918 150198
rect 452534 149940 452562 150198
rect 453178 149940 453206 150198
rect 453822 149940 453850 150198
rect 454466 149940 454494 150198
rect 455110 149940 455138 150198
rect 455754 149940 455782 150198
rect 456398 149940 456426 150198
rect 457042 149940 457070 150198
rect 457686 149940 457714 150198
rect 458238 150198 458312 150226
rect 458836 150226 458864 152118
rect 459480 150226 459508 153138
rect 459572 152998 459600 158714
rect 459560 152992 459612 152998
rect 459560 152934 459612 152940
rect 459664 152658 459692 159326
rect 461320 159254 461348 163200
rect 461308 159248 461360 159254
rect 461308 159190 461360 159196
rect 462148 159186 462176 163200
rect 462136 159180 462188 159186
rect 462136 159122 462188 159128
rect 462976 159118 463004 163200
rect 462964 159112 463016 159118
rect 462964 159054 463016 159060
rect 463332 159044 463384 159050
rect 463332 158986 463384 158992
rect 461860 158976 461912 158982
rect 461860 158918 461912 158924
rect 461872 153202 461900 158918
rect 462964 158908 463016 158914
rect 462964 158850 463016 158856
rect 461860 153196 461912 153202
rect 461860 153138 461912 153144
rect 462976 153134 463004 158850
rect 460756 153128 460808 153134
rect 460756 153070 460808 153076
rect 462964 153128 463016 153134
rect 462964 153070 463016 153076
rect 459652 152652 459704 152658
rect 459652 152594 459704 152600
rect 460112 152584 460164 152590
rect 460112 152526 460164 152532
rect 460124 150226 460152 152526
rect 460768 150226 460796 153070
rect 463344 153066 463372 158986
rect 463804 158914 463832 163200
rect 464160 159520 464212 159526
rect 464160 159462 464212 159468
rect 463792 158908 463844 158914
rect 463792 158850 463844 158856
rect 463332 153060 463384 153066
rect 463332 153002 463384 153008
rect 464172 152930 464200 159462
rect 464528 159316 464580 159322
rect 464528 159258 464580 159264
rect 464160 152924 464212 152930
rect 464160 152866 464212 152872
rect 464540 152862 464568 159258
rect 464632 158846 464660 163200
rect 465080 159928 465132 159934
rect 465080 159870 465132 159876
rect 464620 158840 464672 158846
rect 464620 158782 464672 158788
rect 465092 152998 465120 159870
rect 465552 158778 465580 163200
rect 466380 158982 466408 163200
rect 467208 159866 467236 163200
rect 467196 159860 467248 159866
rect 467196 159802 467248 159808
rect 468036 159662 468064 163200
rect 466460 159656 466512 159662
rect 466460 159598 466512 159604
rect 468024 159656 468076 159662
rect 468024 159598 468076 159604
rect 466368 158976 466420 158982
rect 466368 158918 466420 158924
rect 465540 158772 465592 158778
rect 465540 158714 465592 158720
rect 466472 153202 466500 159598
rect 466644 159588 466696 159594
rect 466644 159530 466696 159536
rect 465908 153196 465960 153202
rect 465908 153138 465960 153144
rect 466460 153196 466512 153202
rect 466460 153138 466512 153144
rect 464620 152992 464672 152998
rect 464620 152934 464672 152940
rect 465080 152992 465132 152998
rect 465080 152934 465132 152940
rect 464528 152856 464580 152862
rect 464528 152798 464580 152804
rect 463976 152720 464028 152726
rect 463976 152662 464028 152668
rect 463332 152040 463384 152046
rect 463332 151982 463384 151988
rect 461400 151972 461452 151978
rect 461400 151914 461452 151920
rect 461412 150226 461440 151914
rect 462688 151904 462740 151910
rect 462688 151846 462740 151852
rect 462044 151836 462096 151842
rect 462044 151778 462096 151784
rect 462056 150226 462084 151778
rect 462700 150226 462728 151846
rect 463344 150226 463372 151982
rect 463988 150226 464016 152662
rect 464632 150226 464660 152934
rect 465264 152652 465316 152658
rect 465264 152594 465316 152600
rect 465276 150226 465304 152594
rect 465920 150226 465948 153138
rect 466656 153066 466684 159530
rect 468864 159526 468892 163200
rect 468852 159520 468904 159526
rect 468852 159462 468904 159468
rect 469692 159390 469720 163200
rect 470520 159594 470548 163200
rect 471440 159798 471468 163200
rect 471428 159792 471480 159798
rect 471428 159734 471480 159740
rect 470508 159588 470560 159594
rect 470508 159530 470560 159536
rect 469680 159384 469732 159390
rect 469680 159326 469732 159332
rect 468024 159248 468076 159254
rect 468024 159190 468076 159196
rect 467932 159180 467984 159186
rect 467932 159122 467984 159128
rect 467196 153128 467248 153134
rect 467196 153070 467248 153076
rect 466552 153060 466604 153066
rect 466552 153002 466604 153008
rect 466644 153060 466696 153066
rect 466644 153002 466696 153008
rect 466564 150226 466592 153002
rect 467208 150226 467236 153070
rect 467840 152924 467892 152930
rect 467840 152866 467892 152872
rect 467852 150226 467880 152866
rect 467944 151842 467972 159122
rect 468036 151910 468064 159190
rect 472268 159118 472296 163200
rect 469220 159112 469272 159118
rect 469220 159054 469272 159060
rect 472256 159112 472308 159118
rect 472256 159054 472308 159060
rect 469128 152992 469180 152998
rect 469128 152934 469180 152940
rect 468392 152856 468444 152862
rect 468392 152798 468444 152804
rect 468024 151904 468076 151910
rect 468024 151846 468076 151852
rect 467932 151836 467984 151842
rect 468404 151814 468432 152798
rect 468404 151786 468524 151814
rect 467932 151778 467984 151784
rect 468496 150226 468524 151786
rect 469140 150226 469168 152934
rect 469232 151978 469260 159054
rect 472532 158976 472584 158982
rect 472532 158918 472584 158924
rect 471244 158908 471296 158914
rect 471244 158850 471296 158856
rect 471256 153202 471284 158850
rect 471612 158840 471664 158846
rect 471612 158782 471664 158788
rect 469772 153196 469824 153202
rect 469772 153138 469824 153144
rect 471244 153196 471296 153202
rect 471244 153138 471296 153144
rect 469220 151972 469272 151978
rect 469220 151914 469272 151920
rect 469784 150226 469812 153138
rect 471624 153134 471652 158782
rect 472440 158772 472492 158778
rect 472440 158714 472492 158720
rect 471612 153128 471664 153134
rect 471612 153070 471664 153076
rect 472452 153066 472480 158714
rect 470416 153060 470468 153066
rect 470416 153002 470468 153008
rect 472440 153060 472492 153066
rect 472440 153002 472492 153008
rect 470428 150226 470456 153002
rect 472544 152998 472572 158918
rect 473096 158778 473124 163200
rect 473360 159860 473412 159866
rect 473360 159802 473412 159808
rect 473084 158772 473136 158778
rect 473084 158714 473136 158720
rect 472992 153196 473044 153202
rect 472992 153138 473044 153144
rect 472532 152992 472584 152998
rect 472532 152934 472584 152940
rect 472348 151972 472400 151978
rect 472348 151914 472400 151920
rect 471060 151904 471112 151910
rect 471060 151846 471112 151852
rect 471072 150226 471100 151846
rect 471704 151836 471756 151842
rect 471704 151778 471756 151784
rect 471716 150226 471744 151778
rect 472360 150226 472388 151914
rect 473004 150226 473032 153138
rect 473372 152930 473400 159802
rect 473924 159050 473952 163200
rect 473912 159044 473964 159050
rect 473912 158986 473964 158992
rect 474752 158914 474780 163200
rect 474832 159520 474884 159526
rect 474832 159462 474884 159468
rect 474740 158908 474792 158914
rect 474740 158850 474792 158856
rect 474844 153202 474872 159462
rect 475580 158982 475608 163200
rect 476028 159656 476080 159662
rect 476028 159598 476080 159604
rect 475568 158976 475620 158982
rect 475568 158918 475620 158924
rect 474832 153196 474884 153202
rect 474832 153138 474884 153144
rect 473636 153128 473688 153134
rect 473636 153070 473688 153076
rect 473360 152924 473412 152930
rect 473360 152866 473412 152872
rect 473648 150226 473676 153070
rect 474280 153060 474332 153066
rect 474280 153002 474332 153008
rect 474292 150226 474320 153002
rect 474924 152992 474976 152998
rect 474924 152934 474976 152940
rect 474936 150226 474964 152934
rect 475568 152924 475620 152930
rect 475568 152866 475620 152872
rect 475580 150226 475608 152866
rect 476040 151814 476068 159598
rect 476120 159588 476172 159594
rect 476120 159530 476172 159536
rect 476132 153134 476160 159530
rect 476408 158846 476436 163200
rect 477328 159526 477356 163200
rect 477684 159792 477736 159798
rect 477684 159734 477736 159740
rect 477316 159520 477368 159526
rect 477316 159462 477368 159468
rect 477408 159384 477460 159390
rect 477408 159326 477460 159332
rect 476396 158840 476448 158846
rect 476396 158782 476448 158788
rect 476856 153196 476908 153202
rect 476856 153138 476908 153144
rect 476120 153128 476172 153134
rect 476120 153070 476172 153076
rect 476040 151786 476252 151814
rect 476224 150226 476252 151786
rect 476868 150226 476896 153138
rect 477420 151814 477448 159326
rect 477420 151786 477540 151814
rect 477512 150226 477540 151786
rect 458836 150198 458910 150226
rect 459480 150198 459554 150226
rect 460124 150198 460198 150226
rect 460768 150198 460842 150226
rect 461412 150198 461486 150226
rect 462056 150198 462130 150226
rect 462700 150198 462774 150226
rect 463344 150198 463418 150226
rect 463988 150198 464062 150226
rect 464632 150198 464706 150226
rect 465276 150198 465350 150226
rect 465920 150198 465994 150226
rect 466564 150198 466638 150226
rect 467208 150198 467282 150226
rect 467852 150198 467926 150226
rect 468496 150198 468570 150226
rect 469140 150198 469214 150226
rect 469784 150198 469858 150226
rect 470428 150198 470502 150226
rect 471072 150198 471146 150226
rect 471716 150198 471790 150226
rect 472360 150198 472434 150226
rect 473004 150198 473078 150226
rect 473648 150198 473722 150226
rect 474292 150198 474366 150226
rect 474936 150198 475010 150226
rect 475580 150198 475654 150226
rect 476224 150198 476298 150226
rect 476868 150198 476942 150226
rect 477512 150198 477586 150226
rect 477696 150210 477724 159734
rect 478156 159390 478184 163200
rect 478984 159934 479012 163200
rect 478972 159928 479024 159934
rect 478972 159870 479024 159876
rect 479812 159594 479840 163200
rect 479800 159588 479852 159594
rect 479800 159530 479852 159536
rect 478144 159384 478196 159390
rect 478144 159326 478196 159332
rect 479432 159112 479484 159118
rect 479432 159054 479484 159060
rect 478972 158772 479024 158778
rect 478972 158714 479024 158720
rect 478144 153128 478196 153134
rect 478144 153070 478196 153076
rect 478156 150226 478184 153070
rect 458238 149940 458266 150198
rect 458882 149940 458910 150198
rect 459526 149940 459554 150198
rect 460170 149940 460198 150198
rect 460814 149940 460842 150198
rect 461458 149940 461486 150198
rect 462102 149940 462130 150198
rect 462746 149940 462774 150198
rect 463390 149940 463418 150198
rect 464034 149940 464062 150198
rect 464678 149940 464706 150198
rect 465322 149940 465350 150198
rect 465966 149940 465994 150198
rect 466610 149940 466638 150198
rect 467254 149940 467282 150198
rect 467898 149940 467926 150198
rect 468542 149940 468570 150198
rect 469186 149940 469214 150198
rect 469830 149940 469858 150198
rect 470474 149940 470502 150198
rect 471118 149940 471146 150198
rect 471762 149940 471790 150198
rect 472406 149940 472434 150198
rect 473050 149940 473078 150198
rect 473694 149940 473722 150198
rect 474338 149940 474366 150198
rect 474982 149940 475010 150198
rect 475626 149940 475654 150198
rect 476270 149940 476298 150198
rect 476914 149940 476942 150198
rect 477558 149940 477586 150198
rect 477684 150204 477736 150210
rect 478156 150198 478230 150226
rect 478984 150210 479012 158714
rect 479444 150226 479472 159054
rect 480640 159050 480668 163200
rect 480260 159044 480312 159050
rect 480260 158986 480312 158992
rect 480628 159044 480680 159050
rect 480628 158986 480680 158992
rect 480272 151814 480300 158986
rect 481468 158914 481496 163200
rect 482008 158976 482060 158982
rect 482008 158918 482060 158924
rect 481364 158908 481416 158914
rect 481364 158850 481416 158856
rect 481456 158908 481508 158914
rect 481456 158850 481508 158856
rect 480272 151786 480760 151814
rect 480732 150226 480760 151786
rect 481376 150226 481404 158850
rect 481640 158840 481692 158846
rect 481640 158782 481692 158788
rect 477684 150146 477736 150152
rect 478202 149940 478230 150198
rect 478834 150204 478886 150210
rect 478834 150146 478886 150152
rect 478972 150204 479024 150210
rect 479444 150198 479518 150226
rect 478972 150146 479024 150152
rect 478846 149940 478874 150146
rect 479490 149940 479518 150198
rect 480122 150204 480174 150210
rect 480732 150198 480806 150226
rect 481376 150198 481450 150226
rect 481652 150210 481680 158782
rect 482020 150226 482048 158918
rect 482296 158778 482324 163200
rect 482284 158772 482336 158778
rect 482284 158714 482336 158720
rect 483216 152998 483244 163200
rect 483296 159520 483348 159526
rect 483296 159462 483348 159468
rect 483204 152992 483256 152998
rect 483204 152934 483256 152940
rect 483308 150226 483336 159462
rect 483940 159384 483992 159390
rect 483940 159326 483992 159332
rect 483952 150226 483980 159326
rect 484044 153066 484072 163200
rect 484584 159928 484636 159934
rect 484584 159870 484636 159876
rect 484032 153060 484084 153066
rect 484032 153002 484084 153008
rect 484596 150226 484624 159870
rect 484872 153134 484900 163200
rect 485228 159588 485280 159594
rect 485228 159530 485280 159536
rect 484860 153128 484912 153134
rect 484860 153070 484912 153076
rect 485240 150226 485268 159530
rect 485700 153202 485728 163200
rect 485872 159044 485924 159050
rect 485872 158986 485924 158992
rect 485688 153196 485740 153202
rect 485688 153138 485740 153144
rect 485884 150226 485912 158986
rect 486424 158908 486476 158914
rect 486424 158850 486476 158856
rect 486436 151814 486464 158850
rect 486528 152046 486556 163200
rect 487252 158772 487304 158778
rect 487252 158714 487304 158720
rect 486516 152040 486568 152046
rect 486516 151982 486568 151988
rect 486436 151786 486556 151814
rect 486528 150226 486556 151786
rect 487264 150226 487292 158714
rect 487356 151978 487384 163200
rect 488184 163146 488212 163200
rect 488276 163146 488304 163254
rect 488184 163118 488304 163146
rect 488356 153060 488408 153066
rect 488356 153002 488408 153008
rect 487804 152992 487856 152998
rect 487804 152934 487856 152940
rect 487344 151972 487396 151978
rect 487344 151914 487396 151920
rect 480122 150146 480174 150152
rect 480134 149940 480162 150146
rect 480778 149940 480806 150198
rect 481422 149940 481450 150198
rect 481640 150204 481692 150210
rect 482020 150198 482094 150226
rect 481640 150146 481692 150152
rect 482066 149940 482094 150198
rect 482698 150204 482750 150210
rect 483308 150198 483382 150226
rect 483952 150198 484026 150226
rect 484596 150198 484670 150226
rect 485240 150198 485314 150226
rect 485884 150198 485958 150226
rect 486528 150198 486602 150226
rect 482698 150146 482750 150152
rect 482710 149940 482738 150146
rect 483354 149940 483382 150198
rect 483998 149940 484026 150198
rect 484642 149940 484670 150198
rect 485286 149940 485314 150198
rect 485930 149940 485958 150198
rect 486574 149940 486602 150198
rect 487218 150198 487292 150226
rect 487816 150226 487844 152934
rect 487816 150198 487890 150226
rect 487218 149940 487246 150198
rect 487862 149940 487890 150198
rect 488368 150192 488396 153002
rect 488460 151842 488488 163254
rect 489090 163200 489146 164400
rect 489918 163200 489974 164400
rect 490746 163200 490802 164400
rect 491574 163200 491630 164400
rect 492402 163200 492458 164400
rect 493230 163200 493286 164400
rect 494058 163200 494114 164400
rect 494978 163200 495034 164400
rect 495084 163254 495296 163282
rect 489000 153128 489052 153134
rect 489000 153070 489052 153076
rect 488448 151836 488500 151842
rect 488448 151778 488500 151784
rect 489012 150226 489040 153070
rect 489104 151910 489132 163200
rect 489644 153196 489696 153202
rect 489644 153138 489696 153144
rect 489092 151904 489144 151910
rect 489092 151846 489144 151852
rect 489656 150226 489684 153138
rect 489932 153134 489960 163200
rect 490760 153202 490788 163200
rect 490748 153196 490800 153202
rect 490748 153138 490800 153144
rect 489920 153128 489972 153134
rect 489920 153070 489972 153076
rect 491588 152998 491616 163200
rect 492416 153066 492444 163200
rect 493244 153134 493272 163200
rect 494072 153202 494100 163200
rect 494992 163146 495020 163200
rect 495084 163146 495112 163254
rect 494992 163118 495112 163146
rect 493508 153196 493560 153202
rect 493508 153138 493560 153144
rect 494060 153196 494112 153202
rect 494060 153138 494112 153144
rect 492864 153128 492916 153134
rect 492864 153070 492916 153076
rect 493232 153128 493284 153134
rect 493232 153070 493284 153076
rect 492404 153060 492456 153066
rect 492404 153002 492456 153008
rect 491576 152992 491628 152998
rect 491576 152934 491628 152940
rect 490288 152040 490340 152046
rect 490288 151982 490340 151988
rect 490300 150226 490328 151982
rect 490932 151972 490984 151978
rect 490932 151914 490984 151920
rect 490944 150226 490972 151914
rect 492220 151904 492272 151910
rect 492220 151846 492272 151852
rect 491576 151836 491628 151842
rect 491576 151778 491628 151784
rect 491588 150226 491616 151778
rect 492232 150226 492260 151846
rect 492876 150226 492904 153070
rect 493520 150226 493548 153138
rect 495268 153066 495296 163254
rect 495806 163200 495862 164400
rect 496634 163200 496690 164400
rect 497462 163200 497518 164400
rect 498290 163200 498346 164400
rect 499118 163200 499174 164400
rect 499224 163254 499528 163282
rect 495820 153134 495848 163200
rect 496648 153202 496676 163200
rect 496084 153196 496136 153202
rect 496084 153138 496136 153144
rect 496636 153196 496688 153202
rect 496636 153138 496688 153144
rect 495440 153128 495492 153134
rect 495440 153070 495492 153076
rect 495808 153128 495860 153134
rect 495808 153070 495860 153076
rect 494796 153060 494848 153066
rect 494796 153002 494848 153008
rect 495256 153060 495308 153066
rect 495256 153002 495308 153008
rect 494152 152992 494204 152998
rect 494152 152934 494204 152940
rect 494164 150226 494192 152934
rect 494808 150226 494836 153002
rect 495452 150226 495480 153070
rect 496096 150226 496124 153138
rect 497476 153134 497504 163200
rect 498304 153202 498332 163200
rect 499132 163146 499160 163200
rect 499224 163146 499252 163254
rect 499132 163118 499252 163146
rect 498016 153196 498068 153202
rect 498016 153138 498068 153144
rect 498292 153196 498344 153202
rect 498292 153138 498344 153144
rect 499304 153196 499356 153202
rect 499304 153138 499356 153144
rect 497372 153128 497424 153134
rect 497372 153070 497424 153076
rect 497464 153128 497516 153134
rect 497464 153070 497516 153076
rect 496636 153060 496688 153066
rect 496636 153002 496688 153008
rect 496648 151814 496676 153002
rect 496648 151786 496768 151814
rect 496740 150226 496768 151786
rect 497384 150226 497412 153070
rect 498028 150226 498056 153138
rect 498660 153128 498712 153134
rect 498660 153070 498712 153076
rect 498672 150226 498700 153070
rect 499316 150226 499344 153138
rect 499500 151910 499528 163254
rect 499946 163200 500002 164400
rect 500866 163200 500922 164400
rect 500972 163254 501644 163282
rect 499960 158846 499988 163200
rect 499948 158840 500000 158846
rect 499948 158782 500000 158788
rect 500592 158840 500644 158846
rect 500592 158782 500644 158788
rect 499488 151904 499540 151910
rect 499488 151846 499540 151852
rect 499948 151904 500000 151910
rect 499948 151846 500000 151852
rect 499960 150226 499988 151846
rect 500604 150226 500632 158782
rect 500880 151814 500908 163200
rect 500972 153202 501000 163254
rect 501616 163146 501644 163254
rect 501694 163200 501750 164400
rect 502522 163200 502578 164400
rect 503350 163200 503406 164400
rect 503824 163254 504128 163282
rect 501708 163146 501736 163200
rect 501616 163118 501736 163146
rect 500960 153196 501012 153202
rect 500960 153138 501012 153144
rect 501880 153196 501932 153202
rect 501880 153138 501932 153144
rect 500880 151786 501276 151814
rect 501248 150226 501276 151786
rect 501892 150226 501920 153138
rect 502536 150226 502564 163200
rect 503364 151814 503392 163200
rect 503272 151786 503392 151814
rect 503272 150226 503300 151786
rect 489012 150198 489086 150226
rect 489656 150198 489730 150226
rect 490300 150198 490374 150226
rect 490944 150198 491018 150226
rect 491588 150198 491662 150226
rect 492232 150198 492306 150226
rect 492876 150198 492950 150226
rect 493520 150198 493594 150226
rect 494164 150198 494238 150226
rect 494808 150198 494882 150226
rect 495452 150198 495526 150226
rect 496096 150198 496170 150226
rect 496740 150198 496814 150226
rect 497384 150198 497458 150226
rect 498028 150198 498102 150226
rect 498672 150198 498746 150226
rect 499316 150198 499390 150226
rect 499960 150198 500034 150226
rect 500604 150198 500678 150226
rect 501248 150198 501322 150226
rect 501892 150198 501966 150226
rect 502536 150198 502610 150226
rect 488368 150164 488534 150192
rect 488506 149940 488534 150164
rect 489058 149940 489086 150198
rect 489702 149940 489730 150198
rect 490346 149940 490374 150198
rect 490990 149940 491018 150198
rect 491634 149940 491662 150198
rect 492278 149940 492306 150198
rect 492922 149940 492950 150198
rect 493566 149940 493594 150198
rect 494210 149940 494238 150198
rect 494854 149940 494882 150198
rect 495498 149940 495526 150198
rect 496142 149940 496170 150198
rect 496786 149940 496814 150198
rect 497430 149940 497458 150198
rect 498074 149940 498102 150198
rect 498718 149940 498746 150198
rect 499362 149940 499390 150198
rect 500006 149940 500034 150198
rect 500650 149940 500678 150198
rect 501294 149940 501322 150198
rect 501938 149940 501966 150198
rect 502582 149940 502610 150198
rect 503226 150198 503300 150226
rect 503824 150226 503852 163254
rect 504100 163146 504128 163254
rect 504178 163200 504234 164400
rect 505006 163200 505062 164400
rect 505112 163254 505784 163282
rect 504192 163146 504220 163200
rect 504100 163118 504220 163146
rect 505020 158778 505048 163200
rect 504456 158772 504508 158778
rect 504456 158714 504508 158720
rect 505008 158772 505060 158778
rect 505008 158714 505060 158720
rect 504468 150226 504496 158714
rect 505112 150226 505140 163254
rect 505756 163146 505784 163254
rect 505834 163200 505890 164400
rect 506492 163254 506704 163282
rect 505848 163146 505876 163200
rect 505756 163118 505876 163146
rect 506296 158840 506348 158846
rect 506296 158782 506348 158788
rect 505836 158772 505888 158778
rect 505836 158714 505888 158720
rect 505848 150226 505876 158714
rect 506308 151814 506336 158782
rect 506492 158778 506520 163254
rect 506676 163146 506704 163254
rect 506754 163200 506810 164400
rect 507582 163200 507638 164400
rect 508410 163200 508466 164400
rect 509238 163200 509294 164400
rect 510066 163200 510122 164400
rect 510894 163200 510950 164400
rect 511722 163200 511778 164400
rect 512012 163254 512592 163282
rect 506768 163146 506796 163200
rect 506676 163118 506796 163146
rect 507124 159044 507176 159050
rect 507124 158986 507176 158992
rect 506480 158772 506532 158778
rect 506480 158714 506532 158720
rect 506308 151786 506428 151814
rect 503824 150198 503898 150226
rect 504468 150198 504542 150226
rect 505112 150198 505186 150226
rect 503226 149940 503254 150198
rect 503870 149940 503898 150198
rect 504514 149940 504542 150198
rect 505158 149940 505186 150198
rect 505802 150198 505876 150226
rect 506400 150226 506428 151786
rect 507136 150226 507164 158986
rect 507596 158846 507624 163200
rect 508424 159050 508452 163200
rect 508412 159044 508464 159050
rect 508412 158986 508464 158992
rect 508412 158908 508464 158914
rect 508412 158850 508464 158856
rect 507584 158840 507636 158846
rect 507584 158782 507636 158788
rect 507676 151972 507728 151978
rect 507676 151914 507728 151920
rect 506400 150198 506474 150226
rect 505802 149940 505830 150198
rect 506446 149940 506474 150198
rect 507090 150198 507164 150226
rect 507688 150226 507716 151914
rect 508424 150226 508452 158850
rect 509252 151978 509280 163200
rect 510080 158914 510108 163200
rect 510068 158908 510120 158914
rect 510068 158850 510120 158856
rect 509700 158772 509752 158778
rect 509700 158714 509752 158720
rect 509240 151972 509292 151978
rect 509240 151914 509292 151920
rect 509056 151836 509108 151842
rect 509056 151778 509108 151784
rect 509068 150226 509096 151778
rect 509712 150226 509740 158714
rect 510344 152856 510396 152862
rect 510344 152798 510396 152804
rect 510356 150226 510384 152798
rect 510908 151842 510936 163200
rect 511736 158778 511764 163200
rect 511724 158772 511776 158778
rect 511724 158714 511776 158720
rect 511632 153196 511684 153202
rect 511632 153138 511684 153144
rect 510988 153128 511040 153134
rect 510988 153070 511040 153076
rect 510896 151836 510948 151842
rect 510896 151778 510948 151784
rect 511000 150226 511028 153070
rect 511644 150226 511672 153138
rect 512012 152862 512040 163254
rect 512564 163146 512592 163254
rect 512642 163200 512698 164400
rect 513470 163200 513526 164400
rect 513760 163254 514248 163282
rect 512656 163146 512684 163200
rect 512564 163118 512684 163146
rect 513484 153134 513512 163200
rect 513760 153202 513788 163254
rect 514220 163146 514248 163254
rect 514298 163200 514354 164400
rect 514864 163254 515076 163282
rect 514312 163146 514340 163200
rect 514220 163118 514340 163146
rect 513748 153196 513800 153202
rect 513748 153138 513800 153144
rect 514208 153196 514260 153202
rect 514208 153138 514260 153144
rect 513472 153128 513524 153134
rect 513472 153070 513524 153076
rect 513564 153128 513616 153134
rect 513564 153070 513616 153076
rect 512276 153060 512328 153066
rect 512276 153002 512328 153008
rect 512000 152856 512052 152862
rect 512000 152798 512052 152804
rect 512288 150226 512316 153002
rect 512920 152992 512972 152998
rect 512920 152934 512972 152940
rect 512932 150226 512960 152934
rect 513576 150226 513604 153070
rect 514220 150226 514248 153138
rect 514864 153066 514892 163254
rect 515048 163146 515076 163254
rect 515126 163200 515182 164400
rect 515954 163200 516010 164400
rect 516152 163254 516732 163282
rect 515140 163146 515168 163200
rect 515048 163118 515168 163146
rect 514944 158772 514996 158778
rect 514944 158714 514996 158720
rect 514852 153060 514904 153066
rect 514852 153002 514904 153008
rect 514956 151814 514984 158714
rect 515968 152998 515996 163200
rect 516152 153134 516180 163254
rect 516704 163146 516732 163254
rect 516782 163200 516838 164400
rect 517610 163200 517666 164400
rect 518530 163200 518586 164400
rect 519004 163254 519308 163282
rect 516796 163146 516824 163200
rect 516704 163118 516824 163146
rect 517624 161474 517652 163200
rect 517532 161446 517652 161474
rect 517532 158794 517560 161446
rect 518072 159520 518124 159526
rect 518072 159462 518124 159468
rect 517440 158766 517560 158794
rect 517440 153202 517468 158766
rect 517428 153196 517480 153202
rect 517428 153138 517480 153144
rect 516140 153128 516192 153134
rect 516140 153070 516192 153076
rect 515956 152992 516008 152998
rect 515956 152934 516008 152940
rect 516692 152176 516744 152182
rect 516692 152118 516744 152124
rect 515496 152108 515548 152114
rect 515496 152050 515548 152056
rect 514864 151786 514984 151814
rect 514864 150226 514892 151786
rect 515508 150226 515536 152050
rect 515956 152040 516008 152046
rect 515956 151982 516008 151988
rect 515968 151814 515996 151982
rect 515968 151786 516088 151814
rect 507688 150198 507762 150226
rect 507090 149940 507118 150198
rect 507734 149940 507762 150198
rect 508378 150198 508452 150226
rect 509022 150198 509096 150226
rect 509666 150198 509740 150226
rect 510310 150198 510384 150226
rect 510954 150198 511028 150226
rect 511598 150198 511672 150226
rect 512242 150198 512316 150226
rect 512886 150198 512960 150226
rect 513530 150198 513604 150226
rect 514174 150198 514248 150226
rect 514818 150198 514892 150226
rect 515462 150198 515536 150226
rect 516060 150226 516088 151786
rect 516704 150226 516732 152118
rect 517428 151972 517480 151978
rect 517428 151914 517480 151920
rect 517440 150226 517468 151914
rect 518084 150226 518112 159462
rect 518544 158778 518572 163200
rect 518716 159384 518768 159390
rect 518716 159326 518768 159332
rect 518532 158772 518584 158778
rect 518532 158714 518584 158720
rect 518728 150226 518756 159326
rect 519004 152114 519032 163254
rect 519280 163146 519308 163254
rect 519358 163200 519414 164400
rect 519924 163254 520136 163282
rect 519372 163146 519400 163200
rect 519280 163118 519400 163146
rect 519726 163160 519782 163169
rect 519726 163095 519782 163104
rect 519542 161664 519598 161673
rect 519542 161599 519598 161608
rect 518992 152108 519044 152114
rect 518992 152050 519044 152056
rect 519450 151056 519506 151065
rect 519450 150991 519506 151000
rect 516060 150198 516134 150226
rect 516704 150198 516778 150226
rect 508378 149940 508406 150198
rect 509022 149940 509050 150198
rect 509666 149940 509694 150198
rect 510310 149940 510338 150198
rect 510954 149940 510982 150198
rect 511598 149940 511626 150198
rect 512242 149940 512270 150198
rect 512886 149940 512914 150198
rect 513530 149940 513558 150198
rect 514174 149940 514202 150198
rect 514818 149940 514846 150198
rect 515462 149940 515490 150198
rect 516106 149940 516134 150198
rect 516750 149940 516778 150198
rect 517394 150198 517468 150226
rect 518038 150198 518112 150226
rect 518682 150198 518756 150226
rect 517394 149940 517422 150198
rect 518038 149940 518066 150198
rect 518682 149940 518710 150198
rect 519358 143440 519414 143449
rect 519358 143375 519414 143384
rect 519266 138952 519322 138961
rect 519266 138887 519322 138896
rect 519280 127401 519308 138887
rect 519372 131481 519400 143375
rect 519464 138417 519492 150991
rect 519556 147937 519584 161599
rect 519634 160168 519690 160177
rect 519634 160103 519690 160112
rect 519542 147928 519598 147937
rect 519542 147863 519598 147872
rect 519648 146577 519676 160103
rect 519740 149297 519768 163095
rect 519818 158672 519874 158681
rect 519818 158607 519874 158616
rect 519726 149288 519782 149297
rect 519726 149223 519782 149232
rect 519726 148064 519782 148073
rect 519726 147999 519782 148008
rect 519634 146568 519690 146577
rect 519634 146503 519690 146512
rect 519542 144936 519598 144945
rect 519542 144871 519598 144880
rect 519450 138408 519506 138417
rect 519450 138343 519506 138352
rect 519556 132977 519584 144871
rect 519740 135697 519768 147999
rect 519832 145217 519860 158607
rect 519924 152046 519952 163254
rect 520108 163146 520136 163254
rect 520186 163200 520242 164400
rect 520292 163254 520964 163282
rect 520200 163146 520228 163200
rect 520108 163118 520228 163146
rect 520186 157176 520242 157185
rect 520186 157111 520242 157120
rect 520094 155680 520150 155689
rect 520094 155615 520150 155624
rect 520002 154048 520058 154057
rect 520002 153983 520058 153992
rect 519912 152040 519964 152046
rect 519912 151982 519964 151988
rect 519910 149560 519966 149569
rect 519910 149495 519966 149504
rect 519818 145208 519874 145217
rect 519818 145143 519874 145152
rect 519924 137057 519952 149495
rect 520016 141137 520044 153983
rect 520108 142497 520136 155615
rect 520200 143857 520228 157111
rect 520292 152182 520320 163254
rect 520936 163146 520964 163254
rect 521014 163200 521070 164400
rect 521842 163200 521898 164400
rect 522670 163200 522726 164400
rect 523498 163200 523554 164400
rect 521028 163146 521056 163200
rect 520936 163118 521056 163146
rect 521856 161474 521884 163200
rect 521672 161446 521884 161474
rect 521672 158794 521700 161446
rect 522684 159526 522712 163200
rect 522672 159520 522724 159526
rect 522672 159462 522724 159468
rect 523512 159390 523540 163200
rect 523500 159384 523552 159390
rect 523500 159326 523552 159332
rect 521580 158766 521700 158794
rect 521014 152552 521070 152561
rect 521014 152487 521070 152496
rect 520280 152176 520332 152182
rect 520280 152118 520332 152124
rect 520922 146568 520978 146577
rect 520922 146503 520978 146512
rect 520186 143848 520242 143857
rect 520186 143783 520242 143792
rect 520094 142488 520150 142497
rect 520094 142423 520150 142432
rect 520186 141944 520242 141953
rect 520186 141879 520242 141888
rect 520002 141128 520058 141137
rect 520002 141063 520058 141072
rect 520002 140448 520058 140457
rect 520002 140383 520058 140392
rect 519910 137048 519966 137057
rect 519910 136983 519966 136992
rect 519910 135824 519966 135833
rect 519910 135759 519966 135768
rect 519726 135688 519782 135697
rect 519726 135623 519782 135632
rect 519634 134328 519690 134337
rect 519634 134263 519690 134272
rect 519542 132968 519598 132977
rect 519542 132903 519598 132912
rect 519358 131472 519414 131481
rect 519358 131407 519414 131416
rect 519542 129840 519598 129849
rect 519542 129775 519598 129784
rect 519266 127392 519322 127401
rect 519266 127327 519322 127336
rect 519450 126712 519506 126721
rect 519450 126647 519506 126656
rect 519358 125216 519414 125225
rect 519358 125151 519414 125160
rect 117228 118040 117280 118046
rect 117228 117982 117280 117988
rect 519372 115161 519400 125151
rect 519464 116521 519492 126647
rect 519556 119241 519584 129775
rect 519648 123321 519676 134263
rect 519726 132832 519782 132841
rect 519726 132767 519782 132776
rect 519634 123312 519690 123321
rect 519634 123247 519690 123256
rect 519740 121961 519768 132767
rect 519818 131336 519874 131345
rect 519818 131271 519874 131280
rect 519726 121952 519782 121961
rect 519726 121887 519782 121896
rect 519634 120728 519690 120737
rect 519634 120663 519690 120672
rect 519542 119232 519598 119241
rect 519542 119167 519598 119176
rect 519450 116512 519506 116521
rect 519450 116447 519506 116456
rect 519358 115152 519414 115161
rect 519358 115087 519414 115096
rect 519542 114608 519598 114617
rect 519542 114543 519598 114552
rect 519556 105505 519584 114543
rect 519648 110945 519676 120663
rect 519832 120601 519860 131271
rect 519924 124681 519952 135759
rect 520016 128761 520044 140383
rect 520094 137456 520150 137465
rect 520094 137391 520150 137400
rect 520002 128752 520058 128761
rect 520002 128687 520058 128696
rect 520002 128344 520058 128353
rect 520002 128279 520058 128288
rect 519910 124672 519966 124681
rect 519910 124607 519966 124616
rect 519818 120592 519874 120601
rect 519818 120527 519874 120536
rect 519726 119232 519782 119241
rect 519726 119167 519782 119176
rect 519634 110936 519690 110945
rect 519634 110871 519690 110880
rect 519740 109585 519768 119167
rect 520016 117881 520044 128279
rect 520108 126041 520136 137391
rect 520200 130121 520228 141879
rect 520936 134473 520964 146503
rect 521028 139777 521056 152487
rect 521580 151978 521608 158766
rect 521568 151972 521620 151978
rect 521568 151914 521620 151920
rect 521014 139768 521070 139777
rect 521014 139703 521070 139712
rect 520922 134464 520978 134473
rect 520922 134399 520978 134408
rect 520186 130112 520242 130121
rect 520186 130047 520242 130056
rect 520094 126032 520150 126041
rect 520094 125967 520150 125976
rect 520094 123720 520150 123729
rect 520094 123655 520150 123664
rect 520002 117872 520058 117881
rect 520002 117807 520058 117816
rect 519818 117600 519874 117609
rect 519818 117535 519874 117544
rect 519726 109576 519782 109585
rect 519726 109511 519782 109520
rect 519832 108225 519860 117535
rect 519910 116104 519966 116113
rect 519910 116039 519966 116048
rect 519818 108216 519874 108225
rect 519818 108151 519874 108160
rect 519924 106865 519952 116039
rect 520108 113801 520136 123655
rect 520186 122224 520242 122233
rect 520186 122159 520242 122168
rect 520094 113792 520150 113801
rect 520094 113727 520150 113736
rect 520200 112305 520228 122159
rect 521014 113112 521070 113121
rect 521014 113047 521070 113056
rect 520186 112296 520242 112305
rect 520186 112231 520242 112240
rect 520922 110120 520978 110129
rect 520922 110055 520978 110064
rect 519910 106856 519966 106865
rect 519910 106791 519966 106800
rect 519542 105496 519598 105505
rect 519542 105431 519598 105440
rect 520278 105496 520334 105505
rect 520278 105431 520334 105440
rect 117134 104816 117190 104825
rect 117134 104751 117190 104760
rect 117042 102912 117098 102921
rect 117042 102847 117098 102856
rect 116950 101008 117006 101017
rect 116950 100943 117006 100952
rect 519818 99376 519874 99385
rect 519818 99311 519874 99320
rect 116858 99104 116914 99113
rect 116858 99039 116914 99048
rect 519726 97880 519782 97889
rect 519726 97815 519782 97824
rect 116766 97200 116822 97209
rect 116766 97135 116822 97144
rect 116674 95296 116730 95305
rect 116674 95231 116730 95240
rect 519266 94888 519322 94897
rect 519266 94823 519322 94832
rect 116582 93392 116638 93401
rect 116582 93327 116638 93336
rect 116124 92472 116176 92478
rect 116124 92414 116176 92420
rect 116136 91361 116164 92414
rect 116122 91352 116178 91361
rect 116122 91287 116178 91296
rect 116124 89684 116176 89690
rect 116124 89626 116176 89632
rect 116136 89457 116164 89626
rect 116122 89448 116178 89457
rect 116122 89383 116178 89392
rect 116032 88324 116084 88330
rect 116032 88266 116084 88272
rect 116044 87553 116072 88266
rect 519280 87689 519308 94823
rect 519450 91896 519506 91905
rect 519450 91831 519506 91840
rect 519266 87680 519322 87689
rect 519266 87615 519322 87624
rect 116030 87544 116086 87553
rect 116030 87479 116086 87488
rect 114466 87272 114522 87281
rect 114466 87207 114468 87216
rect 114520 87207 114522 87216
rect 116492 87236 116544 87242
rect 114468 87178 114520 87184
rect 116492 87178 116544 87184
rect 116216 86964 116268 86970
rect 116216 86906 116268 86912
rect 116228 85649 116256 86906
rect 116214 85640 116270 85649
rect 116214 85575 116270 85584
rect 116308 82816 116360 82822
rect 116308 82758 116360 82764
rect 116320 81841 116348 82758
rect 116306 81832 116362 81841
rect 116306 81767 116362 81776
rect 114192 80028 114244 80034
rect 114192 79970 114244 79976
rect 115940 80028 115992 80034
rect 115940 79970 115992 79976
rect 115952 79937 115980 79970
rect 115938 79928 115994 79937
rect 115938 79863 115994 79872
rect 116504 78033 116532 87178
rect 519464 84969 519492 91831
rect 519740 90409 519768 97815
rect 519832 91769 519860 99311
rect 520292 97345 520320 105431
rect 520738 102504 520794 102513
rect 520738 102439 520794 102448
rect 520278 97336 520334 97345
rect 520278 97271 520334 97280
rect 520094 96384 520150 96393
rect 520094 96319 520150 96328
rect 520002 93392 520058 93401
rect 520002 93327 520058 93336
rect 519818 91760 519874 91769
rect 519818 91695 519874 91704
rect 519726 90400 519782 90409
rect 519726 90335 519782 90344
rect 519910 90264 519966 90273
rect 519910 90199 519966 90208
rect 519726 87272 519782 87281
rect 519726 87207 519782 87216
rect 519450 84960 519506 84969
rect 519450 84895 519506 84904
rect 519266 84280 519322 84289
rect 519266 84215 519322 84224
rect 116584 83972 116636 83978
rect 116584 83914 116636 83920
rect 116596 83745 116624 83914
rect 116582 83736 116638 83745
rect 116582 83671 116638 83680
rect 519280 78169 519308 84215
rect 519450 81152 519506 81161
rect 519450 81087 519506 81096
rect 519266 78160 519322 78169
rect 519266 78095 519322 78104
rect 116490 78024 116546 78033
rect 116490 77959 116546 77968
rect 519464 75313 519492 81087
rect 519740 80889 519768 87207
rect 519818 85776 519874 85785
rect 519818 85711 519874 85720
rect 519726 80880 519782 80889
rect 519726 80815 519782 80824
rect 519634 79656 519690 79665
rect 519634 79591 519690 79600
rect 519450 75304 519506 75313
rect 519450 75239 519506 75248
rect 116674 74080 116730 74089
rect 116674 74015 116730 74024
rect 116582 72176 116638 72185
rect 116582 72111 116638 72120
rect 116596 71806 116624 72111
rect 114192 71800 114244 71806
rect 114192 71742 114244 71748
rect 116584 71800 116636 71806
rect 116584 71742 116636 71748
rect 114100 69080 114152 69086
rect 114100 69022 114152 69028
rect 114008 67652 114060 67658
rect 114008 67594 114060 67600
rect 113916 66292 113968 66298
rect 113916 66234 113968 66240
rect 113824 63572 113876 63578
rect 113824 63514 113876 63520
rect 109684 41472 109736 41478
rect 109684 41414 109736 41420
rect 109592 3052 109644 3058
rect 109592 2994 109644 3000
rect 2504 2916 2556 2922
rect 2504 2858 2556 2864
rect 2516 2666 2544 2858
rect 109604 2689 109632 2994
rect 39118 2680 39174 2689
rect 2516 2638 2714 2666
rect 32772 2644 32824 2650
rect 53470 2680 53526 2689
rect 39330 2650 39712 2666
rect 39330 2644 39724 2650
rect 39330 2638 39672 2644
rect 39118 2615 39120 2624
rect 32772 2586 32824 2592
rect 39172 2615 39174 2624
rect 39120 2586 39172 2592
rect 39672 2586 39724 2592
rect 40316 2644 40368 2650
rect 42642 2638 42840 2666
rect 49358 2650 49648 2666
rect 40316 2586 40368 2592
rect 6012 1426 6040 2108
rect 9324 1465 9352 2108
rect 12636 1601 12664 2108
rect 15948 1737 15976 2108
rect 19352 1873 19380 2108
rect 19338 1864 19394 1873
rect 19338 1799 19394 1808
rect 15934 1728 15990 1737
rect 15934 1663 15990 1672
rect 12622 1592 12678 1601
rect 12622 1527 12678 1536
rect 22664 1494 22692 2108
rect 25976 1562 26004 2108
rect 29288 1630 29316 2108
rect 32692 1698 32720 2108
rect 32680 1692 32732 1698
rect 32680 1634 32732 1640
rect 29276 1624 29328 1630
rect 29276 1566 29328 1572
rect 25964 1556 26016 1562
rect 25964 1498 26016 1504
rect 22652 1488 22704 1494
rect 9310 1456 9366 1465
rect 6000 1420 6052 1426
rect 22652 1430 22704 1436
rect 9310 1391 9366 1400
rect 6000 1362 6052 1368
rect 32784 800 32812 2586
rect 36018 2514 36400 2530
rect 40328 2514 40356 2586
rect 42812 2553 42840 2638
rect 47492 2644 47544 2650
rect 47492 2586 47544 2592
rect 49148 2644 49200 2650
rect 49358 2644 49660 2650
rect 49358 2638 49608 2644
rect 49148 2586 49200 2592
rect 49608 2586 49660 2592
rect 50896 2644 50948 2650
rect 50896 2586 50948 2592
rect 53012 2644 53064 2650
rect 81254 2680 81310 2689
rect 62698 2650 62804 2666
rect 53470 2615 53472 2624
rect 53012 2586 53064 2592
rect 53524 2615 53526 2624
rect 53656 2644 53708 2650
rect 53472 2586 53524 2592
rect 53656 2586 53708 2592
rect 57520 2644 57572 2650
rect 57520 2586 57572 2592
rect 58624 2644 58676 2650
rect 58624 2586 58676 2592
rect 58716 2644 58768 2650
rect 58716 2586 58768 2592
rect 62396 2644 62448 2650
rect 62698 2644 62816 2650
rect 62698 2638 62764 2644
rect 62396 2586 62448 2592
rect 62764 2586 62816 2592
rect 63040 2644 63092 2650
rect 63040 2586 63092 2592
rect 63132 2644 63184 2650
rect 63132 2586 63184 2592
rect 65524 2644 65576 2650
rect 65524 2586 65576 2592
rect 78036 2644 78088 2650
rect 78036 2586 78088 2592
rect 78128 2644 78180 2650
rect 78128 2586 78180 2592
rect 78496 2644 78548 2650
rect 78496 2586 78548 2592
rect 79692 2644 79744 2650
rect 79692 2586 79744 2592
rect 79784 2644 79836 2650
rect 79784 2586 79836 2592
rect 81164 2644 81216 2650
rect 106094 2680 106150 2689
rect 81254 2615 81256 2624
rect 81164 2586 81216 2592
rect 81308 2615 81310 2624
rect 81348 2644 81400 2650
rect 81256 2586 81308 2592
rect 81348 2586 81400 2592
rect 82084 2644 82136 2650
rect 82084 2586 82136 2592
rect 82176 2644 82228 2650
rect 82176 2586 82228 2592
rect 82268 2644 82320 2650
rect 82268 2586 82320 2592
rect 98276 2644 98328 2650
rect 106094 2615 106096 2624
rect 98276 2586 98328 2592
rect 106148 2615 106150 2624
rect 109590 2680 109646 2689
rect 109590 2615 109646 2624
rect 106096 2586 106148 2592
rect 46296 2576 46348 2582
rect 42798 2544 42854 2553
rect 36018 2508 36412 2514
rect 36018 2502 36360 2508
rect 36360 2450 36412 2456
rect 40316 2508 40368 2514
rect 46046 2524 46296 2530
rect 46046 2518 46348 2524
rect 46046 2502 46336 2518
rect 42798 2479 42854 2488
rect 40316 2450 40368 2456
rect 47504 2242 47532 2586
rect 49160 2417 49188 2586
rect 50908 2553 50936 2586
rect 50894 2544 50950 2553
rect 50894 2479 50950 2488
rect 52920 2440 52972 2446
rect 49146 2408 49202 2417
rect 52670 2388 52920 2394
rect 52670 2382 52972 2388
rect 52670 2366 52960 2382
rect 49146 2343 49202 2352
rect 53024 2310 53052 2586
rect 53668 2446 53696 2586
rect 56232 2576 56284 2582
rect 55982 2524 56232 2530
rect 55982 2518 56284 2524
rect 55982 2502 56272 2518
rect 53656 2440 53708 2446
rect 53656 2382 53708 2388
rect 53012 2304 53064 2310
rect 53012 2246 53064 2252
rect 47492 2236 47544 2242
rect 47492 2178 47544 2184
rect 57532 2174 57560 2586
rect 58636 2553 58664 2586
rect 58622 2544 58678 2553
rect 58622 2479 58678 2488
rect 58728 2242 58756 2586
rect 59728 2440 59780 2446
rect 59386 2388 59728 2394
rect 62408 2417 62436 2586
rect 63052 2417 63080 2586
rect 59386 2382 59780 2388
rect 62394 2408 62450 2417
rect 59386 2366 59768 2382
rect 62394 2343 62450 2352
rect 63038 2408 63094 2417
rect 63038 2343 63094 2352
rect 63144 2242 63172 2586
rect 65536 2446 65564 2586
rect 73988 2576 74040 2582
rect 74080 2576 74132 2582
rect 74040 2536 74080 2564
rect 73988 2518 74040 2524
rect 74080 2518 74132 2524
rect 76656 2576 76708 2582
rect 76656 2518 76708 2524
rect 65524 2440 65576 2446
rect 66352 2440 66404 2446
rect 65524 2382 65576 2388
rect 66010 2388 66352 2394
rect 66010 2382 66404 2388
rect 66010 2366 66392 2382
rect 76668 2310 76696 2518
rect 78048 2417 78076 2586
rect 78034 2408 78090 2417
rect 78034 2343 78090 2352
rect 76564 2304 76616 2310
rect 69322 2242 69704 2258
rect 76564 2246 76616 2252
rect 76656 2304 76708 2310
rect 78140 2281 78168 2586
rect 76656 2246 76708 2252
rect 78126 2272 78182 2281
rect 58716 2236 58768 2242
rect 58716 2178 58768 2184
rect 63132 2236 63184 2242
rect 69322 2236 69716 2242
rect 69322 2230 69664 2236
rect 63132 2178 63184 2184
rect 69664 2178 69716 2184
rect 76576 2174 76604 2246
rect 78126 2207 78182 2216
rect 57520 2168 57572 2174
rect 57520 2110 57572 2116
rect 76564 2168 76616 2174
rect 76564 2110 76616 2116
rect 72712 1834 72740 2108
rect 72700 1828 72752 1834
rect 72700 1770 72752 1776
rect 76024 1766 76052 2108
rect 78508 2106 78536 2586
rect 79416 2576 79468 2582
rect 79600 2576 79652 2582
rect 79468 2536 79600 2564
rect 79416 2518 79468 2524
rect 79600 2518 79652 2524
rect 79704 2281 79732 2586
rect 79796 2417 79824 2586
rect 79782 2408 79838 2417
rect 81176 2378 81204 2586
rect 79782 2343 79838 2352
rect 81164 2372 81216 2378
rect 81164 2314 81216 2320
rect 79690 2272 79746 2281
rect 79690 2207 79746 2216
rect 81360 2174 81388 2586
rect 82096 2446 82124 2586
rect 82084 2440 82136 2446
rect 82084 2382 82136 2388
rect 82188 2242 82216 2586
rect 82280 2553 82308 2586
rect 82266 2544 82322 2553
rect 82266 2479 82322 2488
rect 96002 2242 96384 2258
rect 82176 2236 82228 2242
rect 96002 2236 96396 2242
rect 96002 2230 96344 2236
rect 82176 2178 82228 2184
rect 96344 2178 96396 2184
rect 81348 2168 81400 2174
rect 93032 2168 93084 2174
rect 81348 2110 81400 2116
rect 78496 2100 78548 2106
rect 78496 2042 78548 2048
rect 79336 1902 79364 2108
rect 82648 1970 82676 2108
rect 86066 2094 86448 2122
rect 89378 2106 89668 2122
rect 92690 2116 93032 2122
rect 92690 2110 93084 2116
rect 89378 2100 89680 2106
rect 89378 2094 89628 2100
rect 86420 2038 86448 2094
rect 92690 2094 93072 2110
rect 89628 2042 89680 2048
rect 86408 2032 86460 2038
rect 86408 1974 86460 1980
rect 82636 1964 82688 1970
rect 82636 1906 82688 1912
rect 79324 1896 79376 1902
rect 79324 1838 79376 1844
rect 76012 1760 76064 1766
rect 76012 1702 76064 1708
rect 98288 800 98316 2586
rect 109342 2514 109632 2530
rect 109342 2508 109644 2514
rect 109342 2502 109592 2508
rect 109592 2450 109644 2456
rect 106188 2440 106240 2446
rect 102718 2378 103008 2394
rect 106030 2388 106188 2394
rect 106030 2382 106240 2388
rect 102718 2372 103020 2378
rect 102718 2366 102968 2372
rect 106030 2366 106228 2382
rect 102968 2314 103020 2320
rect 99656 2304 99708 2310
rect 99406 2252 99656 2258
rect 99406 2246 99708 2252
rect 99406 2230 99696 2246
rect 109696 1834 109724 41414
rect 111064 34536 111116 34542
rect 111064 34478 111116 34484
rect 109776 4208 109828 4214
rect 109776 4150 109828 4156
rect 109684 1828 109736 1834
rect 109684 1770 109736 1776
rect 109788 1426 109816 4150
rect 111076 3942 111104 34478
rect 112444 33176 112496 33182
rect 112444 33118 112496 33124
rect 111156 23520 111208 23526
rect 111156 23462 111208 23468
rect 111064 3936 111116 3942
rect 111064 3878 111116 3884
rect 111168 3534 111196 23462
rect 111248 22160 111300 22166
rect 111248 22102 111300 22108
rect 111156 3528 111208 3534
rect 111156 3470 111208 3476
rect 111260 3466 111288 22102
rect 112456 3874 112484 33118
rect 112536 31816 112588 31822
rect 112536 31758 112588 31764
rect 112444 3868 112496 3874
rect 112444 3810 112496 3816
rect 112548 3806 112576 31758
rect 112628 29028 112680 29034
rect 112628 28970 112680 28976
rect 112536 3800 112588 3806
rect 112536 3742 112588 3748
rect 112640 3738 112668 28970
rect 112720 27668 112772 27674
rect 112720 27610 112772 27616
rect 112628 3732 112680 3738
rect 112628 3674 112680 3680
rect 112732 3670 112760 27610
rect 112812 24880 112864 24886
rect 112812 24822 112864 24828
rect 112720 3664 112772 3670
rect 112720 3606 112772 3612
rect 112824 3602 112852 24822
rect 113836 7721 113864 63514
rect 113928 19009 113956 66234
rect 114020 30433 114048 67594
rect 114112 41857 114140 69022
rect 114204 53145 114232 71742
rect 116306 70272 116362 70281
rect 116306 70207 116362 70216
rect 116320 69086 116348 70207
rect 116308 69080 116360 69086
rect 116308 69022 116360 69028
rect 116122 68368 116178 68377
rect 116122 68303 116178 68312
rect 116136 67658 116164 68303
rect 116124 67652 116176 67658
rect 116124 67594 116176 67600
rect 116582 66464 116638 66473
rect 116582 66399 116638 66408
rect 116596 66298 116624 66399
rect 116584 66292 116636 66298
rect 116584 66234 116636 66240
rect 116688 64874 116716 74015
rect 519648 73953 519676 79591
rect 519832 79529 519860 85711
rect 519924 83609 519952 90199
rect 520016 86329 520044 93327
rect 520108 89049 520136 96319
rect 520752 94489 520780 102439
rect 520936 101425 520964 110055
rect 521028 104145 521056 113047
rect 521106 111616 521162 111625
rect 521106 111551 521162 111560
rect 521014 104136 521070 104145
rect 521014 104071 521070 104080
rect 521120 102785 521148 111551
rect 521198 108488 521254 108497
rect 521198 108423 521254 108432
rect 521106 102776 521162 102785
rect 521106 102711 521162 102720
rect 520922 101416 520978 101425
rect 520922 101351 520978 101360
rect 521106 101008 521162 101017
rect 521106 100943 521162 100952
rect 520738 94480 520794 94489
rect 520738 94415 520794 94424
rect 521120 93129 521148 100943
rect 521212 100065 521240 108423
rect 521474 106992 521530 107001
rect 521474 106927 521530 106936
rect 521290 104000 521346 104009
rect 521290 103935 521346 103944
rect 521198 100056 521254 100065
rect 521198 99991 521254 100000
rect 521304 95985 521332 103935
rect 521488 98705 521516 106927
rect 521474 98696 521530 98705
rect 521474 98631 521530 98640
rect 521290 95976 521346 95985
rect 521290 95911 521346 95920
rect 521106 93120 521162 93129
rect 521106 93055 521162 93064
rect 520094 89040 520150 89049
rect 520094 88975 520150 88984
rect 520186 88768 520242 88777
rect 520186 88703 520242 88712
rect 520002 86320 520058 86329
rect 520002 86255 520058 86264
rect 519910 83600 519966 83609
rect 519910 83535 519966 83544
rect 520094 82784 520150 82793
rect 520094 82719 520150 82728
rect 519818 79520 519874 79529
rect 519818 79455 519874 79464
rect 519726 78160 519782 78169
rect 519726 78095 519782 78104
rect 519634 73944 519690 73953
rect 519634 73879 519690 73888
rect 519740 72593 519768 78095
rect 520108 76809 520136 82719
rect 520200 82249 520228 88703
rect 520186 82240 520242 82249
rect 520186 82175 520242 82184
rect 520094 76800 520150 76809
rect 520094 76735 520150 76744
rect 520002 76664 520058 76673
rect 520002 76599 520058 76608
rect 519818 75168 519874 75177
rect 519818 75103 519874 75112
rect 519726 72584 519782 72593
rect 519726 72519 519782 72528
rect 519832 69873 519860 75103
rect 519910 73672 519966 73681
rect 519910 73607 519966 73616
rect 519818 69864 519874 69873
rect 519818 69799 519874 69808
rect 519634 69048 519690 69057
rect 519634 68983 519690 68992
rect 116596 64846 116716 64874
rect 116596 64598 116624 64846
rect 114468 64592 114520 64598
rect 114466 64560 114468 64569
rect 116584 64592 116636 64598
rect 114520 64560 114522 64569
rect 114466 64495 114522 64504
rect 116214 64560 116270 64569
rect 116584 64534 116636 64540
rect 116214 64495 116270 64504
rect 116228 63578 116256 64495
rect 519648 64433 519676 68983
rect 519924 68513 519952 73607
rect 520016 71233 520044 76599
rect 520094 72040 520150 72049
rect 520094 71975 520150 71984
rect 520002 71224 520058 71233
rect 520002 71159 520058 71168
rect 519910 68504 519966 68513
rect 519910 68439 519966 68448
rect 520108 67153 520136 71975
rect 520186 70544 520242 70553
rect 520186 70479 520242 70488
rect 520094 67144 520150 67153
rect 520094 67079 520150 67088
rect 520200 65793 520228 70479
rect 520462 67552 520518 67561
rect 520462 67487 520518 67496
rect 520370 66056 520426 66065
rect 520370 65991 520426 66000
rect 520186 65784 520242 65793
rect 520186 65719 520242 65728
rect 519634 64424 519690 64433
rect 519634 64359 519690 64368
rect 116216 63572 116268 63578
rect 116216 63514 116268 63520
rect 116582 62656 116638 62665
rect 116582 62591 116638 62600
rect 114190 53136 114246 53145
rect 114190 53071 114246 53080
rect 116490 47152 116546 47161
rect 116490 47087 116546 47096
rect 116214 45248 116270 45257
rect 116214 45183 116270 45192
rect 114098 41848 114154 41857
rect 114098 41783 114154 41792
rect 116124 41472 116176 41478
rect 116122 41440 116124 41449
rect 116176 41440 116178 41449
rect 116122 41375 116178 41384
rect 114100 38684 114152 38690
rect 114100 38626 114152 38632
rect 114006 30424 114062 30433
rect 114006 30359 114062 30368
rect 113914 19000 113970 19009
rect 113914 18935 113970 18944
rect 113822 7712 113878 7721
rect 113822 7647 113878 7656
rect 112812 3596 112864 3602
rect 112812 3538 112864 3544
rect 111248 3460 111300 3466
rect 111248 3402 111300 3408
rect 114112 3330 114140 38626
rect 116228 38554 116256 45183
rect 116306 43344 116362 43353
rect 116306 43279 116362 43288
rect 116216 38548 116268 38554
rect 116216 38490 116268 38496
rect 116214 37632 116270 37641
rect 116214 37567 116270 37576
rect 116228 37330 116256 37567
rect 114192 37324 114244 37330
rect 114192 37266 114244 37272
rect 116216 37324 116268 37330
rect 116216 37266 116268 37272
rect 114204 3398 114232 37266
rect 116122 35728 116178 35737
rect 116122 35663 116178 35672
rect 116136 34542 116164 35663
rect 116124 34536 116176 34542
rect 116124 34478 116176 34484
rect 116122 33824 116178 33833
rect 116122 33759 116178 33768
rect 116136 33182 116164 33759
rect 116124 33176 116176 33182
rect 116124 33118 116176 33124
rect 116124 31816 116176 31822
rect 116122 31784 116124 31793
rect 116176 31784 116178 31793
rect 116122 31719 116178 31728
rect 116122 29880 116178 29889
rect 116122 29815 116178 29824
rect 116136 29034 116164 29815
rect 116124 29028 116176 29034
rect 116124 28970 116176 28976
rect 116122 27976 116178 27985
rect 116122 27911 116178 27920
rect 116136 27674 116164 27911
rect 116124 27668 116176 27674
rect 116124 27610 116176 27616
rect 116122 26072 116178 26081
rect 116122 26007 116178 26016
rect 116136 24886 116164 26007
rect 116124 24880 116176 24886
rect 116124 24822 116176 24828
rect 116122 24168 116178 24177
rect 116122 24103 116178 24112
rect 116136 23526 116164 24103
rect 116124 23520 116176 23526
rect 116124 23462 116176 23468
rect 116030 22264 116086 22273
rect 116030 22199 116086 22208
rect 116044 22166 116072 22199
rect 116032 22160 116084 22166
rect 116032 22102 116084 22108
rect 116214 20360 116270 20369
rect 116214 20295 116270 20304
rect 116122 18456 116178 18465
rect 116122 18391 116178 18400
rect 116032 16516 116084 16522
rect 116032 16458 116084 16464
rect 115938 14512 115994 14521
rect 115938 14447 115994 14456
rect 115952 5234 115980 14447
rect 115940 5228 115992 5234
rect 115940 5170 115992 5176
rect 115940 5092 115992 5098
rect 115940 5034 115992 5040
rect 114192 3392 114244 3398
rect 114192 3334 114244 3340
rect 114100 3324 114152 3330
rect 114100 3266 114152 3272
rect 115952 1630 115980 5034
rect 116044 1698 116072 16458
rect 116136 5098 116164 18391
rect 116228 16522 116256 20295
rect 116216 16516 116268 16522
rect 116216 16458 116268 16464
rect 116214 16416 116270 16425
rect 116214 16351 116270 16360
rect 116228 11898 116256 16351
rect 116216 11892 116268 11898
rect 116216 11834 116268 11840
rect 116320 11778 116348 43279
rect 116398 39536 116454 39545
rect 116398 39471 116454 39480
rect 116412 38690 116440 39471
rect 116400 38684 116452 38690
rect 116400 38626 116452 38632
rect 116400 38548 116452 38554
rect 116400 38490 116452 38496
rect 116228 11750 116348 11778
rect 116124 5092 116176 5098
rect 116124 5034 116176 5040
rect 116122 4992 116178 5001
rect 116122 4927 116178 4936
rect 116136 4214 116164 4927
rect 116124 4208 116176 4214
rect 116124 4150 116176 4156
rect 116122 3088 116178 3097
rect 116122 3023 116178 3032
rect 116136 2922 116164 3023
rect 116124 2916 116176 2922
rect 116124 2858 116176 2864
rect 116228 1766 116256 11750
rect 116308 11688 116360 11694
rect 116308 11630 116360 11636
rect 116320 5370 116348 11630
rect 116308 5364 116360 5370
rect 116308 5306 116360 5312
rect 116308 5228 116360 5234
rect 116308 5170 116360 5176
rect 116216 1760 116268 1766
rect 116216 1702 116268 1708
rect 116032 1692 116084 1698
rect 116032 1634 116084 1640
rect 115940 1624 115992 1630
rect 115940 1566 115992 1572
rect 116320 1494 116348 5170
rect 116412 1902 116440 38490
rect 116504 1970 116532 47087
rect 116596 2514 116624 62591
rect 520384 61713 520412 65991
rect 520476 63073 520504 67487
rect 520738 64560 520794 64569
rect 520738 64495 520794 64504
rect 520462 63064 520518 63073
rect 520462 62999 520518 63008
rect 520370 61704 520426 61713
rect 520370 61639 520426 61648
rect 116674 60616 116730 60625
rect 116674 60551 116730 60560
rect 116584 2508 116636 2514
rect 116584 2450 116636 2456
rect 116688 2446 116716 60551
rect 520752 60353 520780 64495
rect 521106 62928 521162 62937
rect 521106 62863 521162 62872
rect 521014 61432 521070 61441
rect 521014 61367 521070 61376
rect 520738 60344 520794 60353
rect 520738 60279 520794 60288
rect 520738 59936 520794 59945
rect 520738 59871 520794 59880
rect 116766 58712 116822 58721
rect 116766 58647 116822 58656
rect 116676 2440 116728 2446
rect 116676 2382 116728 2388
rect 116780 2378 116808 58647
rect 520370 56944 520426 56953
rect 520370 56879 520426 56888
rect 116858 56808 116914 56817
rect 116858 56743 116914 56752
rect 116768 2372 116820 2378
rect 116768 2314 116820 2320
rect 116872 2310 116900 56743
rect 520278 55448 520334 55457
rect 520278 55383 520334 55392
rect 116950 54904 117006 54913
rect 116950 54839 117006 54848
rect 116964 11506 116992 54839
rect 519082 53816 519138 53825
rect 519082 53751 519138 53760
rect 117042 53000 117098 53009
rect 117042 52935 117098 52944
rect 117056 11642 117084 52935
rect 117134 51096 117190 51105
rect 117134 51031 117190 51040
rect 117148 11778 117176 51031
rect 519096 50697 519124 53751
rect 519910 52320 519966 52329
rect 519910 52255 519966 52264
rect 519082 50688 519138 50697
rect 519082 50623 519138 50632
rect 519924 49337 519952 52255
rect 520292 52057 520320 55383
rect 520384 53417 520412 56879
rect 520752 56137 520780 59871
rect 521028 57497 521056 61367
rect 521120 58993 521148 62863
rect 521106 58984 521162 58993
rect 521106 58919 521162 58928
rect 521106 58440 521162 58449
rect 521106 58375 521162 58384
rect 521014 57488 521070 57497
rect 521014 57423 521070 57432
rect 520738 56128 520794 56137
rect 520738 56063 520794 56072
rect 521120 54777 521148 58375
rect 521106 54768 521162 54777
rect 521106 54703 521162 54712
rect 520370 53408 520426 53417
rect 520370 53343 520426 53352
rect 520278 52048 520334 52057
rect 520278 51983 520334 51992
rect 520002 50824 520058 50833
rect 520002 50759 520058 50768
rect 519910 49328 519966 49337
rect 519910 49263 519966 49272
rect 117226 49192 117282 49201
rect 117226 49127 117282 49136
rect 117240 11914 117268 49127
rect 520016 47977 520044 50759
rect 520186 49328 520242 49337
rect 520186 49263 520242 49272
rect 520002 47968 520058 47977
rect 520002 47903 520058 47912
rect 519266 47832 519322 47841
rect 519266 47767 519322 47776
rect 519280 45257 519308 47767
rect 520200 46617 520228 49263
rect 520186 46608 520242 46617
rect 520186 46543 520242 46552
rect 519910 46336 519966 46345
rect 519910 46271 519966 46280
rect 519266 45248 519322 45257
rect 519266 45183 519322 45192
rect 519818 44704 519874 44713
rect 519818 44639 519874 44648
rect 519832 42537 519860 44639
rect 519924 43897 519952 46271
rect 519910 43888 519966 43897
rect 519910 43823 519966 43832
rect 520094 43208 520150 43217
rect 520094 43143 520150 43152
rect 519818 42528 519874 42537
rect 519818 42463 519874 42472
rect 520108 41177 520136 43143
rect 520186 41712 520242 41721
rect 520186 41647 520242 41656
rect 520094 41168 520150 41177
rect 520094 41103 520150 41112
rect 519818 40216 519874 40225
rect 519818 40151 519874 40160
rect 519832 38321 519860 40151
rect 520200 39817 520228 41647
rect 520186 39808 520242 39817
rect 520186 39743 520242 39752
rect 520186 38720 520242 38729
rect 520186 38655 520242 38664
rect 519818 38312 519874 38321
rect 519818 38247 519874 38256
rect 520200 36961 520228 38655
rect 521106 37224 521162 37233
rect 521106 37159 521162 37168
rect 520186 36952 520242 36961
rect 520186 36887 520242 36896
rect 521120 36009 521148 37159
rect 521106 36000 521162 36009
rect 521106 35935 521162 35944
rect 520922 35592 520978 35601
rect 520922 35527 520978 35536
rect 520936 34649 520964 35527
rect 520922 34640 520978 34649
rect 520922 34575 520978 34584
rect 520830 34096 520886 34105
rect 520830 34031 520886 34040
rect 520844 33289 520872 34031
rect 520830 33280 520886 33289
rect 520830 33215 520886 33224
rect 521106 32600 521162 32609
rect 521106 32535 521162 32544
rect 521120 31793 521148 32535
rect 521106 31784 521162 31793
rect 521106 31719 521162 31728
rect 521106 31104 521162 31113
rect 521106 31039 521162 31048
rect 521120 30433 521148 31039
rect 521106 30424 521162 30433
rect 521106 30359 521162 30368
rect 521106 29608 521162 29617
rect 521106 29543 521162 29552
rect 521120 28801 521148 29543
rect 521106 28792 521162 28801
rect 521106 28727 521162 28736
rect 521106 20496 521162 20505
rect 521106 20431 521162 20440
rect 521120 19825 521148 20431
rect 521106 19816 521162 19825
rect 521106 19751 521162 19760
rect 521106 15056 521162 15065
rect 521106 14991 521162 15000
rect 521120 14385 521148 14991
rect 521106 14376 521162 14385
rect 521106 14311 521162 14320
rect 521106 13696 521162 13705
rect 521106 13631 521162 13640
rect 521120 12889 521148 13631
rect 521106 12880 521162 12889
rect 521106 12815 521162 12824
rect 519634 12336 519690 12345
rect 519634 12271 519690 12280
rect 117240 11886 117360 11914
rect 117148 11750 117268 11778
rect 117056 11614 117176 11642
rect 116964 11478 117084 11506
rect 116952 11416 117004 11422
rect 116952 11358 117004 11364
rect 116964 5506 116992 11358
rect 116952 5500 117004 5506
rect 116952 5442 117004 5448
rect 116952 5364 117004 5370
rect 116952 5306 117004 5312
rect 116860 2304 116912 2310
rect 116860 2246 116912 2252
rect 116492 1964 116544 1970
rect 116492 1906 116544 1912
rect 116400 1896 116452 1902
rect 116400 1838 116452 1844
rect 116964 1562 116992 5306
rect 117056 2242 117084 11478
rect 117148 5658 117176 11614
rect 117240 5794 117268 11750
rect 117332 11422 117360 11886
rect 117320 11416 117372 11422
rect 519648 11393 519676 12271
rect 117320 11358 117372 11364
rect 519634 11384 519690 11393
rect 519634 11319 519690 11328
rect 521106 10976 521162 10985
rect 521106 10911 521162 10920
rect 521120 9897 521148 10911
rect 521106 9888 521162 9897
rect 521106 9823 521162 9832
rect 521106 9616 521162 9625
rect 521106 9551 521162 9560
rect 521120 8265 521148 9551
rect 520370 8256 520426 8265
rect 520370 8191 520426 8200
rect 521106 8256 521162 8265
rect 521106 8191 521162 8200
rect 520384 6769 520412 8191
rect 521106 6896 521162 6905
rect 521106 6831 521162 6840
rect 520370 6760 520426 6769
rect 520370 6695 520426 6704
rect 117240 5766 117360 5794
rect 117148 5630 117268 5658
rect 117136 5500 117188 5506
rect 117136 5442 117188 5448
rect 117044 2236 117096 2242
rect 117044 2178 117096 2184
rect 117148 2038 117176 5442
rect 117240 2174 117268 5630
rect 117228 2168 117280 2174
rect 117228 2110 117280 2116
rect 117332 2106 117360 5766
rect 521014 5536 521070 5545
rect 521014 5471 521070 5480
rect 521028 3777 521056 5471
rect 521120 5273 521148 6831
rect 521106 5264 521162 5273
rect 521106 5199 521162 5208
rect 521106 4176 521162 4185
rect 521106 4111 521162 4120
rect 521014 3768 521070 3777
rect 521014 3703 521070 3712
rect 117964 3052 118016 3058
rect 117964 2994 118016 3000
rect 117688 2984 117740 2990
rect 117688 2926 117740 2932
rect 117320 2100 117372 2106
rect 117320 2042 117372 2048
rect 117136 2032 117188 2038
rect 117136 1974 117188 1980
rect 116952 1556 117004 1562
rect 116952 1498 117004 1504
rect 117700 1494 117728 2926
rect 116308 1488 116360 1494
rect 116308 1430 116360 1436
rect 117688 1488 117740 1494
rect 117688 1430 117740 1436
rect 117976 1426 118004 2994
rect 520002 2816 520058 2825
rect 520002 2751 520058 2760
rect 443656 2650 443992 2666
rect 493612 2650 493948 2666
rect 294788 2644 294840 2650
rect 294788 2586 294840 2592
rect 425796 2644 425848 2650
rect 425796 2586 425848 2592
rect 443644 2644 443992 2650
rect 443696 2638 443992 2644
rect 491300 2644 491352 2650
rect 443644 2586 443696 2592
rect 491300 2586 491352 2592
rect 493600 2644 493948 2650
rect 493652 2638 493948 2644
rect 493600 2586 493652 2592
rect 143644 2094 143980 2122
rect 193600 2094 193936 2122
rect 243648 2094 243984 2122
rect 293604 2094 293940 2122
rect 143644 1494 143672 2094
rect 143632 1488 143684 1494
rect 143632 1430 143684 1436
rect 163778 1456 163834 1465
rect 109776 1420 109828 1426
rect 109776 1362 109828 1368
rect 117964 1420 118016 1426
rect 193600 1426 193628 2094
rect 229282 1592 229338 1601
rect 229282 1527 229338 1536
rect 163778 1391 163834 1400
rect 193588 1420 193640 1426
rect 117964 1362 118016 1368
rect 163792 800 163820 1391
rect 193588 1362 193640 1368
rect 229296 800 229324 1527
rect 243648 1465 243676 2094
rect 293604 1601 293632 2094
rect 293590 1592 293646 1601
rect 293590 1527 293646 1536
rect 243634 1456 243690 1465
rect 294800 1426 294828 2586
rect 343652 2094 343988 2122
rect 393608 2094 393944 2122
rect 343652 1426 343680 2094
rect 393608 1465 393636 2094
rect 360290 1456 360346 1465
rect 243634 1391 243690 1400
rect 294788 1420 294840 1426
rect 294788 1362 294840 1368
rect 343640 1420 343692 1426
rect 360290 1391 360346 1400
rect 393594 1456 393650 1465
rect 393594 1391 393650 1400
rect 343640 1362 343692 1368
rect 294800 800 294828 1362
rect 360304 800 360332 1391
rect 425808 800 425836 2586
rect 491312 800 491340 2586
rect 32770 -400 32826 800
rect 98274 -400 98330 800
rect 163778 -400 163834 800
rect 229282 -400 229338 800
rect 294786 -400 294842 800
rect 360290 -400 360346 800
rect 425794 -400 425850 800
rect 491298 -400 491354 800
rect 520016 785 520044 2751
rect 521120 2281 521148 4111
rect 521106 2272 521162 2281
rect 521106 2207 521162 2216
rect 520002 776 520058 785
rect 520002 711 520058 720
<< via2 >>
rect 16302 159432 16358 159488
rect 17130 153856 17186 153912
rect 20534 153720 20590 153776
rect 23018 159296 23074 159352
rect 28078 156712 28134 156768
rect 29826 159568 29882 159624
rect 31482 156576 31538 156632
rect 33966 157936 34022 157992
rect 40682 158208 40738 158264
rect 44086 158072 44142 158128
rect 42430 156848 42486 156904
rect 27250 153992 27306 154048
rect 49146 156984 49202 157040
rect 57518 158344 57574 158400
rect 55034 154264 55090 154320
rect 51630 154128 51686 154184
rect 12990 152496 13046 152552
rect 9586 152360 9642 152416
rect 61750 155216 61806 155272
rect 65982 157120 66038 157176
rect 76010 155624 76066 155680
rect 69294 155488 69350 155544
rect 68466 155352 68522 155408
rect 85302 155760 85358 155816
rect 89718 154400 89774 154456
rect 92018 155896 92074 155952
rect 104622 158480 104678 158536
rect 113086 157256 113142 157312
rect 116398 153584 116454 153640
rect 95790 149504 95846 149560
rect 102690 149504 102746 149560
rect 99286 149368 99342 149424
rect 102874 149368 102930 149424
rect 113822 144200 113878 144256
rect 115938 148996 115940 149016
rect 115940 148996 115992 149016
rect 115992 148996 115994 149016
rect 115938 148960 115994 148996
rect 116122 147056 116178 147112
rect 116030 145152 116086 145208
rect 116214 143248 116270 143304
rect 116490 141344 116546 141400
rect 115938 139440 115994 139496
rect 116398 137536 116454 137592
rect 115938 135496 115994 135552
rect 116122 133592 116178 133648
rect 113914 132776 113970 132832
rect 116122 131688 116178 131744
rect 116122 129784 116178 129840
rect 116122 127880 116178 127936
rect 116030 125976 116086 126032
rect 116122 124108 116124 124128
rect 116124 124108 116176 124128
rect 116176 124108 116178 124128
rect 116122 124072 116178 124108
rect 115938 122168 115994 122224
rect 114006 121352 114062 121408
rect 116122 120128 116178 120184
rect 116122 118224 116178 118280
rect 116122 116320 116178 116376
rect 116122 114452 116124 114472
rect 116124 114452 116176 114472
rect 116176 114452 116178 114472
rect 116122 114416 116178 114452
rect 115938 112512 115994 112568
rect 116122 110608 116178 110664
rect 114098 110064 114154 110120
rect 116122 108704 116178 108760
rect 116490 106800 116546 106856
rect 114190 98640 114246 98696
rect 120538 158908 120594 158944
rect 120538 158888 120540 158908
rect 120540 158888 120592 158908
rect 120592 158888 120594 158908
rect 119434 153584 119490 153640
rect 121550 158888 121606 158944
rect 122654 159160 122710 159216
rect 122838 159160 122894 159216
rect 127070 159432 127126 159488
rect 126426 152632 126482 152688
rect 126242 152360 126298 152416
rect 127070 153040 127126 153096
rect 128818 152496 128874 152552
rect 132038 153856 132094 153912
rect 131394 153040 131450 153096
rect 134614 153720 134670 153776
rect 135442 159296 135498 159352
rect 137374 159468 137376 159488
rect 137376 159468 137428 159488
rect 137428 159468 137430 159488
rect 137374 159432 137430 159468
rect 137098 153856 137154 153912
rect 138018 159432 138074 159488
rect 137650 153856 137706 153912
rect 139398 159568 139454 159624
rect 139950 156712 140006 156768
rect 139766 153992 139822 154048
rect 142986 156576 143042 156632
rect 143630 152632 143686 152688
rect 144918 157936 144974 157992
rect 149610 158208 149666 158264
rect 152554 158072 152610 158128
rect 150714 156848 150770 156904
rect 157154 159588 157210 159624
rect 157154 159568 157156 159588
rect 157156 159568 157208 159588
rect 157208 159568 157210 159588
rect 157338 159568 157394 159624
rect 156418 156984 156474 157040
rect 158350 154128 158406 154184
rect 160926 154264 160982 154320
rect 162858 158344 162914 158400
rect 166078 155216 166134 155272
rect 169298 157120 169354 157176
rect 171138 155488 171194 155544
rect 171230 155352 171286 155408
rect 177026 155624 177082 155680
rect 184018 155760 184074 155816
rect 185214 154284 185270 154320
rect 185214 154264 185216 154284
rect 185216 154264 185268 154284
rect 185268 154264 185270 154284
rect 186226 154980 186228 155000
rect 186228 154980 186280 155000
rect 186280 154980 186282 155000
rect 186226 154944 186282 154980
rect 186594 154980 186596 155000
rect 186596 154980 186648 155000
rect 186648 154980 186650 155000
rect 186594 154944 186650 154980
rect 187238 154400 187294 154456
rect 188342 153448 188398 153504
rect 189170 155896 189226 155952
rect 191470 154264 191526 154320
rect 192390 153448 192446 153504
rect 198738 158480 198794 158536
rect 204718 159296 204774 159352
rect 204258 157256 204314 157312
rect 212354 153720 212410 153776
rect 227442 152360 227498 152416
rect 274546 159432 274602 159488
rect 275190 159296 275246 159352
rect 278686 159060 278688 159080
rect 278688 159060 278740 159080
rect 278740 159060 278742 159080
rect 278686 159024 278742 159060
rect 280066 159060 280068 159080
rect 280068 159060 280120 159080
rect 280120 159060 280122 159080
rect 280066 159024 280122 159060
rect 280986 153720 281042 153776
rect 292578 152360 292634 152416
rect 313462 152360 313518 152416
rect 328550 159432 328606 159488
rect 357438 152360 357494 152416
rect 408314 152360 408370 152416
rect 430578 152360 430634 152416
rect 431866 152360 431922 152416
rect 448610 152360 448666 152416
rect 519726 163104 519782 163160
rect 519542 161608 519598 161664
rect 519450 151000 519506 151056
rect 519358 143384 519414 143440
rect 519266 138896 519322 138952
rect 519634 160112 519690 160168
rect 519542 147872 519598 147928
rect 519818 158616 519874 158672
rect 519726 149232 519782 149288
rect 519726 148008 519782 148064
rect 519634 146512 519690 146568
rect 519542 144880 519598 144936
rect 519450 138352 519506 138408
rect 520186 157120 520242 157176
rect 520094 155624 520150 155680
rect 520002 153992 520058 154048
rect 519910 149504 519966 149560
rect 519818 145152 519874 145208
rect 521014 152496 521070 152552
rect 520922 146512 520978 146568
rect 520186 143792 520242 143848
rect 520094 142432 520150 142488
rect 520186 141888 520242 141944
rect 520002 141072 520058 141128
rect 520002 140392 520058 140448
rect 519910 136992 519966 137048
rect 519910 135768 519966 135824
rect 519726 135632 519782 135688
rect 519634 134272 519690 134328
rect 519542 132912 519598 132968
rect 519358 131416 519414 131472
rect 519542 129784 519598 129840
rect 519266 127336 519322 127392
rect 519450 126656 519506 126712
rect 519358 125160 519414 125216
rect 519726 132776 519782 132832
rect 519634 123256 519690 123312
rect 519818 131280 519874 131336
rect 519726 121896 519782 121952
rect 519634 120672 519690 120728
rect 519542 119176 519598 119232
rect 519450 116456 519506 116512
rect 519358 115096 519414 115152
rect 519542 114552 519598 114608
rect 520094 137400 520150 137456
rect 520002 128696 520058 128752
rect 520002 128288 520058 128344
rect 519910 124616 519966 124672
rect 519818 120536 519874 120592
rect 519726 119176 519782 119232
rect 519634 110880 519690 110936
rect 521014 139712 521070 139768
rect 520922 134408 520978 134464
rect 520186 130056 520242 130112
rect 520094 125976 520150 126032
rect 520094 123664 520150 123720
rect 520002 117816 520058 117872
rect 519818 117544 519874 117600
rect 519726 109520 519782 109576
rect 519910 116048 519966 116104
rect 519818 108160 519874 108216
rect 520186 122168 520242 122224
rect 520094 113736 520150 113792
rect 521014 113056 521070 113112
rect 520186 112240 520242 112296
rect 520922 110064 520978 110120
rect 519910 106800 519966 106856
rect 519542 105440 519598 105496
rect 520278 105440 520334 105496
rect 117134 104760 117190 104816
rect 117042 102856 117098 102912
rect 116950 100952 117006 101008
rect 519818 99320 519874 99376
rect 116858 99048 116914 99104
rect 519726 97824 519782 97880
rect 116766 97144 116822 97200
rect 116674 95240 116730 95296
rect 519266 94832 519322 94888
rect 116582 93336 116638 93392
rect 116122 91296 116178 91352
rect 116122 89392 116178 89448
rect 519450 91840 519506 91896
rect 519266 87624 519322 87680
rect 116030 87488 116086 87544
rect 114466 87236 114522 87272
rect 114466 87216 114468 87236
rect 114468 87216 114520 87236
rect 114520 87216 114522 87236
rect 116214 85584 116270 85640
rect 116306 81776 116362 81832
rect 115938 79872 115994 79928
rect 520738 102448 520794 102504
rect 520278 97280 520334 97336
rect 520094 96328 520150 96384
rect 520002 93336 520058 93392
rect 519818 91704 519874 91760
rect 519726 90344 519782 90400
rect 519910 90208 519966 90264
rect 519726 87216 519782 87272
rect 519450 84904 519506 84960
rect 519266 84224 519322 84280
rect 116582 83680 116638 83736
rect 519450 81096 519506 81152
rect 519266 78104 519322 78160
rect 116490 77968 116546 78024
rect 519818 85720 519874 85776
rect 519726 80824 519782 80880
rect 519634 79600 519690 79656
rect 519450 75248 519506 75304
rect 116674 74024 116730 74080
rect 116582 72120 116638 72176
rect 39118 2644 39174 2680
rect 39118 2624 39120 2644
rect 39120 2624 39172 2644
rect 39172 2624 39174 2644
rect 19338 1808 19394 1864
rect 15934 1672 15990 1728
rect 12622 1536 12678 1592
rect 9310 1400 9366 1456
rect 53470 2644 53526 2680
rect 53470 2624 53472 2644
rect 53472 2624 53524 2644
rect 53524 2624 53526 2644
rect 81254 2644 81310 2680
rect 81254 2624 81256 2644
rect 81256 2624 81308 2644
rect 81308 2624 81310 2644
rect 106094 2644 106150 2680
rect 106094 2624 106096 2644
rect 106096 2624 106148 2644
rect 106148 2624 106150 2644
rect 109590 2624 109646 2680
rect 42798 2488 42854 2544
rect 50894 2488 50950 2544
rect 49146 2352 49202 2408
rect 58622 2488 58678 2544
rect 62394 2352 62450 2408
rect 63038 2352 63094 2408
rect 78034 2352 78090 2408
rect 78126 2216 78182 2272
rect 79782 2352 79838 2408
rect 79690 2216 79746 2272
rect 82266 2488 82322 2544
rect 116306 70216 116362 70272
rect 116122 68312 116178 68368
rect 116582 66408 116638 66464
rect 521106 111560 521162 111616
rect 521014 104080 521070 104136
rect 521198 108432 521254 108488
rect 521106 102720 521162 102776
rect 520922 101360 520978 101416
rect 521106 100952 521162 101008
rect 520738 94424 520794 94480
rect 521474 106936 521530 106992
rect 521290 103944 521346 104000
rect 521198 100000 521254 100056
rect 521474 98640 521530 98696
rect 521290 95920 521346 95976
rect 521106 93064 521162 93120
rect 520094 88984 520150 89040
rect 520186 88712 520242 88768
rect 520002 86264 520058 86320
rect 519910 83544 519966 83600
rect 520094 82728 520150 82784
rect 519818 79464 519874 79520
rect 519726 78104 519782 78160
rect 519634 73888 519690 73944
rect 520186 82184 520242 82240
rect 520094 76744 520150 76800
rect 520002 76608 520058 76664
rect 519818 75112 519874 75168
rect 519726 72528 519782 72584
rect 519910 73616 519966 73672
rect 519818 69808 519874 69864
rect 519634 68992 519690 69048
rect 114466 64540 114468 64560
rect 114468 64540 114520 64560
rect 114520 64540 114522 64560
rect 114466 64504 114522 64540
rect 116214 64504 116270 64560
rect 520094 71984 520150 72040
rect 520002 71168 520058 71224
rect 519910 68448 519966 68504
rect 520186 70488 520242 70544
rect 520094 67088 520150 67144
rect 520462 67496 520518 67552
rect 520370 66000 520426 66056
rect 520186 65728 520242 65784
rect 519634 64368 519690 64424
rect 116582 62600 116638 62656
rect 114190 53080 114246 53136
rect 116490 47096 116546 47152
rect 116214 45192 116270 45248
rect 114098 41792 114154 41848
rect 116122 41420 116124 41440
rect 116124 41420 116176 41440
rect 116176 41420 116178 41440
rect 116122 41384 116178 41420
rect 114006 30368 114062 30424
rect 113914 18944 113970 19000
rect 113822 7656 113878 7712
rect 116306 43288 116362 43344
rect 116214 37576 116270 37632
rect 116122 35672 116178 35728
rect 116122 33768 116178 33824
rect 116122 31764 116124 31784
rect 116124 31764 116176 31784
rect 116176 31764 116178 31784
rect 116122 31728 116178 31764
rect 116122 29824 116178 29880
rect 116122 27920 116178 27976
rect 116122 26016 116178 26072
rect 116122 24112 116178 24168
rect 116030 22208 116086 22264
rect 116214 20304 116270 20360
rect 116122 18400 116178 18456
rect 115938 14456 115994 14512
rect 116214 16360 116270 16416
rect 116398 39480 116454 39536
rect 116122 4936 116178 4992
rect 116122 3032 116178 3088
rect 520738 64504 520794 64560
rect 520462 63008 520518 63064
rect 520370 61648 520426 61704
rect 116674 60560 116730 60616
rect 521106 62872 521162 62928
rect 521014 61376 521070 61432
rect 520738 60288 520794 60344
rect 520738 59880 520794 59936
rect 116766 58656 116822 58712
rect 520370 56888 520426 56944
rect 116858 56752 116914 56808
rect 520278 55392 520334 55448
rect 116950 54848 117006 54904
rect 519082 53760 519138 53816
rect 117042 52944 117098 53000
rect 117134 51040 117190 51096
rect 519910 52264 519966 52320
rect 519082 50632 519138 50688
rect 521106 58928 521162 58984
rect 521106 58384 521162 58440
rect 521014 57432 521070 57488
rect 520738 56072 520794 56128
rect 521106 54712 521162 54768
rect 520370 53352 520426 53408
rect 520278 51992 520334 52048
rect 520002 50768 520058 50824
rect 519910 49272 519966 49328
rect 117226 49136 117282 49192
rect 520186 49272 520242 49328
rect 520002 47912 520058 47968
rect 519266 47776 519322 47832
rect 520186 46552 520242 46608
rect 519910 46280 519966 46336
rect 519266 45192 519322 45248
rect 519818 44648 519874 44704
rect 519910 43832 519966 43888
rect 520094 43152 520150 43208
rect 519818 42472 519874 42528
rect 520186 41656 520242 41712
rect 520094 41112 520150 41168
rect 519818 40160 519874 40216
rect 520186 39752 520242 39808
rect 520186 38664 520242 38720
rect 519818 38256 519874 38312
rect 521106 37168 521162 37224
rect 520186 36896 520242 36952
rect 521106 35944 521162 36000
rect 520922 35536 520978 35592
rect 520922 34584 520978 34640
rect 520830 34040 520886 34096
rect 520830 33224 520886 33280
rect 521106 32544 521162 32600
rect 521106 31728 521162 31784
rect 521106 31048 521162 31104
rect 521106 30368 521162 30424
rect 521106 29552 521162 29608
rect 521106 28736 521162 28792
rect 521106 20440 521162 20496
rect 521106 19760 521162 19816
rect 521106 15000 521162 15056
rect 521106 14320 521162 14376
rect 521106 13640 521162 13696
rect 521106 12824 521162 12880
rect 519634 12280 519690 12336
rect 519634 11328 519690 11384
rect 521106 10920 521162 10976
rect 521106 9832 521162 9888
rect 521106 9560 521162 9616
rect 520370 8200 520426 8256
rect 521106 8200 521162 8256
rect 521106 6840 521162 6896
rect 520370 6704 520426 6760
rect 521014 5480 521070 5536
rect 521106 5208 521162 5264
rect 521106 4120 521162 4176
rect 521014 3712 521070 3768
rect 520002 2760 520058 2816
rect 163778 1400 163834 1456
rect 229282 1536 229338 1592
rect 293590 1536 293646 1592
rect 243634 1400 243690 1456
rect 360290 1400 360346 1456
rect 393594 1400 393650 1456
rect 521106 2216 521162 2272
rect 520002 720 520058 776
<< metal3 >>
rect 519721 163162 519787 163165
rect 523200 163162 524400 163192
rect 519721 163160 524400 163162
rect 519721 163104 519726 163160
rect 519782 163104 524400 163160
rect 519721 163102 524400 163104
rect 519721 163099 519787 163102
rect 523200 163072 524400 163102
rect 519537 161666 519603 161669
rect 523200 161666 524400 161696
rect 519537 161664 524400 161666
rect 519537 161608 519542 161664
rect 519598 161608 524400 161664
rect 519537 161606 524400 161608
rect 519537 161603 519603 161606
rect 523200 161576 524400 161606
rect 519629 160170 519695 160173
rect 523200 160170 524400 160200
rect 519629 160168 524400 160170
rect 519629 160112 519634 160168
rect 519690 160112 524400 160168
rect 519629 160110 524400 160112
rect 519629 160107 519695 160110
rect 523200 160080 524400 160110
rect 29821 159626 29887 159629
rect 139393 159626 139459 159629
rect 29821 159624 139459 159626
rect 29821 159568 29826 159624
rect 29882 159568 139398 159624
rect 139454 159568 139459 159624
rect 29821 159566 139459 159568
rect 29821 159563 29887 159566
rect 139393 159563 139459 159566
rect 157149 159626 157215 159629
rect 157333 159626 157399 159629
rect 157149 159624 157399 159626
rect 157149 159568 157154 159624
rect 157210 159568 157338 159624
rect 157394 159568 157399 159624
rect 157149 159566 157399 159568
rect 157149 159563 157215 159566
rect 157333 159563 157399 159566
rect 16297 159490 16363 159493
rect 127065 159490 127131 159493
rect 16297 159488 127131 159490
rect 16297 159432 16302 159488
rect 16358 159432 127070 159488
rect 127126 159432 127131 159488
rect 16297 159430 127131 159432
rect 16297 159427 16363 159430
rect 127065 159427 127131 159430
rect 137369 159490 137435 159493
rect 138013 159490 138079 159493
rect 137369 159488 138079 159490
rect 137369 159432 137374 159488
rect 137430 159432 138018 159488
rect 138074 159432 138079 159488
rect 137369 159430 138079 159432
rect 137369 159427 137435 159430
rect 138013 159427 138079 159430
rect 274541 159490 274607 159493
rect 328545 159490 328611 159493
rect 274541 159488 328611 159490
rect 274541 159432 274546 159488
rect 274602 159432 328550 159488
rect 328606 159432 328611 159488
rect 274541 159430 328611 159432
rect 274541 159427 274607 159430
rect 328545 159427 328611 159430
rect 23013 159354 23079 159357
rect 135437 159354 135503 159357
rect 23013 159352 135503 159354
rect 23013 159296 23018 159352
rect 23074 159296 135442 159352
rect 135498 159296 135503 159352
rect 23013 159294 135503 159296
rect 23013 159291 23079 159294
rect 135437 159291 135503 159294
rect 204713 159354 204779 159357
rect 275185 159354 275251 159357
rect 204713 159352 275251 159354
rect 204713 159296 204718 159352
rect 204774 159296 275190 159352
rect 275246 159296 275251 159352
rect 204713 159294 275251 159296
rect 204713 159291 204779 159294
rect 275185 159291 275251 159294
rect 122649 159218 122715 159221
rect 122833 159218 122899 159221
rect 122649 159216 122899 159218
rect 122649 159160 122654 159216
rect 122710 159160 122838 159216
rect 122894 159160 122899 159216
rect 122649 159158 122899 159160
rect 122649 159155 122715 159158
rect 122833 159155 122899 159158
rect 278681 159082 278747 159085
rect 280061 159082 280127 159085
rect 278681 159080 280127 159082
rect 278681 159024 278686 159080
rect 278742 159024 280066 159080
rect 280122 159024 280127 159080
rect 278681 159022 280127 159024
rect 278681 159019 278747 159022
rect 280061 159019 280127 159022
rect 120533 158946 120599 158949
rect 121545 158946 121611 158949
rect 120533 158944 121611 158946
rect 120533 158888 120538 158944
rect 120594 158888 121550 158944
rect 121606 158888 121611 158944
rect 120533 158886 121611 158888
rect 120533 158883 120599 158886
rect 121545 158883 121611 158886
rect 519813 158674 519879 158677
rect 523200 158674 524400 158704
rect 519813 158672 524400 158674
rect 519813 158616 519818 158672
rect 519874 158616 524400 158672
rect 519813 158614 524400 158616
rect 519813 158611 519879 158614
rect 523200 158584 524400 158614
rect 104617 158538 104683 158541
rect 198733 158538 198799 158541
rect 104617 158536 198799 158538
rect 104617 158480 104622 158536
rect 104678 158480 198738 158536
rect 198794 158480 198799 158536
rect 104617 158478 198799 158480
rect 104617 158475 104683 158478
rect 198733 158475 198799 158478
rect 57513 158402 57579 158405
rect 162853 158402 162919 158405
rect 57513 158400 162919 158402
rect 57513 158344 57518 158400
rect 57574 158344 162858 158400
rect 162914 158344 162919 158400
rect 57513 158342 162919 158344
rect 57513 158339 57579 158342
rect 162853 158339 162919 158342
rect 40677 158266 40743 158269
rect 149605 158266 149671 158269
rect 40677 158264 149671 158266
rect 40677 158208 40682 158264
rect 40738 158208 149610 158264
rect 149666 158208 149671 158264
rect 40677 158206 149671 158208
rect 40677 158203 40743 158206
rect 149605 158203 149671 158206
rect 44081 158130 44147 158133
rect 152549 158130 152615 158133
rect 44081 158128 152615 158130
rect 44081 158072 44086 158128
rect 44142 158072 152554 158128
rect 152610 158072 152615 158128
rect 44081 158070 152615 158072
rect 44081 158067 44147 158070
rect 152549 158067 152615 158070
rect 33961 157994 34027 157997
rect 144913 157994 144979 157997
rect 33961 157992 144979 157994
rect 33961 157936 33966 157992
rect 34022 157936 144918 157992
rect 144974 157936 144979 157992
rect 33961 157934 144979 157936
rect 33961 157931 34027 157934
rect 144913 157931 144979 157934
rect 113081 157314 113147 157317
rect 204253 157314 204319 157317
rect 113081 157312 204319 157314
rect 113081 157256 113086 157312
rect 113142 157256 204258 157312
rect 204314 157256 204319 157312
rect 113081 157254 204319 157256
rect 113081 157251 113147 157254
rect 204253 157251 204319 157254
rect 65977 157178 66043 157181
rect 169293 157178 169359 157181
rect 65977 157176 169359 157178
rect 65977 157120 65982 157176
rect 66038 157120 169298 157176
rect 169354 157120 169359 157176
rect 65977 157118 169359 157120
rect 65977 157115 66043 157118
rect 169293 157115 169359 157118
rect 520181 157178 520247 157181
rect 523200 157178 524400 157208
rect 520181 157176 524400 157178
rect 520181 157120 520186 157176
rect 520242 157120 524400 157176
rect 520181 157118 524400 157120
rect 520181 157115 520247 157118
rect 523200 157088 524400 157118
rect 49141 157042 49207 157045
rect 156413 157042 156479 157045
rect 49141 157040 156479 157042
rect 49141 156984 49146 157040
rect 49202 156984 156418 157040
rect 156474 156984 156479 157040
rect 49141 156982 156479 156984
rect 49141 156979 49207 156982
rect 156413 156979 156479 156982
rect 42425 156906 42491 156909
rect 150709 156906 150775 156909
rect 42425 156904 150775 156906
rect 42425 156848 42430 156904
rect 42486 156848 150714 156904
rect 150770 156848 150775 156904
rect 42425 156846 150775 156848
rect 42425 156843 42491 156846
rect 150709 156843 150775 156846
rect 28073 156770 28139 156773
rect 139945 156770 140011 156773
rect 28073 156768 140011 156770
rect 28073 156712 28078 156768
rect 28134 156712 139950 156768
rect 140006 156712 140011 156768
rect 28073 156710 140011 156712
rect 28073 156707 28139 156710
rect 139945 156707 140011 156710
rect 31477 156634 31543 156637
rect 142981 156634 143047 156637
rect 31477 156632 143047 156634
rect 31477 156576 31482 156632
rect 31538 156576 142986 156632
rect 143042 156576 143047 156632
rect 31477 156574 143047 156576
rect 31477 156571 31543 156574
rect 142981 156571 143047 156574
rect 92013 155954 92079 155957
rect 189165 155954 189231 155957
rect 92013 155952 189231 155954
rect 92013 155896 92018 155952
rect 92074 155896 189170 155952
rect 189226 155896 189231 155952
rect 92013 155894 189231 155896
rect 92013 155891 92079 155894
rect 189165 155891 189231 155894
rect 85297 155818 85363 155821
rect 184013 155818 184079 155821
rect 85297 155816 184079 155818
rect 85297 155760 85302 155816
rect 85358 155760 184018 155816
rect 184074 155760 184079 155816
rect 85297 155758 184079 155760
rect 85297 155755 85363 155758
rect 184013 155755 184079 155758
rect 76005 155682 76071 155685
rect 177021 155682 177087 155685
rect 76005 155680 177087 155682
rect 76005 155624 76010 155680
rect 76066 155624 177026 155680
rect 177082 155624 177087 155680
rect 76005 155622 177087 155624
rect 76005 155619 76071 155622
rect 177021 155619 177087 155622
rect 520089 155682 520155 155685
rect 523200 155682 524400 155712
rect 520089 155680 524400 155682
rect 520089 155624 520094 155680
rect 520150 155624 524400 155680
rect 520089 155622 524400 155624
rect 520089 155619 520155 155622
rect 523200 155592 524400 155622
rect 69289 155546 69355 155549
rect 171133 155546 171199 155549
rect 69289 155544 171199 155546
rect 69289 155488 69294 155544
rect 69350 155488 171138 155544
rect 171194 155488 171199 155544
rect 69289 155486 171199 155488
rect 69289 155483 69355 155486
rect 171133 155483 171199 155486
rect 68461 155410 68527 155413
rect 171225 155410 171291 155413
rect 68461 155408 171291 155410
rect 68461 155352 68466 155408
rect 68522 155352 171230 155408
rect 171286 155352 171291 155408
rect 68461 155350 171291 155352
rect 68461 155347 68527 155350
rect 171225 155347 171291 155350
rect 61745 155274 61811 155277
rect 166073 155274 166139 155277
rect 61745 155272 166139 155274
rect 61745 155216 61750 155272
rect 61806 155216 166078 155272
rect 166134 155216 166139 155272
rect 61745 155214 166139 155216
rect 61745 155211 61811 155214
rect 166073 155211 166139 155214
rect 186221 155002 186287 155005
rect 186589 155002 186655 155005
rect 186221 155000 186655 155002
rect 186221 154944 186226 155000
rect 186282 154944 186594 155000
rect 186650 154944 186655 155000
rect 186221 154942 186655 154944
rect 186221 154939 186287 154942
rect 186589 154939 186655 154942
rect 89713 154458 89779 154461
rect 187233 154458 187299 154461
rect 89713 154456 187299 154458
rect 89713 154400 89718 154456
rect 89774 154400 187238 154456
rect 187294 154400 187299 154456
rect 89713 154398 187299 154400
rect 89713 154395 89779 154398
rect 187233 154395 187299 154398
rect 55029 154322 55095 154325
rect 160921 154322 160987 154325
rect 55029 154320 160987 154322
rect 55029 154264 55034 154320
rect 55090 154264 160926 154320
rect 160982 154264 160987 154320
rect 55029 154262 160987 154264
rect 55029 154259 55095 154262
rect 160921 154259 160987 154262
rect 185209 154322 185275 154325
rect 191465 154322 191531 154325
rect 185209 154320 191531 154322
rect 185209 154264 185214 154320
rect 185270 154264 191470 154320
rect 191526 154264 191531 154320
rect 185209 154262 191531 154264
rect 185209 154259 185275 154262
rect 191465 154259 191531 154262
rect 51625 154186 51691 154189
rect 158345 154186 158411 154189
rect 51625 154184 158411 154186
rect 51625 154128 51630 154184
rect 51686 154128 158350 154184
rect 158406 154128 158411 154184
rect 51625 154126 158411 154128
rect 51625 154123 51691 154126
rect 158345 154123 158411 154126
rect 27245 154050 27311 154053
rect 139761 154050 139827 154053
rect 27245 154048 139827 154050
rect 27245 153992 27250 154048
rect 27306 153992 139766 154048
rect 139822 153992 139827 154048
rect 27245 153990 139827 153992
rect 27245 153987 27311 153990
rect 139761 153987 139827 153990
rect 519997 154050 520063 154053
rect 523200 154050 524400 154080
rect 519997 154048 524400 154050
rect 519997 153992 520002 154048
rect 520058 153992 524400 154048
rect 519997 153990 524400 153992
rect 519997 153987 520063 153990
rect 523200 153960 524400 153990
rect 17125 153914 17191 153917
rect 132033 153914 132099 153917
rect 17125 153912 132099 153914
rect 17125 153856 17130 153912
rect 17186 153856 132038 153912
rect 132094 153856 132099 153912
rect 17125 153854 132099 153856
rect 17125 153851 17191 153854
rect 132033 153851 132099 153854
rect 137093 153914 137159 153917
rect 137645 153914 137711 153917
rect 137093 153912 137711 153914
rect 137093 153856 137098 153912
rect 137154 153856 137650 153912
rect 137706 153856 137711 153912
rect 137093 153854 137711 153856
rect 137093 153851 137159 153854
rect 137645 153851 137711 153854
rect 20529 153778 20595 153781
rect 134609 153778 134675 153781
rect 20529 153776 134675 153778
rect 20529 153720 20534 153776
rect 20590 153720 134614 153776
rect 134670 153720 134675 153776
rect 20529 153718 134675 153720
rect 20529 153715 20595 153718
rect 134609 153715 134675 153718
rect 212349 153778 212415 153781
rect 280981 153778 281047 153781
rect 212349 153776 281047 153778
rect 212349 153720 212354 153776
rect 212410 153720 280986 153776
rect 281042 153720 281047 153776
rect 212349 153718 281047 153720
rect 212349 153715 212415 153718
rect 280981 153715 281047 153718
rect 116393 153642 116459 153645
rect 119429 153642 119495 153645
rect 116393 153640 119495 153642
rect 116393 153584 116398 153640
rect 116454 153584 119434 153640
rect 119490 153584 119495 153640
rect 116393 153582 119495 153584
rect 116393 153579 116459 153582
rect 119429 153579 119495 153582
rect 188337 153506 188403 153509
rect 192385 153506 192451 153509
rect 188337 153504 192451 153506
rect 188337 153448 188342 153504
rect 188398 153448 192390 153504
rect 192446 153448 192451 153504
rect 188337 153446 192451 153448
rect 188337 153443 188403 153446
rect 192385 153443 192451 153446
rect 127065 153098 127131 153101
rect 131389 153098 131455 153101
rect 127065 153096 131455 153098
rect 127065 153040 127070 153096
rect 127126 153040 131394 153096
rect 131450 153040 131455 153096
rect 127065 153038 131455 153040
rect 127065 153035 127131 153038
rect 131389 153035 131455 153038
rect 126421 152690 126487 152693
rect 143625 152690 143691 152693
rect 126421 152688 143691 152690
rect 126421 152632 126426 152688
rect 126482 152632 143630 152688
rect 143686 152632 143691 152688
rect 126421 152630 143691 152632
rect 126421 152627 126487 152630
rect 143625 152627 143691 152630
rect 12985 152554 13051 152557
rect 128813 152554 128879 152557
rect 12985 152552 128879 152554
rect 12985 152496 12990 152552
rect 13046 152496 128818 152552
rect 128874 152496 128879 152552
rect 12985 152494 128879 152496
rect 12985 152491 13051 152494
rect 128813 152491 128879 152494
rect 521009 152554 521075 152557
rect 523200 152554 524400 152584
rect 521009 152552 524400 152554
rect 521009 152496 521014 152552
rect 521070 152496 524400 152552
rect 521009 152494 524400 152496
rect 521009 152491 521075 152494
rect 523200 152464 524400 152494
rect 9581 152418 9647 152421
rect 126237 152418 126303 152421
rect 9581 152416 126303 152418
rect 9581 152360 9586 152416
rect 9642 152360 126242 152416
rect 126298 152360 126303 152416
rect 9581 152358 126303 152360
rect 9581 152355 9647 152358
rect 126237 152355 126303 152358
rect 227437 152418 227503 152421
rect 292573 152418 292639 152421
rect 227437 152416 292639 152418
rect 227437 152360 227442 152416
rect 227498 152360 292578 152416
rect 292634 152360 292639 152416
rect 227437 152358 292639 152360
rect 227437 152355 227503 152358
rect 292573 152355 292639 152358
rect 313457 152418 313523 152421
rect 357433 152418 357499 152421
rect 313457 152416 357499 152418
rect 313457 152360 313462 152416
rect 313518 152360 357438 152416
rect 357494 152360 357499 152416
rect 313457 152358 357499 152360
rect 313457 152355 313523 152358
rect 357433 152355 357499 152358
rect 408309 152418 408375 152421
rect 430573 152418 430639 152421
rect 408309 152416 430639 152418
rect 408309 152360 408314 152416
rect 408370 152360 430578 152416
rect 430634 152360 430639 152416
rect 408309 152358 430639 152360
rect 408309 152355 408375 152358
rect 430573 152355 430639 152358
rect 431861 152418 431927 152421
rect 448605 152418 448671 152421
rect 431861 152416 448671 152418
rect 431861 152360 431866 152416
rect 431922 152360 448610 152416
rect 448666 152360 448671 152416
rect 431861 152358 448671 152360
rect 431861 152355 431927 152358
rect 448605 152355 448671 152358
rect 519445 151058 519511 151061
rect 523200 151058 524400 151088
rect 519445 151056 524400 151058
rect 519445 151000 519450 151056
rect 519506 151000 524400 151056
rect 519445 150998 524400 151000
rect 519445 150995 519511 150998
rect 523200 150968 524400 150998
rect 95785 149562 95851 149565
rect 102685 149562 102751 149565
rect 95785 149560 102751 149562
rect 95785 149504 95790 149560
rect 95846 149504 102690 149560
rect 102746 149504 102751 149560
rect 95785 149502 102751 149504
rect 95785 149499 95851 149502
rect 102685 149499 102751 149502
rect 519905 149562 519971 149565
rect 523200 149562 524400 149592
rect 519905 149560 524400 149562
rect 519905 149504 519910 149560
rect 519966 149504 524400 149560
rect 519905 149502 524400 149504
rect 519905 149499 519971 149502
rect 523200 149472 524400 149502
rect 99281 149426 99347 149429
rect 102869 149426 102935 149429
rect 99281 149424 102935 149426
rect 99281 149368 99286 149424
rect 99342 149368 102874 149424
rect 102930 149368 102935 149424
rect 99281 149366 102935 149368
rect 99281 149363 99347 149366
rect 102869 149363 102935 149366
rect 519721 149290 519787 149293
rect 518788 149288 519787 149290
rect 518788 149232 519726 149288
rect 519782 149232 519787 149288
rect 518788 149230 519787 149232
rect 519721 149227 519787 149230
rect 115933 149018 115999 149021
rect 115933 149016 119140 149018
rect 115933 148960 115938 149016
rect 115994 148960 119140 149016
rect 115933 148958 119140 148960
rect 115933 148955 115999 148958
rect 519721 148066 519787 148069
rect 523200 148066 524400 148096
rect 519721 148064 524400 148066
rect 519721 148008 519726 148064
rect 519782 148008 524400 148064
rect 519721 148006 524400 148008
rect 519721 148003 519787 148006
rect 523200 147976 524400 148006
rect 519537 147930 519603 147933
rect 518788 147928 519603 147930
rect 518788 147872 519542 147928
rect 519598 147872 519603 147928
rect 518788 147870 519603 147872
rect 519537 147867 519603 147870
rect 116117 147114 116183 147117
rect 116117 147112 119140 147114
rect 116117 147056 116122 147112
rect 116178 147056 119140 147112
rect 116117 147054 119140 147056
rect 116117 147051 116183 147054
rect 519629 146570 519695 146573
rect 518788 146568 519695 146570
rect 518788 146512 519634 146568
rect 519690 146512 519695 146568
rect 518788 146510 519695 146512
rect 519629 146507 519695 146510
rect 520917 146570 520983 146573
rect 523200 146570 524400 146600
rect 520917 146568 524400 146570
rect 520917 146512 520922 146568
rect 520978 146512 524400 146568
rect 520917 146510 524400 146512
rect 520917 146507 520983 146510
rect 523200 146480 524400 146510
rect 116025 145210 116091 145213
rect 519813 145210 519879 145213
rect 116025 145208 119140 145210
rect 116025 145152 116030 145208
rect 116086 145152 119140 145208
rect 116025 145150 119140 145152
rect 518788 145208 519879 145210
rect 518788 145152 519818 145208
rect 519874 145152 519879 145208
rect 518788 145150 519879 145152
rect 116025 145147 116091 145150
rect 519813 145147 519879 145150
rect 519537 144938 519603 144941
rect 523200 144938 524400 144968
rect 519537 144936 524400 144938
rect 519537 144880 519542 144936
rect 519598 144880 524400 144936
rect 519537 144878 524400 144880
rect 519537 144875 519603 144878
rect 523200 144848 524400 144878
rect 113817 144258 113883 144261
rect 110860 144256 113883 144258
rect 110860 144200 113822 144256
rect 113878 144200 113883 144256
rect 110860 144198 113883 144200
rect 113817 144195 113883 144198
rect 520181 143850 520247 143853
rect 518788 143848 520247 143850
rect 518788 143792 520186 143848
rect 520242 143792 520247 143848
rect 518788 143790 520247 143792
rect 520181 143787 520247 143790
rect 519353 143442 519419 143445
rect 523200 143442 524400 143472
rect 519353 143440 524400 143442
rect 519353 143384 519358 143440
rect 519414 143384 524400 143440
rect 519353 143382 524400 143384
rect 519353 143379 519419 143382
rect 523200 143352 524400 143382
rect 116209 143306 116275 143309
rect 116209 143304 119140 143306
rect 116209 143248 116214 143304
rect 116270 143248 119140 143304
rect 116209 143246 119140 143248
rect 116209 143243 116275 143246
rect 520089 142490 520155 142493
rect 518788 142488 520155 142490
rect 518788 142432 520094 142488
rect 520150 142432 520155 142488
rect 518788 142430 520155 142432
rect 520089 142427 520155 142430
rect 520181 141946 520247 141949
rect 523200 141946 524400 141976
rect 520181 141944 524400 141946
rect 520181 141888 520186 141944
rect 520242 141888 524400 141944
rect 520181 141886 524400 141888
rect 520181 141883 520247 141886
rect 523200 141856 524400 141886
rect 116485 141402 116551 141405
rect 116485 141400 119140 141402
rect 116485 141344 116490 141400
rect 116546 141344 119140 141400
rect 116485 141342 119140 141344
rect 116485 141339 116551 141342
rect 519997 141130 520063 141133
rect 518788 141128 520063 141130
rect 518788 141072 520002 141128
rect 520058 141072 520063 141128
rect 518788 141070 520063 141072
rect 519997 141067 520063 141070
rect 519997 140450 520063 140453
rect 523200 140450 524400 140480
rect 519997 140448 524400 140450
rect 519997 140392 520002 140448
rect 520058 140392 524400 140448
rect 519997 140390 524400 140392
rect 519997 140387 520063 140390
rect 523200 140360 524400 140390
rect 521009 139770 521075 139773
rect 518788 139768 521075 139770
rect 518788 139712 521014 139768
rect 521070 139712 521075 139768
rect 518788 139710 521075 139712
rect 521009 139707 521075 139710
rect 115933 139498 115999 139501
rect 115933 139496 119140 139498
rect 115933 139440 115938 139496
rect 115994 139440 119140 139496
rect 115933 139438 119140 139440
rect 115933 139435 115999 139438
rect 519261 138954 519327 138957
rect 523200 138954 524400 138984
rect 519261 138952 524400 138954
rect 519261 138896 519266 138952
rect 519322 138896 524400 138952
rect 519261 138894 524400 138896
rect 519261 138891 519327 138894
rect 523200 138864 524400 138894
rect 519445 138410 519511 138413
rect 518788 138408 519511 138410
rect 518788 138352 519450 138408
rect 519506 138352 519511 138408
rect 518788 138350 519511 138352
rect 519445 138347 519511 138350
rect 116393 137594 116459 137597
rect 116393 137592 119140 137594
rect 116393 137536 116398 137592
rect 116454 137536 119140 137592
rect 116393 137534 119140 137536
rect 116393 137531 116459 137534
rect 520089 137458 520155 137461
rect 523200 137458 524400 137488
rect 520089 137456 524400 137458
rect 520089 137400 520094 137456
rect 520150 137400 524400 137456
rect 520089 137398 524400 137400
rect 520089 137395 520155 137398
rect 523200 137368 524400 137398
rect 519905 137050 519971 137053
rect 518788 137048 519971 137050
rect 518788 136992 519910 137048
rect 519966 136992 519971 137048
rect 518788 136990 519971 136992
rect 519905 136987 519971 136990
rect 519905 135826 519971 135829
rect 523200 135826 524400 135856
rect 519905 135824 524400 135826
rect 519905 135768 519910 135824
rect 519966 135768 524400 135824
rect 519905 135766 524400 135768
rect 519905 135763 519971 135766
rect 523200 135736 524400 135766
rect 519721 135690 519787 135693
rect 518788 135688 519787 135690
rect 518788 135632 519726 135688
rect 519782 135632 519787 135688
rect 518788 135630 519787 135632
rect 519721 135627 519787 135630
rect 115933 135554 115999 135557
rect 115933 135552 119140 135554
rect 115933 135496 115938 135552
rect 115994 135496 119140 135552
rect 115933 135494 119140 135496
rect 115933 135491 115999 135494
rect 520917 134466 520983 134469
rect 518758 134464 520983 134466
rect 518758 134408 520922 134464
rect 520978 134408 520983 134464
rect 518758 134406 520983 134408
rect 518758 134300 518818 134406
rect 520917 134403 520983 134406
rect 519629 134330 519695 134333
rect 523200 134330 524400 134360
rect 519629 134328 524400 134330
rect 519629 134272 519634 134328
rect 519690 134272 524400 134328
rect 519629 134270 524400 134272
rect 519629 134267 519695 134270
rect 523200 134240 524400 134270
rect 116117 133650 116183 133653
rect 116117 133648 119140 133650
rect 116117 133592 116122 133648
rect 116178 133592 119140 133648
rect 116117 133590 119140 133592
rect 116117 133587 116183 133590
rect 519537 132970 519603 132973
rect 518788 132968 519603 132970
rect 518788 132912 519542 132968
rect 519598 132912 519603 132968
rect 518788 132910 519603 132912
rect 519537 132907 519603 132910
rect 113909 132834 113975 132837
rect 110860 132832 113975 132834
rect 110860 132776 113914 132832
rect 113970 132776 113975 132832
rect 110860 132774 113975 132776
rect 113909 132771 113975 132774
rect 519721 132834 519787 132837
rect 523200 132834 524400 132864
rect 519721 132832 524400 132834
rect 519721 132776 519726 132832
rect 519782 132776 524400 132832
rect 519721 132774 524400 132776
rect 519721 132771 519787 132774
rect 523200 132744 524400 132774
rect 116117 131746 116183 131749
rect 116117 131744 119140 131746
rect 116117 131688 116122 131744
rect 116178 131688 119140 131744
rect 116117 131686 119140 131688
rect 116117 131683 116183 131686
rect 519353 131474 519419 131477
rect 518788 131472 519419 131474
rect 518788 131416 519358 131472
rect 519414 131416 519419 131472
rect 518788 131414 519419 131416
rect 519353 131411 519419 131414
rect 519813 131338 519879 131341
rect 523200 131338 524400 131368
rect 519813 131336 524400 131338
rect 519813 131280 519818 131336
rect 519874 131280 524400 131336
rect 519813 131278 524400 131280
rect 519813 131275 519879 131278
rect 523200 131248 524400 131278
rect 520181 130114 520247 130117
rect 518788 130112 520247 130114
rect 518788 130056 520186 130112
rect 520242 130056 520247 130112
rect 518788 130054 520247 130056
rect 520181 130051 520247 130054
rect 116117 129842 116183 129845
rect 519537 129842 519603 129845
rect 523200 129842 524400 129872
rect 116117 129840 119140 129842
rect 116117 129784 116122 129840
rect 116178 129784 119140 129840
rect 116117 129782 119140 129784
rect 519537 129840 524400 129842
rect 519537 129784 519542 129840
rect 519598 129784 524400 129840
rect 519537 129782 524400 129784
rect 116117 129779 116183 129782
rect 519537 129779 519603 129782
rect 523200 129752 524400 129782
rect 519997 128754 520063 128757
rect 518788 128752 520063 128754
rect 518788 128696 520002 128752
rect 520058 128696 520063 128752
rect 518788 128694 520063 128696
rect 519997 128691 520063 128694
rect 519997 128346 520063 128349
rect 523200 128346 524400 128376
rect 519997 128344 524400 128346
rect 519997 128288 520002 128344
rect 520058 128288 524400 128344
rect 519997 128286 524400 128288
rect 519997 128283 520063 128286
rect 523200 128256 524400 128286
rect 116117 127938 116183 127941
rect 116117 127936 119140 127938
rect 116117 127880 116122 127936
rect 116178 127880 119140 127936
rect 116117 127878 119140 127880
rect 116117 127875 116183 127878
rect 519261 127394 519327 127397
rect 518788 127392 519327 127394
rect 518788 127336 519266 127392
rect 519322 127336 519327 127392
rect 518788 127334 519327 127336
rect 519261 127331 519327 127334
rect 519445 126714 519511 126717
rect 523200 126714 524400 126744
rect 519445 126712 524400 126714
rect 519445 126656 519450 126712
rect 519506 126656 524400 126712
rect 519445 126654 524400 126656
rect 519445 126651 519511 126654
rect 523200 126624 524400 126654
rect 116025 126034 116091 126037
rect 520089 126034 520155 126037
rect 116025 126032 119140 126034
rect 116025 125976 116030 126032
rect 116086 125976 119140 126032
rect 116025 125974 119140 125976
rect 518788 126032 520155 126034
rect 518788 125976 520094 126032
rect 520150 125976 520155 126032
rect 518788 125974 520155 125976
rect 116025 125971 116091 125974
rect 520089 125971 520155 125974
rect 519353 125218 519419 125221
rect 523200 125218 524400 125248
rect 519353 125216 524400 125218
rect 519353 125160 519358 125216
rect 519414 125160 524400 125216
rect 519353 125158 524400 125160
rect 519353 125155 519419 125158
rect 523200 125128 524400 125158
rect 519905 124674 519971 124677
rect 518788 124672 519971 124674
rect 518788 124616 519910 124672
rect 519966 124616 519971 124672
rect 518788 124614 519971 124616
rect 519905 124611 519971 124614
rect 116117 124130 116183 124133
rect 116117 124128 119140 124130
rect 116117 124072 116122 124128
rect 116178 124072 119140 124128
rect 116117 124070 119140 124072
rect 116117 124067 116183 124070
rect 520089 123722 520155 123725
rect 523200 123722 524400 123752
rect 520089 123720 524400 123722
rect 520089 123664 520094 123720
rect 520150 123664 524400 123720
rect 520089 123662 524400 123664
rect 520089 123659 520155 123662
rect 523200 123632 524400 123662
rect 519629 123314 519695 123317
rect 518788 123312 519695 123314
rect 518788 123256 519634 123312
rect 519690 123256 519695 123312
rect 518788 123254 519695 123256
rect 519629 123251 519695 123254
rect 115933 122226 115999 122229
rect 520181 122226 520247 122229
rect 523200 122226 524400 122256
rect 115933 122224 119140 122226
rect 115933 122168 115938 122224
rect 115994 122168 119140 122224
rect 115933 122166 119140 122168
rect 520181 122224 524400 122226
rect 520181 122168 520186 122224
rect 520242 122168 524400 122224
rect 520181 122166 524400 122168
rect 115933 122163 115999 122166
rect 520181 122163 520247 122166
rect 523200 122136 524400 122166
rect 519721 121954 519787 121957
rect 518788 121952 519787 121954
rect 518788 121896 519726 121952
rect 519782 121896 519787 121952
rect 518788 121894 519787 121896
rect 519721 121891 519787 121894
rect 114001 121410 114067 121413
rect 110860 121408 114067 121410
rect 110860 121352 114006 121408
rect 114062 121352 114067 121408
rect 110860 121350 114067 121352
rect 114001 121347 114067 121350
rect 519629 120730 519695 120733
rect 523200 120730 524400 120760
rect 519629 120728 524400 120730
rect 519629 120672 519634 120728
rect 519690 120672 524400 120728
rect 519629 120670 524400 120672
rect 519629 120667 519695 120670
rect 523200 120640 524400 120670
rect 519813 120594 519879 120597
rect 518788 120592 519879 120594
rect 518788 120536 519818 120592
rect 519874 120536 519879 120592
rect 518788 120534 519879 120536
rect 519813 120531 519879 120534
rect 116117 120186 116183 120189
rect 116117 120184 119140 120186
rect 116117 120128 116122 120184
rect 116178 120128 119140 120184
rect 116117 120126 119140 120128
rect 116117 120123 116183 120126
rect 519537 119234 519603 119237
rect 518788 119232 519603 119234
rect 518788 119176 519542 119232
rect 519598 119176 519603 119232
rect 518788 119174 519603 119176
rect 519537 119171 519603 119174
rect 519721 119234 519787 119237
rect 523200 119234 524400 119264
rect 519721 119232 524400 119234
rect 519721 119176 519726 119232
rect 519782 119176 524400 119232
rect 519721 119174 524400 119176
rect 519721 119171 519787 119174
rect 523200 119144 524400 119174
rect 116117 118282 116183 118285
rect 116117 118280 119140 118282
rect 116117 118224 116122 118280
rect 116178 118224 119140 118280
rect 116117 118222 119140 118224
rect 116117 118219 116183 118222
rect 519997 117874 520063 117877
rect 518788 117872 520063 117874
rect 518788 117816 520002 117872
rect 520058 117816 520063 117872
rect 518788 117814 520063 117816
rect 519997 117811 520063 117814
rect 519813 117602 519879 117605
rect 523200 117602 524400 117632
rect 519813 117600 524400 117602
rect 519813 117544 519818 117600
rect 519874 117544 524400 117600
rect 519813 117542 524400 117544
rect 519813 117539 519879 117542
rect 523200 117512 524400 117542
rect 519445 116514 519511 116517
rect 518788 116512 519511 116514
rect 518788 116456 519450 116512
rect 519506 116456 519511 116512
rect 518788 116454 519511 116456
rect 519445 116451 519511 116454
rect 116117 116378 116183 116381
rect 116117 116376 119140 116378
rect 116117 116320 116122 116376
rect 116178 116320 119140 116376
rect 116117 116318 119140 116320
rect 116117 116315 116183 116318
rect 519905 116106 519971 116109
rect 523200 116106 524400 116136
rect 519905 116104 524400 116106
rect 519905 116048 519910 116104
rect 519966 116048 524400 116104
rect 519905 116046 524400 116048
rect 519905 116043 519971 116046
rect 523200 116016 524400 116046
rect 519353 115154 519419 115157
rect 518788 115152 519419 115154
rect 518788 115096 519358 115152
rect 519414 115096 519419 115152
rect 518788 115094 519419 115096
rect 519353 115091 519419 115094
rect 519537 114610 519603 114613
rect 523200 114610 524400 114640
rect 519537 114608 524400 114610
rect 519537 114552 519542 114608
rect 519598 114552 524400 114608
rect 519537 114550 524400 114552
rect 519537 114547 519603 114550
rect 523200 114520 524400 114550
rect 116117 114474 116183 114477
rect 116117 114472 119140 114474
rect 116117 114416 116122 114472
rect 116178 114416 119140 114472
rect 116117 114414 119140 114416
rect 116117 114411 116183 114414
rect 520089 113794 520155 113797
rect 518788 113792 520155 113794
rect 518788 113736 520094 113792
rect 520150 113736 520155 113792
rect 518788 113734 520155 113736
rect 520089 113731 520155 113734
rect 521009 113114 521075 113117
rect 523200 113114 524400 113144
rect 521009 113112 524400 113114
rect 521009 113056 521014 113112
rect 521070 113056 524400 113112
rect 521009 113054 524400 113056
rect 521009 113051 521075 113054
rect 523200 113024 524400 113054
rect 115933 112570 115999 112573
rect 115933 112568 119140 112570
rect 115933 112512 115938 112568
rect 115994 112512 119140 112568
rect 115933 112510 119140 112512
rect 115933 112507 115999 112510
rect 520181 112298 520247 112301
rect 518788 112296 520247 112298
rect 518788 112240 520186 112296
rect 520242 112240 520247 112296
rect 518788 112238 520247 112240
rect 520181 112235 520247 112238
rect 521101 111618 521167 111621
rect 523200 111618 524400 111648
rect 521101 111616 524400 111618
rect 521101 111560 521106 111616
rect 521162 111560 524400 111616
rect 521101 111558 524400 111560
rect 521101 111555 521167 111558
rect 523200 111528 524400 111558
rect 519629 110938 519695 110941
rect 518788 110936 519695 110938
rect 518788 110880 519634 110936
rect 519690 110880 519695 110936
rect 518788 110878 519695 110880
rect 519629 110875 519695 110878
rect 116117 110666 116183 110669
rect 116117 110664 119140 110666
rect 116117 110608 116122 110664
rect 116178 110608 119140 110664
rect 116117 110606 119140 110608
rect 116117 110603 116183 110606
rect 114093 110122 114159 110125
rect 110860 110120 114159 110122
rect 110860 110064 114098 110120
rect 114154 110064 114159 110120
rect 110860 110062 114159 110064
rect 114093 110059 114159 110062
rect 520917 110122 520983 110125
rect 523200 110122 524400 110152
rect 520917 110120 524400 110122
rect 520917 110064 520922 110120
rect 520978 110064 524400 110120
rect 520917 110062 524400 110064
rect 520917 110059 520983 110062
rect 523200 110032 524400 110062
rect 519721 109578 519787 109581
rect 518788 109576 519787 109578
rect 518788 109520 519726 109576
rect 519782 109520 519787 109576
rect 518788 109518 519787 109520
rect 519721 109515 519787 109518
rect 116117 108762 116183 108765
rect 116117 108760 119140 108762
rect 116117 108704 116122 108760
rect 116178 108704 119140 108760
rect 116117 108702 119140 108704
rect 116117 108699 116183 108702
rect 521193 108490 521259 108493
rect 523200 108490 524400 108520
rect 521193 108488 524400 108490
rect 521193 108432 521198 108488
rect 521254 108432 524400 108488
rect 521193 108430 524400 108432
rect 521193 108427 521259 108430
rect 523200 108400 524400 108430
rect 519813 108218 519879 108221
rect 518788 108216 519879 108218
rect 518788 108160 519818 108216
rect 519874 108160 519879 108216
rect 518788 108158 519879 108160
rect 519813 108155 519879 108158
rect 521469 106994 521535 106997
rect 523200 106994 524400 107024
rect 521469 106992 524400 106994
rect 521469 106936 521474 106992
rect 521530 106936 524400 106992
rect 521469 106934 524400 106936
rect 521469 106931 521535 106934
rect 523200 106904 524400 106934
rect 116485 106858 116551 106861
rect 519905 106858 519971 106861
rect 116485 106856 119140 106858
rect 116485 106800 116490 106856
rect 116546 106800 119140 106856
rect 116485 106798 119140 106800
rect 518788 106856 519971 106858
rect 518788 106800 519910 106856
rect 519966 106800 519971 106856
rect 518788 106798 519971 106800
rect 116485 106795 116551 106798
rect 519905 106795 519971 106798
rect 519537 105498 519603 105501
rect 518788 105496 519603 105498
rect 518788 105440 519542 105496
rect 519598 105440 519603 105496
rect 518788 105438 519603 105440
rect 519537 105435 519603 105438
rect 520273 105498 520339 105501
rect 523200 105498 524400 105528
rect 520273 105496 524400 105498
rect 520273 105440 520278 105496
rect 520334 105440 524400 105496
rect 520273 105438 524400 105440
rect 520273 105435 520339 105438
rect 523200 105408 524400 105438
rect 117129 104818 117195 104821
rect 117129 104816 119140 104818
rect 117129 104760 117134 104816
rect 117190 104760 119140 104816
rect 117129 104758 119140 104760
rect 117129 104755 117195 104758
rect 521009 104138 521075 104141
rect 518788 104136 521075 104138
rect 518788 104080 521014 104136
rect 521070 104080 521075 104136
rect 518788 104078 521075 104080
rect 521009 104075 521075 104078
rect 521285 104002 521351 104005
rect 523200 104002 524400 104032
rect 521285 104000 524400 104002
rect 521285 103944 521290 104000
rect 521346 103944 524400 104000
rect 521285 103942 524400 103944
rect 521285 103939 521351 103942
rect 523200 103912 524400 103942
rect 117037 102914 117103 102917
rect 117037 102912 119140 102914
rect 117037 102856 117042 102912
rect 117098 102856 119140 102912
rect 117037 102854 119140 102856
rect 117037 102851 117103 102854
rect 521101 102778 521167 102781
rect 518788 102776 521167 102778
rect 518788 102720 521106 102776
rect 521162 102720 521167 102776
rect 518788 102718 521167 102720
rect 521101 102715 521167 102718
rect 520733 102506 520799 102509
rect 523200 102506 524400 102536
rect 520733 102504 524400 102506
rect 520733 102448 520738 102504
rect 520794 102448 524400 102504
rect 520733 102446 524400 102448
rect 520733 102443 520799 102446
rect 523200 102416 524400 102446
rect 520917 101418 520983 101421
rect 518788 101416 520983 101418
rect 518788 101360 520922 101416
rect 520978 101360 520983 101416
rect 518788 101358 520983 101360
rect 520917 101355 520983 101358
rect 116945 101010 117011 101013
rect 521101 101010 521167 101013
rect 523200 101010 524400 101040
rect 116945 101008 119140 101010
rect 116945 100952 116950 101008
rect 117006 100952 119140 101008
rect 116945 100950 119140 100952
rect 521101 101008 524400 101010
rect 521101 100952 521106 101008
rect 521162 100952 524400 101008
rect 521101 100950 524400 100952
rect 116945 100947 117011 100950
rect 521101 100947 521167 100950
rect 523200 100920 524400 100950
rect 521193 100058 521259 100061
rect 518788 100056 521259 100058
rect 518788 100000 521198 100056
rect 521254 100000 521259 100056
rect 518788 99998 521259 100000
rect 521193 99995 521259 99998
rect 519813 99378 519879 99381
rect 523200 99378 524400 99408
rect 519813 99376 524400 99378
rect 519813 99320 519818 99376
rect 519874 99320 524400 99376
rect 519813 99318 524400 99320
rect 519813 99315 519879 99318
rect 523200 99288 524400 99318
rect 116853 99106 116919 99109
rect 116853 99104 119140 99106
rect 116853 99048 116858 99104
rect 116914 99048 119140 99104
rect 116853 99046 119140 99048
rect 116853 99043 116919 99046
rect 114185 98698 114251 98701
rect 521469 98698 521535 98701
rect 110860 98696 114251 98698
rect 110860 98640 114190 98696
rect 114246 98640 114251 98696
rect 110860 98638 114251 98640
rect 518788 98696 521535 98698
rect 518788 98640 521474 98696
rect 521530 98640 521535 98696
rect 518788 98638 521535 98640
rect 114185 98635 114251 98638
rect 521469 98635 521535 98638
rect 519721 97882 519787 97885
rect 523200 97882 524400 97912
rect 519721 97880 524400 97882
rect 519721 97824 519726 97880
rect 519782 97824 524400 97880
rect 519721 97822 524400 97824
rect 519721 97819 519787 97822
rect 523200 97792 524400 97822
rect 520273 97338 520339 97341
rect 518788 97336 520339 97338
rect 518788 97280 520278 97336
rect 520334 97280 520339 97336
rect 518788 97278 520339 97280
rect 520273 97275 520339 97278
rect 116761 97202 116827 97205
rect 116761 97200 119140 97202
rect 116761 97144 116766 97200
rect 116822 97144 119140 97200
rect 116761 97142 119140 97144
rect 116761 97139 116827 97142
rect 520089 96386 520155 96389
rect 523200 96386 524400 96416
rect 520089 96384 524400 96386
rect 520089 96328 520094 96384
rect 520150 96328 524400 96384
rect 520089 96326 524400 96328
rect 520089 96323 520155 96326
rect 523200 96296 524400 96326
rect 521285 95978 521351 95981
rect 518788 95976 521351 95978
rect 518788 95920 521290 95976
rect 521346 95920 521351 95976
rect 518788 95918 521351 95920
rect 521285 95915 521351 95918
rect 116669 95298 116735 95301
rect 116669 95296 119140 95298
rect 116669 95240 116674 95296
rect 116730 95240 119140 95296
rect 116669 95238 119140 95240
rect 116669 95235 116735 95238
rect 519261 94890 519327 94893
rect 523200 94890 524400 94920
rect 519261 94888 524400 94890
rect 519261 94832 519266 94888
rect 519322 94832 524400 94888
rect 519261 94830 524400 94832
rect 519261 94827 519327 94830
rect 523200 94800 524400 94830
rect 520733 94482 520799 94485
rect 518788 94480 520799 94482
rect 518788 94424 520738 94480
rect 520794 94424 520799 94480
rect 518788 94422 520799 94424
rect 520733 94419 520799 94422
rect 116577 93394 116643 93397
rect 519997 93394 520063 93397
rect 523200 93394 524400 93424
rect 116577 93392 119140 93394
rect 116577 93336 116582 93392
rect 116638 93336 119140 93392
rect 116577 93334 119140 93336
rect 519997 93392 524400 93394
rect 519997 93336 520002 93392
rect 520058 93336 524400 93392
rect 519997 93334 524400 93336
rect 116577 93331 116643 93334
rect 519997 93331 520063 93334
rect 523200 93304 524400 93334
rect 521101 93122 521167 93125
rect 518788 93120 521167 93122
rect 518788 93064 521106 93120
rect 521162 93064 521167 93120
rect 518788 93062 521167 93064
rect 521101 93059 521167 93062
rect 519445 91898 519511 91901
rect 523200 91898 524400 91928
rect 519445 91896 524400 91898
rect 519445 91840 519450 91896
rect 519506 91840 524400 91896
rect 519445 91838 524400 91840
rect 519445 91835 519511 91838
rect 523200 91808 524400 91838
rect 519813 91762 519879 91765
rect 518788 91760 519879 91762
rect 518788 91704 519818 91760
rect 519874 91704 519879 91760
rect 518788 91702 519879 91704
rect 519813 91699 519879 91702
rect 116117 91354 116183 91357
rect 116117 91352 119140 91354
rect 116117 91296 116122 91352
rect 116178 91296 119140 91352
rect 116117 91294 119140 91296
rect 116117 91291 116183 91294
rect 519721 90402 519787 90405
rect 518788 90400 519787 90402
rect 518788 90344 519726 90400
rect 519782 90344 519787 90400
rect 518788 90342 519787 90344
rect 519721 90339 519787 90342
rect 519905 90266 519971 90269
rect 523200 90266 524400 90296
rect 519905 90264 524400 90266
rect 519905 90208 519910 90264
rect 519966 90208 524400 90264
rect 519905 90206 524400 90208
rect 519905 90203 519971 90206
rect 523200 90176 524400 90206
rect 116117 89450 116183 89453
rect 116117 89448 119140 89450
rect 116117 89392 116122 89448
rect 116178 89392 119140 89448
rect 116117 89390 119140 89392
rect 116117 89387 116183 89390
rect 520089 89042 520155 89045
rect 518788 89040 520155 89042
rect 518788 88984 520094 89040
rect 520150 88984 520155 89040
rect 518788 88982 520155 88984
rect 520089 88979 520155 88982
rect 520181 88770 520247 88773
rect 523200 88770 524400 88800
rect 520181 88768 524400 88770
rect 520181 88712 520186 88768
rect 520242 88712 524400 88768
rect 520181 88710 524400 88712
rect 520181 88707 520247 88710
rect 523200 88680 524400 88710
rect 519261 87682 519327 87685
rect 518788 87680 519327 87682
rect 518788 87624 519266 87680
rect 519322 87624 519327 87680
rect 518788 87622 519327 87624
rect 519261 87619 519327 87622
rect 116025 87546 116091 87549
rect 116025 87544 119140 87546
rect 116025 87488 116030 87544
rect 116086 87488 119140 87544
rect 116025 87486 119140 87488
rect 116025 87483 116091 87486
rect 114461 87274 114527 87277
rect 110860 87272 114527 87274
rect 110860 87216 114466 87272
rect 114522 87216 114527 87272
rect 110860 87214 114527 87216
rect 114461 87211 114527 87214
rect 519721 87274 519787 87277
rect 523200 87274 524400 87304
rect 519721 87272 524400 87274
rect 519721 87216 519726 87272
rect 519782 87216 524400 87272
rect 519721 87214 524400 87216
rect 519721 87211 519787 87214
rect 523200 87184 524400 87214
rect 519997 86322 520063 86325
rect 518788 86320 520063 86322
rect 518788 86264 520002 86320
rect 520058 86264 520063 86320
rect 518788 86262 520063 86264
rect 519997 86259 520063 86262
rect 519813 85778 519879 85781
rect 523200 85778 524400 85808
rect 519813 85776 524400 85778
rect 519813 85720 519818 85776
rect 519874 85720 524400 85776
rect 519813 85718 524400 85720
rect 519813 85715 519879 85718
rect 523200 85688 524400 85718
rect 116209 85642 116275 85645
rect 116209 85640 119140 85642
rect 116209 85584 116214 85640
rect 116270 85584 119140 85640
rect 116209 85582 119140 85584
rect 116209 85579 116275 85582
rect 519445 84962 519511 84965
rect 518788 84960 519511 84962
rect 518788 84904 519450 84960
rect 519506 84904 519511 84960
rect 518788 84902 519511 84904
rect 519445 84899 519511 84902
rect 519261 84282 519327 84285
rect 523200 84282 524400 84312
rect 519261 84280 524400 84282
rect 519261 84224 519266 84280
rect 519322 84224 524400 84280
rect 519261 84222 524400 84224
rect 519261 84219 519327 84222
rect 523200 84192 524400 84222
rect 116577 83738 116643 83741
rect 116577 83736 119140 83738
rect 116577 83680 116582 83736
rect 116638 83680 119140 83736
rect 116577 83678 119140 83680
rect 116577 83675 116643 83678
rect 519905 83602 519971 83605
rect 518788 83600 519971 83602
rect 518788 83544 519910 83600
rect 519966 83544 519971 83600
rect 518788 83542 519971 83544
rect 519905 83539 519971 83542
rect 520089 82786 520155 82789
rect 523200 82786 524400 82816
rect 520089 82784 524400 82786
rect 520089 82728 520094 82784
rect 520150 82728 524400 82784
rect 520089 82726 524400 82728
rect 520089 82723 520155 82726
rect 523200 82696 524400 82726
rect 520181 82242 520247 82245
rect 518788 82240 520247 82242
rect 518788 82184 520186 82240
rect 520242 82184 520247 82240
rect 518788 82182 520247 82184
rect 520181 82179 520247 82182
rect 116301 81834 116367 81837
rect 116301 81832 119140 81834
rect 116301 81776 116306 81832
rect 116362 81776 119140 81832
rect 116301 81774 119140 81776
rect 116301 81771 116367 81774
rect 519445 81154 519511 81157
rect 523200 81154 524400 81184
rect 519445 81152 524400 81154
rect 519445 81096 519450 81152
rect 519506 81096 524400 81152
rect 519445 81094 524400 81096
rect 519445 81091 519511 81094
rect 523200 81064 524400 81094
rect 519721 80882 519787 80885
rect 518788 80880 519787 80882
rect 518788 80824 519726 80880
rect 519782 80824 519787 80880
rect 518788 80822 519787 80824
rect 519721 80819 519787 80822
rect 115933 79930 115999 79933
rect 115933 79928 119140 79930
rect 115933 79872 115938 79928
rect 115994 79872 119140 79928
rect 115933 79870 119140 79872
rect 115933 79867 115999 79870
rect 519629 79658 519695 79661
rect 523200 79658 524400 79688
rect 519629 79656 524400 79658
rect 519629 79600 519634 79656
rect 519690 79600 524400 79656
rect 519629 79598 524400 79600
rect 519629 79595 519695 79598
rect 523200 79568 524400 79598
rect 519813 79522 519879 79525
rect 518788 79520 519879 79522
rect 518788 79464 519818 79520
rect 519874 79464 519879 79520
rect 518788 79462 519879 79464
rect 519813 79459 519879 79462
rect 519261 78162 519327 78165
rect 518788 78160 519327 78162
rect 518788 78104 519266 78160
rect 519322 78104 519327 78160
rect 518788 78102 519327 78104
rect 519261 78099 519327 78102
rect 519721 78162 519787 78165
rect 523200 78162 524400 78192
rect 519721 78160 524400 78162
rect 519721 78104 519726 78160
rect 519782 78104 524400 78160
rect 519721 78102 524400 78104
rect 519721 78099 519787 78102
rect 523200 78072 524400 78102
rect 116485 78026 116551 78029
rect 116485 78024 119140 78026
rect 116485 77968 116490 78024
rect 116546 77968 119140 78024
rect 116485 77966 119140 77968
rect 116485 77963 116551 77966
rect 520089 76802 520155 76805
rect 518788 76800 520155 76802
rect 518788 76744 520094 76800
rect 520150 76744 520155 76800
rect 518788 76742 520155 76744
rect 520089 76739 520155 76742
rect 519997 76666 520063 76669
rect 523200 76666 524400 76696
rect 519997 76664 524400 76666
rect 519997 76608 520002 76664
rect 520058 76608 524400 76664
rect 519997 76606 524400 76608
rect 519997 76603 520063 76606
rect 523200 76576 524400 76606
rect 110860 75926 119140 75986
rect 519445 75306 519511 75309
rect 518788 75304 519511 75306
rect 518788 75248 519450 75304
rect 519506 75248 519511 75304
rect 518788 75246 519511 75248
rect 519445 75243 519511 75246
rect 519813 75170 519879 75173
rect 523200 75170 524400 75200
rect 519813 75168 524400 75170
rect 519813 75112 519818 75168
rect 519874 75112 524400 75168
rect 519813 75110 524400 75112
rect 519813 75107 519879 75110
rect 523200 75080 524400 75110
rect 116669 74082 116735 74085
rect 116669 74080 119140 74082
rect 116669 74024 116674 74080
rect 116730 74024 119140 74080
rect 116669 74022 119140 74024
rect 116669 74019 116735 74022
rect 519629 73946 519695 73949
rect 518788 73944 519695 73946
rect 518788 73888 519634 73944
rect 519690 73888 519695 73944
rect 518788 73886 519695 73888
rect 519629 73883 519695 73886
rect 519905 73674 519971 73677
rect 523200 73674 524400 73704
rect 519905 73672 524400 73674
rect 519905 73616 519910 73672
rect 519966 73616 524400 73672
rect 519905 73614 524400 73616
rect 519905 73611 519971 73614
rect 523200 73584 524400 73614
rect 519721 72586 519787 72589
rect 518788 72584 519787 72586
rect 518788 72528 519726 72584
rect 519782 72528 519787 72584
rect 518788 72526 519787 72528
rect 519721 72523 519787 72526
rect 116577 72178 116643 72181
rect 116577 72176 119140 72178
rect 116577 72120 116582 72176
rect 116638 72120 119140 72176
rect 116577 72118 119140 72120
rect 116577 72115 116643 72118
rect 520089 72042 520155 72045
rect 523200 72042 524400 72072
rect 520089 72040 524400 72042
rect 520089 71984 520094 72040
rect 520150 71984 524400 72040
rect 520089 71982 524400 71984
rect 520089 71979 520155 71982
rect 523200 71952 524400 71982
rect 519997 71226 520063 71229
rect 518788 71224 520063 71226
rect 518788 71168 520002 71224
rect 520058 71168 520063 71224
rect 518788 71166 520063 71168
rect 519997 71163 520063 71166
rect 520181 70546 520247 70549
rect 523200 70546 524400 70576
rect 520181 70544 524400 70546
rect 520181 70488 520186 70544
rect 520242 70488 524400 70544
rect 520181 70486 524400 70488
rect 520181 70483 520247 70486
rect 523200 70456 524400 70486
rect 116301 70274 116367 70277
rect 116301 70272 119140 70274
rect 116301 70216 116306 70272
rect 116362 70216 119140 70272
rect 116301 70214 119140 70216
rect 116301 70211 116367 70214
rect 519813 69866 519879 69869
rect 518788 69864 519879 69866
rect 518788 69808 519818 69864
rect 519874 69808 519879 69864
rect 518788 69806 519879 69808
rect 519813 69803 519879 69806
rect 519629 69050 519695 69053
rect 523200 69050 524400 69080
rect 519629 69048 524400 69050
rect 519629 68992 519634 69048
rect 519690 68992 524400 69048
rect 519629 68990 524400 68992
rect 519629 68987 519695 68990
rect 523200 68960 524400 68990
rect 519905 68506 519971 68509
rect 518788 68504 519971 68506
rect 518788 68448 519910 68504
rect 519966 68448 519971 68504
rect 518788 68446 519971 68448
rect 519905 68443 519971 68446
rect 116117 68370 116183 68373
rect 116117 68368 119140 68370
rect 116117 68312 116122 68368
rect 116178 68312 119140 68368
rect 116117 68310 119140 68312
rect 116117 68307 116183 68310
rect 520457 67554 520523 67557
rect 523200 67554 524400 67584
rect 520457 67552 524400 67554
rect 520457 67496 520462 67552
rect 520518 67496 524400 67552
rect 520457 67494 524400 67496
rect 520457 67491 520523 67494
rect 523200 67464 524400 67494
rect 520089 67146 520155 67149
rect 518788 67144 520155 67146
rect 518788 67088 520094 67144
rect 520150 67088 520155 67144
rect 518788 67086 520155 67088
rect 520089 67083 520155 67086
rect 116577 66466 116643 66469
rect 116577 66464 119140 66466
rect 116577 66408 116582 66464
rect 116638 66408 119140 66464
rect 116577 66406 119140 66408
rect 116577 66403 116643 66406
rect 520365 66058 520431 66061
rect 523200 66058 524400 66088
rect 520365 66056 524400 66058
rect 520365 66000 520370 66056
rect 520426 66000 524400 66056
rect 520365 65998 524400 66000
rect 520365 65995 520431 65998
rect 523200 65968 524400 65998
rect 520181 65786 520247 65789
rect 518788 65784 520247 65786
rect 518788 65728 520186 65784
rect 520242 65728 520247 65784
rect 518788 65726 520247 65728
rect 520181 65723 520247 65726
rect 114461 64562 114527 64565
rect 110860 64560 114527 64562
rect 110860 64504 114466 64560
rect 114522 64504 114527 64560
rect 110860 64502 114527 64504
rect 114461 64499 114527 64502
rect 116209 64562 116275 64565
rect 520733 64562 520799 64565
rect 523200 64562 524400 64592
rect 116209 64560 119140 64562
rect 116209 64504 116214 64560
rect 116270 64504 119140 64560
rect 116209 64502 119140 64504
rect 520733 64560 524400 64562
rect 520733 64504 520738 64560
rect 520794 64504 524400 64560
rect 520733 64502 524400 64504
rect 116209 64499 116275 64502
rect 520733 64499 520799 64502
rect 523200 64472 524400 64502
rect 519629 64426 519695 64429
rect 518788 64424 519695 64426
rect 518788 64368 519634 64424
rect 519690 64368 519695 64424
rect 518788 64366 519695 64368
rect 519629 64363 519695 64366
rect 520457 63066 520523 63069
rect 518788 63064 520523 63066
rect 518788 63008 520462 63064
rect 520518 63008 520523 63064
rect 518788 63006 520523 63008
rect 520457 63003 520523 63006
rect 521101 62930 521167 62933
rect 523200 62930 524400 62960
rect 521101 62928 524400 62930
rect 521101 62872 521106 62928
rect 521162 62872 524400 62928
rect 521101 62870 524400 62872
rect 521101 62867 521167 62870
rect 523200 62840 524400 62870
rect 116577 62658 116643 62661
rect 116577 62656 119140 62658
rect 116577 62600 116582 62656
rect 116638 62600 119140 62656
rect 116577 62598 119140 62600
rect 116577 62595 116643 62598
rect 520365 61706 520431 61709
rect 518788 61704 520431 61706
rect 518788 61648 520370 61704
rect 520426 61648 520431 61704
rect 518788 61646 520431 61648
rect 520365 61643 520431 61646
rect 521009 61434 521075 61437
rect 523200 61434 524400 61464
rect 521009 61432 524400 61434
rect 521009 61376 521014 61432
rect 521070 61376 524400 61432
rect 521009 61374 524400 61376
rect 521009 61371 521075 61374
rect 523200 61344 524400 61374
rect 116669 60618 116735 60621
rect 116669 60616 119140 60618
rect 116669 60560 116674 60616
rect 116730 60560 119140 60616
rect 116669 60558 119140 60560
rect 116669 60555 116735 60558
rect 520733 60346 520799 60349
rect 518788 60344 520799 60346
rect 518788 60288 520738 60344
rect 520794 60288 520799 60344
rect 518788 60286 520799 60288
rect 520733 60283 520799 60286
rect 520733 59938 520799 59941
rect 523200 59938 524400 59968
rect 520733 59936 524400 59938
rect 520733 59880 520738 59936
rect 520794 59880 524400 59936
rect 520733 59878 524400 59880
rect 520733 59875 520799 59878
rect 523200 59848 524400 59878
rect 521101 58986 521167 58989
rect 518788 58984 521167 58986
rect 518788 58928 521106 58984
rect 521162 58928 521167 58984
rect 518788 58926 521167 58928
rect 521101 58923 521167 58926
rect 116761 58714 116827 58717
rect 116761 58712 119140 58714
rect 116761 58656 116766 58712
rect 116822 58656 119140 58712
rect 116761 58654 119140 58656
rect 116761 58651 116827 58654
rect 521101 58442 521167 58445
rect 523200 58442 524400 58472
rect 521101 58440 524400 58442
rect 521101 58384 521106 58440
rect 521162 58384 524400 58440
rect 521101 58382 524400 58384
rect 521101 58379 521167 58382
rect 523200 58352 524400 58382
rect 521009 57490 521075 57493
rect 518788 57488 521075 57490
rect 518788 57432 521014 57488
rect 521070 57432 521075 57488
rect 518788 57430 521075 57432
rect 521009 57427 521075 57430
rect 520365 56946 520431 56949
rect 523200 56946 524400 56976
rect 520365 56944 524400 56946
rect 520365 56888 520370 56944
rect 520426 56888 524400 56944
rect 520365 56886 524400 56888
rect 520365 56883 520431 56886
rect 523200 56856 524400 56886
rect 116853 56810 116919 56813
rect 116853 56808 119140 56810
rect 116853 56752 116858 56808
rect 116914 56752 119140 56808
rect 116853 56750 119140 56752
rect 116853 56747 116919 56750
rect 520733 56130 520799 56133
rect 518788 56128 520799 56130
rect 518788 56072 520738 56128
rect 520794 56072 520799 56128
rect 518788 56070 520799 56072
rect 520733 56067 520799 56070
rect 520273 55450 520339 55453
rect 523200 55450 524400 55480
rect 520273 55448 524400 55450
rect 520273 55392 520278 55448
rect 520334 55392 524400 55448
rect 520273 55390 524400 55392
rect 520273 55387 520339 55390
rect 523200 55360 524400 55390
rect 116945 54906 117011 54909
rect 116945 54904 119140 54906
rect 116945 54848 116950 54904
rect 117006 54848 119140 54904
rect 116945 54846 119140 54848
rect 116945 54843 117011 54846
rect 521101 54770 521167 54773
rect 518788 54768 521167 54770
rect 518788 54712 521106 54768
rect 521162 54712 521167 54768
rect 518788 54710 521167 54712
rect 521101 54707 521167 54710
rect 519077 53818 519143 53821
rect 523200 53818 524400 53848
rect 519077 53816 524400 53818
rect 519077 53760 519082 53816
rect 519138 53760 524400 53816
rect 519077 53758 524400 53760
rect 519077 53755 519143 53758
rect 523200 53728 524400 53758
rect 520365 53410 520431 53413
rect 518788 53408 520431 53410
rect 518788 53352 520370 53408
rect 520426 53352 520431 53408
rect 518788 53350 520431 53352
rect 520365 53347 520431 53350
rect 114185 53138 114251 53141
rect 110860 53136 114251 53138
rect 110860 53080 114190 53136
rect 114246 53080 114251 53136
rect 110860 53078 114251 53080
rect 114185 53075 114251 53078
rect 117037 53002 117103 53005
rect 117037 53000 119140 53002
rect 117037 52944 117042 53000
rect 117098 52944 119140 53000
rect 117037 52942 119140 52944
rect 117037 52939 117103 52942
rect 519905 52322 519971 52325
rect 523200 52322 524400 52352
rect 519905 52320 524400 52322
rect 519905 52264 519910 52320
rect 519966 52264 524400 52320
rect 519905 52262 524400 52264
rect 519905 52259 519971 52262
rect 523200 52232 524400 52262
rect 520273 52050 520339 52053
rect 518788 52048 520339 52050
rect 518788 51992 520278 52048
rect 520334 51992 520339 52048
rect 518788 51990 520339 51992
rect 520273 51987 520339 51990
rect 117129 51098 117195 51101
rect 117129 51096 119140 51098
rect 117129 51040 117134 51096
rect 117190 51040 119140 51096
rect 117129 51038 119140 51040
rect 117129 51035 117195 51038
rect 519997 50826 520063 50829
rect 523200 50826 524400 50856
rect 519997 50824 524400 50826
rect 519997 50768 520002 50824
rect 520058 50768 524400 50824
rect 519997 50766 524400 50768
rect 519997 50763 520063 50766
rect 523200 50736 524400 50766
rect 519077 50690 519143 50693
rect 518788 50688 519143 50690
rect 518788 50632 519082 50688
rect 519138 50632 519143 50688
rect 518788 50630 519143 50632
rect 519077 50627 519143 50630
rect 519905 49330 519971 49333
rect 518788 49328 519971 49330
rect 518788 49272 519910 49328
rect 519966 49272 519971 49328
rect 518788 49270 519971 49272
rect 519905 49267 519971 49270
rect 520181 49330 520247 49333
rect 523200 49330 524400 49360
rect 520181 49328 524400 49330
rect 520181 49272 520186 49328
rect 520242 49272 524400 49328
rect 520181 49270 524400 49272
rect 520181 49267 520247 49270
rect 523200 49240 524400 49270
rect 117221 49194 117287 49197
rect 117221 49192 119140 49194
rect 117221 49136 117226 49192
rect 117282 49136 119140 49192
rect 117221 49134 119140 49136
rect 117221 49131 117287 49134
rect 519997 47970 520063 47973
rect 518788 47968 520063 47970
rect 518788 47912 520002 47968
rect 520058 47912 520063 47968
rect 518788 47910 520063 47912
rect 519997 47907 520063 47910
rect 519261 47834 519327 47837
rect 523200 47834 524400 47864
rect 519261 47832 524400 47834
rect 519261 47776 519266 47832
rect 519322 47776 524400 47832
rect 519261 47774 524400 47776
rect 519261 47771 519327 47774
rect 523200 47744 524400 47774
rect 116485 47154 116551 47157
rect 116485 47152 119140 47154
rect 116485 47096 116490 47152
rect 116546 47096 119140 47152
rect 116485 47094 119140 47096
rect 116485 47091 116551 47094
rect 520181 46610 520247 46613
rect 518788 46608 520247 46610
rect 518788 46552 520186 46608
rect 520242 46552 520247 46608
rect 518788 46550 520247 46552
rect 520181 46547 520247 46550
rect 519905 46338 519971 46341
rect 523200 46338 524400 46368
rect 519905 46336 524400 46338
rect 519905 46280 519910 46336
rect 519966 46280 524400 46336
rect 519905 46278 524400 46280
rect 519905 46275 519971 46278
rect 523200 46248 524400 46278
rect 116209 45250 116275 45253
rect 519261 45250 519327 45253
rect 116209 45248 119140 45250
rect 116209 45192 116214 45248
rect 116270 45192 119140 45248
rect 116209 45190 119140 45192
rect 518788 45248 519327 45250
rect 518788 45192 519266 45248
rect 519322 45192 519327 45248
rect 518788 45190 519327 45192
rect 116209 45187 116275 45190
rect 519261 45187 519327 45190
rect 519813 44706 519879 44709
rect 523200 44706 524400 44736
rect 519813 44704 524400 44706
rect 519813 44648 519818 44704
rect 519874 44648 524400 44704
rect 519813 44646 524400 44648
rect 519813 44643 519879 44646
rect 523200 44616 524400 44646
rect 519905 43890 519971 43893
rect 518788 43888 519971 43890
rect 518788 43832 519910 43888
rect 519966 43832 519971 43888
rect 518788 43830 519971 43832
rect 519905 43827 519971 43830
rect 116301 43346 116367 43349
rect 116301 43344 119140 43346
rect 116301 43288 116306 43344
rect 116362 43288 119140 43344
rect 116301 43286 119140 43288
rect 116301 43283 116367 43286
rect 520089 43210 520155 43213
rect 523200 43210 524400 43240
rect 520089 43208 524400 43210
rect 520089 43152 520094 43208
rect 520150 43152 524400 43208
rect 520089 43150 524400 43152
rect 520089 43147 520155 43150
rect 523200 43120 524400 43150
rect 519813 42530 519879 42533
rect 518788 42528 519879 42530
rect 518788 42472 519818 42528
rect 519874 42472 519879 42528
rect 518788 42470 519879 42472
rect 519813 42467 519879 42470
rect 114093 41850 114159 41853
rect 110860 41848 114159 41850
rect 110860 41792 114098 41848
rect 114154 41792 114159 41848
rect 110860 41790 114159 41792
rect 114093 41787 114159 41790
rect 520181 41714 520247 41717
rect 523200 41714 524400 41744
rect 520181 41712 524400 41714
rect 520181 41656 520186 41712
rect 520242 41656 524400 41712
rect 520181 41654 524400 41656
rect 520181 41651 520247 41654
rect 523200 41624 524400 41654
rect 116117 41442 116183 41445
rect 116117 41440 119140 41442
rect 116117 41384 116122 41440
rect 116178 41384 119140 41440
rect 116117 41382 119140 41384
rect 116117 41379 116183 41382
rect 520089 41170 520155 41173
rect 518788 41168 520155 41170
rect 518788 41112 520094 41168
rect 520150 41112 520155 41168
rect 518788 41110 520155 41112
rect 520089 41107 520155 41110
rect 519813 40218 519879 40221
rect 523200 40218 524400 40248
rect 519813 40216 524400 40218
rect 519813 40160 519818 40216
rect 519874 40160 524400 40216
rect 519813 40158 524400 40160
rect 519813 40155 519879 40158
rect 523200 40128 524400 40158
rect 520181 39810 520247 39813
rect 518788 39808 520247 39810
rect 518788 39752 520186 39808
rect 520242 39752 520247 39808
rect 518788 39750 520247 39752
rect 520181 39747 520247 39750
rect 116393 39538 116459 39541
rect 116393 39536 119140 39538
rect 116393 39480 116398 39536
rect 116454 39480 119140 39536
rect 116393 39478 119140 39480
rect 116393 39475 116459 39478
rect 520181 38722 520247 38725
rect 523200 38722 524400 38752
rect 520181 38720 524400 38722
rect 520181 38664 520186 38720
rect 520242 38664 524400 38720
rect 520181 38662 524400 38664
rect 520181 38659 520247 38662
rect 523200 38632 524400 38662
rect 519813 38314 519879 38317
rect 518788 38312 519879 38314
rect 518788 38256 519818 38312
rect 519874 38256 519879 38312
rect 518788 38254 519879 38256
rect 519813 38251 519879 38254
rect 116209 37634 116275 37637
rect 116209 37632 119140 37634
rect 116209 37576 116214 37632
rect 116270 37576 119140 37632
rect 116209 37574 119140 37576
rect 116209 37571 116275 37574
rect 521101 37226 521167 37229
rect 523200 37226 524400 37256
rect 521101 37224 524400 37226
rect 521101 37168 521106 37224
rect 521162 37168 524400 37224
rect 521101 37166 524400 37168
rect 521101 37163 521167 37166
rect 523200 37136 524400 37166
rect 520181 36954 520247 36957
rect 518788 36952 520247 36954
rect 518788 36896 520186 36952
rect 520242 36896 520247 36952
rect 518788 36894 520247 36896
rect 520181 36891 520247 36894
rect 521101 36002 521167 36005
rect 518758 36000 521167 36002
rect 518758 35944 521106 36000
rect 521162 35944 521167 36000
rect 518758 35942 521167 35944
rect 116117 35730 116183 35733
rect 116117 35728 119140 35730
rect 116117 35672 116122 35728
rect 116178 35672 119140 35728
rect 116117 35670 119140 35672
rect 116117 35667 116183 35670
rect 518758 35564 518818 35942
rect 521101 35939 521167 35942
rect 520917 35594 520983 35597
rect 523200 35594 524400 35624
rect 520917 35592 524400 35594
rect 520917 35536 520922 35592
rect 520978 35536 524400 35592
rect 520917 35534 524400 35536
rect 520917 35531 520983 35534
rect 523200 35504 524400 35534
rect 520917 34642 520983 34645
rect 518758 34640 520983 34642
rect 518758 34584 520922 34640
rect 520978 34584 520983 34640
rect 518758 34582 520983 34584
rect 518758 34204 518818 34582
rect 520917 34579 520983 34582
rect 520825 34098 520891 34101
rect 523200 34098 524400 34128
rect 520825 34096 524400 34098
rect 520825 34040 520830 34096
rect 520886 34040 524400 34096
rect 520825 34038 524400 34040
rect 520825 34035 520891 34038
rect 523200 34008 524400 34038
rect 116117 33826 116183 33829
rect 116117 33824 119140 33826
rect 116117 33768 116122 33824
rect 116178 33768 119140 33824
rect 116117 33766 119140 33768
rect 116117 33763 116183 33766
rect 520825 33282 520891 33285
rect 518758 33280 520891 33282
rect 518758 33224 520830 33280
rect 520886 33224 520891 33280
rect 518758 33222 520891 33224
rect 518758 32844 518818 33222
rect 520825 33219 520891 33222
rect 521101 32602 521167 32605
rect 523200 32602 524400 32632
rect 521101 32600 524400 32602
rect 521101 32544 521106 32600
rect 521162 32544 524400 32600
rect 521101 32542 524400 32544
rect 521101 32539 521167 32542
rect 523200 32512 524400 32542
rect 116117 31786 116183 31789
rect 521101 31786 521167 31789
rect 116117 31784 119140 31786
rect 116117 31728 116122 31784
rect 116178 31728 119140 31784
rect 116117 31726 119140 31728
rect 518758 31784 521167 31786
rect 518758 31728 521106 31784
rect 521162 31728 521167 31784
rect 518758 31726 521167 31728
rect 116117 31723 116183 31726
rect 518758 31484 518818 31726
rect 521101 31723 521167 31726
rect 521101 31106 521167 31109
rect 523200 31106 524400 31136
rect 521101 31104 524400 31106
rect 521101 31048 521106 31104
rect 521162 31048 524400 31104
rect 521101 31046 524400 31048
rect 521101 31043 521167 31046
rect 523200 31016 524400 31046
rect 114001 30426 114067 30429
rect 521101 30426 521167 30429
rect 110860 30424 114067 30426
rect 110860 30368 114006 30424
rect 114062 30368 114067 30424
rect 110860 30366 114067 30368
rect 114001 30363 114067 30366
rect 518758 30424 521167 30426
rect 518758 30368 521106 30424
rect 521162 30368 521167 30424
rect 518758 30366 521167 30368
rect 518758 30124 518818 30366
rect 521101 30363 521167 30366
rect 116117 29882 116183 29885
rect 116117 29880 119140 29882
rect 116117 29824 116122 29880
rect 116178 29824 119140 29880
rect 116117 29822 119140 29824
rect 116117 29819 116183 29822
rect 521101 29610 521167 29613
rect 523200 29610 524400 29640
rect 521101 29608 524400 29610
rect 521101 29552 521106 29608
rect 521162 29552 524400 29608
rect 521101 29550 524400 29552
rect 521101 29547 521167 29550
rect 523200 29520 524400 29550
rect 521101 28794 521167 28797
rect 518788 28792 521167 28794
rect 518788 28736 521106 28792
rect 521162 28736 521167 28792
rect 518788 28734 521167 28736
rect 521101 28731 521167 28734
rect 523200 28114 524400 28144
rect 518850 28054 524400 28114
rect 116117 27978 116183 27981
rect 518850 27978 518910 28054
rect 523200 28024 524400 28054
rect 116117 27976 119140 27978
rect 116117 27920 116122 27976
rect 116178 27920 119140 27976
rect 116117 27918 119140 27920
rect 518758 27918 518910 27978
rect 116117 27915 116183 27918
rect 518758 27404 518818 27918
rect 523200 26482 524400 26512
rect 518850 26422 524400 26482
rect 518850 26346 518910 26422
rect 523200 26392 524400 26422
rect 518758 26286 518910 26346
rect 116117 26074 116183 26077
rect 116117 26072 119140 26074
rect 116117 26016 116122 26072
rect 116178 26016 119140 26072
rect 518758 26044 518818 26286
rect 116117 26014 119140 26016
rect 116117 26011 116183 26014
rect 523200 24986 524400 25016
rect 518758 24926 524400 24986
rect 518758 24684 518818 24926
rect 523200 24896 524400 24926
rect 116117 24170 116183 24173
rect 116117 24168 119140 24170
rect 116117 24112 116122 24168
rect 116178 24112 119140 24168
rect 116117 24110 119140 24112
rect 116117 24107 116183 24110
rect 523200 23490 524400 23520
rect 518758 23430 524400 23490
rect 518758 23324 518818 23430
rect 523200 23400 524400 23430
rect 116025 22266 116091 22269
rect 116025 22264 119140 22266
rect 116025 22208 116030 22264
rect 116086 22208 119140 22264
rect 116025 22206 119140 22208
rect 116025 22203 116091 22206
rect 523200 21994 524400 22024
rect 518788 21934 524400 21994
rect 523200 21904 524400 21934
rect 521101 20498 521167 20501
rect 523200 20498 524400 20528
rect 521101 20496 524400 20498
rect 116209 20362 116275 20365
rect 116209 20360 119140 20362
rect 116209 20304 116214 20360
rect 116270 20304 119140 20360
rect 116209 20302 119140 20304
rect 116209 20299 116275 20302
rect 518758 19818 518818 20468
rect 521101 20440 521106 20496
rect 521162 20440 524400 20496
rect 521101 20438 524400 20440
rect 521101 20435 521167 20438
rect 523200 20408 524400 20438
rect 521101 19818 521167 19821
rect 518758 19816 521167 19818
rect 518758 19760 521106 19816
rect 521162 19760 521167 19816
rect 518758 19758 521167 19760
rect 521101 19755 521167 19758
rect 113909 19002 113975 19005
rect 110860 19000 113975 19002
rect 110860 18944 113914 19000
rect 113970 18944 113975 19000
rect 110860 18942 113975 18944
rect 113909 18939 113975 18942
rect 116117 18458 116183 18461
rect 518758 18458 518818 19108
rect 523200 19002 524400 19032
rect 521150 18942 524400 19002
rect 521150 18458 521210 18942
rect 523200 18912 524400 18942
rect 116117 18456 119140 18458
rect 116117 18400 116122 18456
rect 116178 18400 119140 18456
rect 116117 18398 119140 18400
rect 518758 18398 521210 18458
rect 116117 18395 116183 18398
rect 518758 17098 518818 17748
rect 523200 17370 524400 17400
rect 521150 17310 524400 17370
rect 521150 17098 521210 17310
rect 523200 17280 524400 17310
rect 518758 17038 521210 17098
rect 116209 16418 116275 16421
rect 116209 16416 119140 16418
rect 116209 16360 116214 16416
rect 116270 16360 119140 16416
rect 116209 16358 119140 16360
rect 116209 16355 116275 16358
rect 518758 15738 518818 16388
rect 523200 15874 524400 15904
rect 521104 15814 524400 15874
rect 521104 15738 521164 15814
rect 523200 15784 524400 15814
rect 518758 15678 521164 15738
rect 521101 15058 521167 15061
rect 518788 15056 521167 15058
rect 518788 15000 521106 15056
rect 521162 15000 521167 15056
rect 518788 14998 521167 15000
rect 521101 14995 521167 14998
rect 115933 14514 115999 14517
rect 115933 14512 119140 14514
rect 115933 14456 115938 14512
rect 115994 14456 119140 14512
rect 115933 14454 119140 14456
rect 115933 14451 115999 14454
rect 521101 14378 521167 14381
rect 523200 14378 524400 14408
rect 521101 14376 524400 14378
rect 521101 14320 521106 14376
rect 521162 14320 524400 14376
rect 521101 14318 524400 14320
rect 521101 14315 521167 14318
rect 523200 14288 524400 14318
rect 521101 13698 521167 13701
rect 518788 13696 521167 13698
rect 518788 13640 521106 13696
rect 521162 13640 521167 13696
rect 518788 13638 521167 13640
rect 521101 13635 521167 13638
rect 521101 12882 521167 12885
rect 523200 12882 524400 12912
rect 521101 12880 524400 12882
rect 521101 12824 521106 12880
rect 521162 12824 524400 12880
rect 521101 12822 524400 12824
rect 521101 12819 521167 12822
rect 523200 12792 524400 12822
rect 116526 12548 116532 12612
rect 116596 12610 116602 12612
rect 116596 12550 119140 12610
rect 116596 12548 116602 12550
rect 519629 12338 519695 12341
rect 518788 12336 519695 12338
rect 518788 12280 519634 12336
rect 519690 12280 519695 12336
rect 518788 12278 519695 12280
rect 519629 12275 519695 12278
rect 519629 11386 519695 11389
rect 523200 11386 524400 11416
rect 519629 11384 524400 11386
rect 519629 11328 519634 11384
rect 519690 11328 524400 11384
rect 519629 11326 524400 11328
rect 519629 11323 519695 11326
rect 523200 11296 524400 11326
rect 521101 10978 521167 10981
rect 518788 10976 521167 10978
rect 518788 10920 521106 10976
rect 521162 10920 521167 10976
rect 518788 10918 521167 10920
rect 521101 10915 521167 10918
rect 116710 10644 116716 10708
rect 116780 10706 116786 10708
rect 116780 10646 119140 10706
rect 116780 10644 116786 10646
rect 521101 9890 521167 9893
rect 523200 9890 524400 9920
rect 521101 9888 524400 9890
rect 521101 9832 521106 9888
rect 521162 9832 524400 9888
rect 521101 9830 524400 9832
rect 521101 9827 521167 9830
rect 523200 9800 524400 9830
rect 521101 9618 521167 9621
rect 518788 9616 521167 9618
rect 518788 9560 521106 9616
rect 521162 9560 521167 9616
rect 518788 9558 521167 9560
rect 521101 9555 521167 9558
rect 117262 8740 117268 8804
rect 117332 8802 117338 8804
rect 117332 8742 119140 8802
rect 117332 8740 117338 8742
rect 520365 8258 520431 8261
rect 518788 8256 520431 8258
rect 518788 8200 520370 8256
rect 520426 8200 520431 8256
rect 518788 8198 520431 8200
rect 520365 8195 520431 8198
rect 521101 8258 521167 8261
rect 523200 8258 524400 8288
rect 521101 8256 524400 8258
rect 521101 8200 521106 8256
rect 521162 8200 524400 8256
rect 521101 8198 524400 8200
rect 521101 8195 521167 8198
rect 523200 8168 524400 8198
rect 113817 7714 113883 7717
rect 110860 7712 113883 7714
rect 110860 7656 113822 7712
rect 113878 7656 113883 7712
rect 110860 7654 113883 7656
rect 113817 7651 113883 7654
rect 116158 6836 116164 6900
rect 116228 6898 116234 6900
rect 521101 6898 521167 6901
rect 116228 6838 119140 6898
rect 518788 6896 521167 6898
rect 518788 6840 521106 6896
rect 521162 6840 521167 6896
rect 518788 6838 521167 6840
rect 116228 6836 116234 6838
rect 521101 6835 521167 6838
rect 520365 6762 520431 6765
rect 523200 6762 524400 6792
rect 520365 6760 524400 6762
rect 520365 6704 520370 6760
rect 520426 6704 524400 6760
rect 520365 6702 524400 6704
rect 520365 6699 520431 6702
rect 523200 6672 524400 6702
rect 521009 5538 521075 5541
rect 518788 5536 521075 5538
rect 518788 5480 521014 5536
rect 521070 5480 521075 5536
rect 518788 5478 521075 5480
rect 521009 5475 521075 5478
rect 521101 5266 521167 5269
rect 523200 5266 524400 5296
rect 521101 5264 524400 5266
rect 521101 5208 521106 5264
rect 521162 5208 524400 5264
rect 521101 5206 524400 5208
rect 521101 5203 521167 5206
rect 523200 5176 524400 5206
rect 116117 4994 116183 4997
rect 116117 4992 119140 4994
rect 116117 4936 116122 4992
rect 116178 4936 119140 4992
rect 116117 4934 119140 4936
rect 116117 4931 116183 4934
rect 521101 4178 521167 4181
rect 518788 4176 521167 4178
rect 518788 4120 521106 4176
rect 521162 4120 521167 4176
rect 518788 4118 521167 4120
rect 521101 4115 521167 4118
rect 521009 3770 521075 3773
rect 523200 3770 524400 3800
rect 521009 3768 524400 3770
rect 521009 3712 521014 3768
rect 521070 3712 524400 3768
rect 521009 3710 524400 3712
rect 521009 3707 521075 3710
rect 523200 3680 524400 3710
rect 116117 3090 116183 3093
rect 116117 3088 119140 3090
rect 116117 3032 116122 3088
rect 116178 3032 119140 3088
rect 116117 3030 119140 3032
rect 116117 3027 116183 3030
rect 519997 2818 520063 2821
rect 518788 2816 520063 2818
rect 518788 2760 520002 2816
rect 520058 2760 520063 2816
rect 518788 2758 520063 2760
rect 519997 2755 520063 2758
rect 39113 2682 39179 2685
rect 53465 2682 53531 2685
rect 81249 2682 81315 2685
rect 39113 2680 53531 2682
rect 39113 2624 39118 2680
rect 39174 2624 53470 2680
rect 53526 2624 53531 2680
rect 39113 2622 53531 2624
rect 39113 2619 39179 2622
rect 53465 2619 53531 2622
rect 53790 2680 81315 2682
rect 53790 2624 81254 2680
rect 81310 2624 81315 2680
rect 53790 2622 81315 2624
rect 42793 2546 42859 2549
rect 50889 2546 50955 2549
rect 42793 2544 50955 2546
rect 42793 2488 42798 2544
rect 42854 2488 50894 2544
rect 50950 2488 50955 2544
rect 42793 2486 50955 2488
rect 42793 2483 42859 2486
rect 50889 2483 50955 2486
rect 49141 2410 49207 2413
rect 53790 2410 53850 2622
rect 81249 2619 81315 2622
rect 106089 2682 106155 2685
rect 109585 2682 109651 2685
rect 106089 2680 109651 2682
rect 106089 2624 106094 2680
rect 106150 2624 109590 2680
rect 109646 2624 109651 2680
rect 106089 2622 109651 2624
rect 106089 2619 106155 2622
rect 109585 2619 109651 2622
rect 58617 2546 58683 2549
rect 82261 2546 82327 2549
rect 58617 2544 82327 2546
rect 58617 2488 58622 2544
rect 58678 2488 82266 2544
rect 82322 2488 82327 2544
rect 58617 2486 82327 2488
rect 58617 2483 58683 2486
rect 82261 2483 82327 2486
rect 49141 2408 53850 2410
rect 49141 2352 49146 2408
rect 49202 2352 53850 2408
rect 49141 2350 53850 2352
rect 62389 2410 62455 2413
rect 63033 2410 63099 2413
rect 62389 2408 63099 2410
rect 62389 2352 62394 2408
rect 62450 2352 63038 2408
rect 63094 2352 63099 2408
rect 62389 2350 63099 2352
rect 49141 2347 49207 2350
rect 62389 2347 62455 2350
rect 63033 2347 63099 2350
rect 78029 2410 78095 2413
rect 79777 2410 79843 2413
rect 78029 2408 79843 2410
rect 78029 2352 78034 2408
rect 78090 2352 79782 2408
rect 79838 2352 79843 2408
rect 78029 2350 79843 2352
rect 78029 2347 78095 2350
rect 79777 2347 79843 2350
rect 78121 2274 78187 2277
rect 79685 2274 79751 2277
rect 78121 2272 79751 2274
rect 78121 2216 78126 2272
rect 78182 2216 79690 2272
rect 79746 2216 79751 2272
rect 78121 2214 79751 2216
rect 78121 2211 78187 2214
rect 79685 2211 79751 2214
rect 521101 2274 521167 2277
rect 523200 2274 524400 2304
rect 521101 2272 524400 2274
rect 521101 2216 521106 2272
rect 521162 2216 524400 2272
rect 521101 2214 524400 2216
rect 521101 2211 521167 2214
rect 523200 2184 524400 2214
rect 19333 1866 19399 1869
rect 116526 1866 116532 1868
rect 19333 1864 116532 1866
rect 19333 1808 19338 1864
rect 19394 1808 116532 1864
rect 19333 1806 116532 1808
rect 19333 1803 19399 1806
rect 116526 1804 116532 1806
rect 116596 1804 116602 1868
rect 15929 1730 15995 1733
rect 116710 1730 116716 1732
rect 15929 1728 116716 1730
rect 15929 1672 15934 1728
rect 15990 1672 116716 1728
rect 15929 1670 116716 1672
rect 15929 1667 15995 1670
rect 116710 1668 116716 1670
rect 116780 1668 116786 1732
rect 12617 1594 12683 1597
rect 117262 1594 117268 1596
rect 12617 1592 117268 1594
rect 12617 1536 12622 1592
rect 12678 1536 117268 1592
rect 12617 1534 117268 1536
rect 12617 1531 12683 1534
rect 117262 1532 117268 1534
rect 117332 1532 117338 1596
rect 229277 1594 229343 1597
rect 293585 1594 293651 1597
rect 229277 1592 293651 1594
rect 229277 1536 229282 1592
rect 229338 1536 293590 1592
rect 293646 1536 293651 1592
rect 229277 1534 293651 1536
rect 229277 1531 229343 1534
rect 293585 1531 293651 1534
rect 9305 1458 9371 1461
rect 116158 1458 116164 1460
rect 9305 1456 116164 1458
rect 9305 1400 9310 1456
rect 9366 1400 116164 1456
rect 9305 1398 116164 1400
rect 9305 1395 9371 1398
rect 116158 1396 116164 1398
rect 116228 1396 116234 1460
rect 163773 1458 163839 1461
rect 243629 1458 243695 1461
rect 163773 1456 243695 1458
rect 163773 1400 163778 1456
rect 163834 1400 243634 1456
rect 243690 1400 243695 1456
rect 163773 1398 243695 1400
rect 163773 1395 163839 1398
rect 243629 1395 243695 1398
rect 360285 1458 360351 1461
rect 393589 1458 393655 1461
rect 360285 1456 393655 1458
rect 360285 1400 360290 1456
rect 360346 1400 393594 1456
rect 393650 1400 393655 1456
rect 360285 1398 393655 1400
rect 360285 1395 360351 1398
rect 393589 1395 393655 1398
rect 519997 778 520063 781
rect 523200 778 524400 808
rect 519997 776 524400 778
rect 519997 720 520002 776
rect 520058 720 524400 776
rect 519997 718 524400 720
rect 519997 715 520063 718
rect 523200 688 524400 718
<< via3 >>
rect 116532 12548 116596 12612
rect 116716 10644 116780 10708
rect 117268 8740 117332 8804
rect 116164 6836 116228 6900
rect 116532 1804 116596 1868
rect 116716 1668 116780 1732
rect 117268 1532 117332 1596
rect 116164 1396 116228 1460
<< metal4 >>
rect 1664 144454 1984 144496
rect 1664 144218 1706 144454
rect 1942 144218 1984 144454
rect 1664 144134 1984 144218
rect 1664 143898 1706 144134
rect 1942 143898 1984 144134
rect 1664 143856 1984 143898
rect 109956 144454 110276 144496
rect 109956 144218 109998 144454
rect 110234 144218 110276 144454
rect 109956 144134 110276 144218
rect 109956 143898 109998 144134
rect 110234 143898 110276 144134
rect 109956 143856 110276 143898
rect 119664 144454 119984 144496
rect 119664 144218 119706 144454
rect 119942 144218 119984 144454
rect 119664 144134 119984 144218
rect 119664 143898 119706 144134
rect 119942 143898 119984 144134
rect 119664 143856 119984 143898
rect 517940 144454 518260 144496
rect 517940 144218 517982 144454
rect 518218 144218 518260 144454
rect 517940 144134 518260 144218
rect 517940 143898 517982 144134
rect 518218 143898 518260 144134
rect 517940 143856 518260 143898
rect 1096 131454 1332 131496
rect 1096 131134 1332 131218
rect 1096 130856 1332 130898
rect 110616 131454 110936 131496
rect 110616 131218 110658 131454
rect 110894 131218 110936 131454
rect 110616 131134 110936 131218
rect 110616 130898 110658 131134
rect 110894 130898 110936 131134
rect 110616 130856 110936 130898
rect 119004 131454 119324 131496
rect 119004 131218 119046 131454
rect 119282 131218 119324 131454
rect 119004 131134 119324 131218
rect 119004 130898 119046 131134
rect 119282 130898 119324 131134
rect 119004 130856 119324 130898
rect 518600 131454 518920 131496
rect 518600 131218 518642 131454
rect 518878 131218 518920 131454
rect 518600 131134 518920 131218
rect 518600 130898 518642 131134
rect 518878 130898 518920 131134
rect 518600 130856 518920 130898
rect 1664 118454 1984 118496
rect 1664 118218 1706 118454
rect 1942 118218 1984 118454
rect 1664 118134 1984 118218
rect 1664 117898 1706 118134
rect 1942 117898 1984 118134
rect 1664 117856 1984 117898
rect 109956 118454 110276 118496
rect 109956 118218 109998 118454
rect 110234 118218 110276 118454
rect 109956 118134 110276 118218
rect 109956 117898 109998 118134
rect 110234 117898 110276 118134
rect 109956 117856 110276 117898
rect 119664 118454 119984 118496
rect 119664 118218 119706 118454
rect 119942 118218 119984 118454
rect 119664 118134 119984 118218
rect 119664 117898 119706 118134
rect 119942 117898 119984 118134
rect 119664 117856 119984 117898
rect 517940 118454 518260 118496
rect 517940 118218 517982 118454
rect 518218 118218 518260 118454
rect 517940 118134 518260 118218
rect 517940 117898 517982 118134
rect 518218 117898 518260 118134
rect 517940 117856 518260 117898
rect 1096 105454 1332 105496
rect 1096 105134 1332 105218
rect 1096 104856 1332 104898
rect 110616 105454 110936 105496
rect 110616 105218 110658 105454
rect 110894 105218 110936 105454
rect 110616 105134 110936 105218
rect 110616 104898 110658 105134
rect 110894 104898 110936 105134
rect 110616 104856 110936 104898
rect 119004 105454 119324 105496
rect 119004 105218 119046 105454
rect 119282 105218 119324 105454
rect 119004 105134 119324 105218
rect 119004 104898 119046 105134
rect 119282 104898 119324 105134
rect 119004 104856 119324 104898
rect 518600 105454 518920 105496
rect 518600 105218 518642 105454
rect 518878 105218 518920 105454
rect 518600 105134 518920 105218
rect 518600 104898 518642 105134
rect 518878 104898 518920 105134
rect 518600 104856 518920 104898
rect 1664 92454 1984 92496
rect 1664 92218 1706 92454
rect 1942 92218 1984 92454
rect 1664 92134 1984 92218
rect 1664 91898 1706 92134
rect 1942 91898 1984 92134
rect 1664 91856 1984 91898
rect 109956 92454 110276 92496
rect 109956 92218 109998 92454
rect 110234 92218 110276 92454
rect 109956 92134 110276 92218
rect 109956 91898 109998 92134
rect 110234 91898 110276 92134
rect 109956 91856 110276 91898
rect 119664 92454 119984 92496
rect 119664 92218 119706 92454
rect 119942 92218 119984 92454
rect 119664 92134 119984 92218
rect 119664 91898 119706 92134
rect 119942 91898 119984 92134
rect 119664 91856 119984 91898
rect 517940 92454 518260 92496
rect 517940 92218 517982 92454
rect 518218 92218 518260 92454
rect 517940 92134 518260 92218
rect 517940 91898 517982 92134
rect 518218 91898 518260 92134
rect 517940 91856 518260 91898
rect 1096 79454 1332 79496
rect 1096 79134 1332 79218
rect 1096 78856 1332 78898
rect 110616 79454 110936 79496
rect 110616 79218 110658 79454
rect 110894 79218 110936 79454
rect 110616 79134 110936 79218
rect 110616 78898 110658 79134
rect 110894 78898 110936 79134
rect 110616 78856 110936 78898
rect 119004 79454 119324 79496
rect 119004 79218 119046 79454
rect 119282 79218 119324 79454
rect 119004 79134 119324 79218
rect 119004 78898 119046 79134
rect 119282 78898 119324 79134
rect 119004 78856 119324 78898
rect 518600 79454 518920 79496
rect 518600 79218 518642 79454
rect 518878 79218 518920 79454
rect 518600 79134 518920 79218
rect 518600 78898 518642 79134
rect 518878 78898 518920 79134
rect 518600 78856 518920 78898
rect 1664 66454 1984 66496
rect 1664 66218 1706 66454
rect 1942 66218 1984 66454
rect 1664 66134 1984 66218
rect 1664 65898 1706 66134
rect 1942 65898 1984 66134
rect 1664 65856 1984 65898
rect 109956 66454 110276 66496
rect 109956 66218 109998 66454
rect 110234 66218 110276 66454
rect 109956 66134 110276 66218
rect 109956 65898 109998 66134
rect 110234 65898 110276 66134
rect 109956 65856 110276 65898
rect 119664 66454 119984 66496
rect 119664 66218 119706 66454
rect 119942 66218 119984 66454
rect 119664 66134 119984 66218
rect 119664 65898 119706 66134
rect 119942 65898 119984 66134
rect 119664 65856 119984 65898
rect 517940 66454 518260 66496
rect 517940 66218 517982 66454
rect 518218 66218 518260 66454
rect 517940 66134 518260 66218
rect 517940 65898 517982 66134
rect 518218 65898 518260 66134
rect 517940 65856 518260 65898
rect 1096 53454 1332 53496
rect 1096 53134 1332 53218
rect 1096 52856 1332 52898
rect 110616 53454 110936 53496
rect 110616 53218 110658 53454
rect 110894 53218 110936 53454
rect 110616 53134 110936 53218
rect 110616 52898 110658 53134
rect 110894 52898 110936 53134
rect 110616 52856 110936 52898
rect 119004 53454 119324 53496
rect 119004 53218 119046 53454
rect 119282 53218 119324 53454
rect 119004 53134 119324 53218
rect 119004 52898 119046 53134
rect 119282 52898 119324 53134
rect 119004 52856 119324 52898
rect 518600 53454 518920 53496
rect 518600 53218 518642 53454
rect 518878 53218 518920 53454
rect 518600 53134 518920 53218
rect 518600 52898 518642 53134
rect 518878 52898 518920 53134
rect 518600 52856 518920 52898
rect 1664 40454 1984 40496
rect 1664 40218 1706 40454
rect 1942 40218 1984 40454
rect 1664 40134 1984 40218
rect 1664 39898 1706 40134
rect 1942 39898 1984 40134
rect 1664 39856 1984 39898
rect 109956 40454 110276 40496
rect 109956 40218 109998 40454
rect 110234 40218 110276 40454
rect 109956 40134 110276 40218
rect 109956 39898 109998 40134
rect 110234 39898 110276 40134
rect 109956 39856 110276 39898
rect 119664 40454 119984 40496
rect 119664 40218 119706 40454
rect 119942 40218 119984 40454
rect 119664 40134 119984 40218
rect 119664 39898 119706 40134
rect 119942 39898 119984 40134
rect 119664 39856 119984 39898
rect 517940 40454 518260 40496
rect 517940 40218 517982 40454
rect 518218 40218 518260 40454
rect 517940 40134 518260 40218
rect 517940 39898 517982 40134
rect 518218 39898 518260 40134
rect 517940 39856 518260 39898
rect 1096 27454 1332 27496
rect 1096 27134 1332 27218
rect 1096 26856 1332 26898
rect 110616 27454 110936 27496
rect 110616 27218 110658 27454
rect 110894 27218 110936 27454
rect 110616 27134 110936 27218
rect 110616 26898 110658 27134
rect 110894 26898 110936 27134
rect 110616 26856 110936 26898
rect 119004 27454 119324 27496
rect 119004 27218 119046 27454
rect 119282 27218 119324 27454
rect 119004 27134 119324 27218
rect 119004 26898 119046 27134
rect 119282 26898 119324 27134
rect 119004 26856 119324 26898
rect 518600 27454 518920 27496
rect 518600 27218 518642 27454
rect 518878 27218 518920 27454
rect 518600 27134 518920 27218
rect 518600 26898 518642 27134
rect 518878 26898 518920 27134
rect 518600 26856 518920 26898
rect 1664 14454 1984 14496
rect 1664 14218 1706 14454
rect 1942 14218 1984 14454
rect 1664 14134 1984 14218
rect 1664 13898 1706 14134
rect 1942 13898 1984 14134
rect 1664 13856 1984 13898
rect 109956 14454 110276 14496
rect 109956 14218 109998 14454
rect 110234 14218 110276 14454
rect 109956 14134 110276 14218
rect 109956 13898 109998 14134
rect 110234 13898 110276 14134
rect 109956 13856 110276 13898
rect 119664 14454 119984 14496
rect 119664 14218 119706 14454
rect 119942 14218 119984 14454
rect 119664 14134 119984 14218
rect 119664 13898 119706 14134
rect 119942 13898 119984 14134
rect 119664 13856 119984 13898
rect 517940 14454 518260 14496
rect 517940 14218 517982 14454
rect 518218 14218 518260 14454
rect 517940 14134 518260 14218
rect 517940 13898 517982 14134
rect 518218 13898 518260 14134
rect 517940 13856 518260 13898
rect 116531 12612 116597 12613
rect 116531 12548 116532 12612
rect 116596 12548 116597 12612
rect 116531 12547 116597 12548
rect 116163 6900 116229 6901
rect 116163 6836 116164 6900
rect 116228 6836 116229 6900
rect 116163 6835 116229 6836
rect 116166 1461 116226 6835
rect 116534 1869 116594 12547
rect 116715 10708 116781 10709
rect 116715 10644 116716 10708
rect 116780 10644 116781 10708
rect 116715 10643 116781 10644
rect 116531 1868 116597 1869
rect 116531 1804 116532 1868
rect 116596 1804 116597 1868
rect 116531 1803 116597 1804
rect 116718 1733 116778 10643
rect 117267 8804 117333 8805
rect 117267 8740 117268 8804
rect 117332 8740 117333 8804
rect 117267 8739 117333 8740
rect 116715 1732 116781 1733
rect 116715 1668 116716 1732
rect 116780 1668 116781 1732
rect 116715 1667 116781 1668
rect 117270 1597 117330 8739
rect 117267 1596 117333 1597
rect 117267 1532 117268 1596
rect 117332 1532 117333 1596
rect 117267 1531 117333 1532
rect 116163 1460 116229 1461
rect 116163 1396 116164 1460
rect 116228 1396 116229 1460
rect 116163 1395 116229 1396
<< via4 >>
rect 1706 144218 1942 144454
rect 1706 143898 1942 144134
rect 109998 144218 110234 144454
rect 109998 143898 110234 144134
rect 119706 144218 119942 144454
rect 119706 143898 119942 144134
rect 517982 144218 518218 144454
rect 517982 143898 518218 144134
rect 1096 131218 1332 131454
rect 1096 130898 1332 131134
rect 110658 131218 110894 131454
rect 110658 130898 110894 131134
rect 119046 131218 119282 131454
rect 119046 130898 119282 131134
rect 518642 131218 518878 131454
rect 518642 130898 518878 131134
rect 1706 118218 1942 118454
rect 1706 117898 1942 118134
rect 109998 118218 110234 118454
rect 109998 117898 110234 118134
rect 119706 118218 119942 118454
rect 119706 117898 119942 118134
rect 517982 118218 518218 118454
rect 517982 117898 518218 118134
rect 1096 105218 1332 105454
rect 1096 104898 1332 105134
rect 110658 105218 110894 105454
rect 110658 104898 110894 105134
rect 119046 105218 119282 105454
rect 119046 104898 119282 105134
rect 518642 105218 518878 105454
rect 518642 104898 518878 105134
rect 1706 92218 1942 92454
rect 1706 91898 1942 92134
rect 109998 92218 110234 92454
rect 109998 91898 110234 92134
rect 119706 92218 119942 92454
rect 119706 91898 119942 92134
rect 517982 92218 518218 92454
rect 517982 91898 518218 92134
rect 1096 79218 1332 79454
rect 1096 78898 1332 79134
rect 110658 79218 110894 79454
rect 110658 78898 110894 79134
rect 119046 79218 119282 79454
rect 119046 78898 119282 79134
rect 518642 79218 518878 79454
rect 518642 78898 518878 79134
rect 1706 66218 1942 66454
rect 1706 65898 1942 66134
rect 109998 66218 110234 66454
rect 109998 65898 110234 66134
rect 119706 66218 119942 66454
rect 119706 65898 119942 66134
rect 517982 66218 518218 66454
rect 517982 65898 518218 66134
rect 1096 53218 1332 53454
rect 1096 52898 1332 53134
rect 110658 53218 110894 53454
rect 110658 52898 110894 53134
rect 119046 53218 119282 53454
rect 119046 52898 119282 53134
rect 518642 53218 518878 53454
rect 518642 52898 518878 53134
rect 1706 40218 1942 40454
rect 1706 39898 1942 40134
rect 109998 40218 110234 40454
rect 109998 39898 110234 40134
rect 119706 40218 119942 40454
rect 119706 39898 119942 40134
rect 517982 40218 518218 40454
rect 517982 39898 518218 40134
rect 1096 27218 1332 27454
rect 1096 26898 1332 27134
rect 110658 27218 110894 27454
rect 110658 26898 110894 27134
rect 119046 27218 119282 27454
rect 119046 26898 119282 27134
rect 518642 27218 518878 27454
rect 518642 26898 518878 27134
rect 1706 14218 1942 14454
rect 1706 13898 1942 14134
rect 109998 14218 110234 14454
rect 109998 13898 110234 14134
rect 119706 14218 119942 14454
rect 119706 13898 119942 14134
rect 517982 14218 518218 14454
rect 517982 13898 518218 14134
<< metal5 >>
rect 1104 156856 522836 157496
rect 1104 144454 2200 144496
rect 1104 144218 1706 144454
rect 1942 144218 2200 144454
rect 1104 144134 2200 144218
rect 1104 143898 1706 144134
rect 1942 143898 2200 144134
rect 1104 143856 2200 143898
rect 109800 144454 120200 144496
rect 109800 144218 109998 144454
rect 110234 144218 119706 144454
rect 119942 144218 120200 144454
rect 109800 144134 120200 144218
rect 109800 143898 109998 144134
rect 110234 143898 119706 144134
rect 119942 143898 120200 144134
rect 109800 143856 120200 143898
rect 517800 144454 522836 144496
rect 517800 144218 517982 144454
rect 518218 144218 522836 144454
rect 517800 144134 522836 144218
rect 517800 143898 517982 144134
rect 518218 143898 522836 144134
rect 517800 143856 522836 143898
rect 1072 131454 2200 131496
rect 1072 131218 1096 131454
rect 1332 131218 2200 131454
rect 1072 131134 2200 131218
rect 1072 130898 1096 131134
rect 1332 130898 2200 131134
rect 1072 130856 2200 130898
rect 109800 131454 120200 131496
rect 109800 131218 110658 131454
rect 110894 131218 119046 131454
rect 119282 131218 120200 131454
rect 109800 131134 120200 131218
rect 109800 130898 110658 131134
rect 110894 130898 119046 131134
rect 119282 130898 120200 131134
rect 109800 130856 120200 130898
rect 517800 131454 522836 131496
rect 517800 131218 518642 131454
rect 518878 131218 522836 131454
rect 517800 131134 522836 131218
rect 517800 130898 518642 131134
rect 518878 130898 522836 131134
rect 517800 130856 522836 130898
rect 1104 118454 2200 118496
rect 1104 118218 1706 118454
rect 1942 118218 2200 118454
rect 1104 118134 2200 118218
rect 1104 117898 1706 118134
rect 1942 117898 2200 118134
rect 1104 117856 2200 117898
rect 109800 118454 120200 118496
rect 109800 118218 109998 118454
rect 110234 118218 119706 118454
rect 119942 118218 120200 118454
rect 109800 118134 120200 118218
rect 109800 117898 109998 118134
rect 110234 117898 119706 118134
rect 119942 117898 120200 118134
rect 109800 117856 120200 117898
rect 517800 118454 522836 118496
rect 517800 118218 517982 118454
rect 518218 118218 522836 118454
rect 517800 118134 522836 118218
rect 517800 117898 517982 118134
rect 518218 117898 522836 118134
rect 517800 117856 522836 117898
rect 1072 105454 2200 105496
rect 1072 105218 1096 105454
rect 1332 105218 2200 105454
rect 1072 105134 2200 105218
rect 1072 104898 1096 105134
rect 1332 104898 2200 105134
rect 1072 104856 2200 104898
rect 109800 105454 120200 105496
rect 109800 105218 110658 105454
rect 110894 105218 119046 105454
rect 119282 105218 120200 105454
rect 109800 105134 120200 105218
rect 109800 104898 110658 105134
rect 110894 104898 119046 105134
rect 119282 104898 120200 105134
rect 109800 104856 120200 104898
rect 517800 105454 522836 105496
rect 517800 105218 518642 105454
rect 518878 105218 522836 105454
rect 517800 105134 522836 105218
rect 517800 104898 518642 105134
rect 518878 104898 522836 105134
rect 517800 104856 522836 104898
rect 1104 92454 2200 92496
rect 1104 92218 1706 92454
rect 1942 92218 2200 92454
rect 1104 92134 2200 92218
rect 1104 91898 1706 92134
rect 1942 91898 2200 92134
rect 1104 91856 2200 91898
rect 109800 92454 120200 92496
rect 109800 92218 109998 92454
rect 110234 92218 119706 92454
rect 119942 92218 120200 92454
rect 109800 92134 120200 92218
rect 109800 91898 109998 92134
rect 110234 91898 119706 92134
rect 119942 91898 120200 92134
rect 109800 91856 120200 91898
rect 517800 92454 522836 92496
rect 517800 92218 517982 92454
rect 518218 92218 522836 92454
rect 517800 92134 522836 92218
rect 517800 91898 517982 92134
rect 518218 91898 522836 92134
rect 517800 91856 522836 91898
rect 1072 79454 2200 79496
rect 1072 79218 1096 79454
rect 1332 79218 2200 79454
rect 1072 79134 2200 79218
rect 1072 78898 1096 79134
rect 1332 78898 2200 79134
rect 1072 78856 2200 78898
rect 109800 79454 120200 79496
rect 109800 79218 110658 79454
rect 110894 79218 119046 79454
rect 119282 79218 120200 79454
rect 109800 79134 120200 79218
rect 109800 78898 110658 79134
rect 110894 78898 119046 79134
rect 119282 78898 120200 79134
rect 109800 78856 120200 78898
rect 517800 79454 522836 79496
rect 517800 79218 518642 79454
rect 518878 79218 522836 79454
rect 517800 79134 522836 79218
rect 517800 78898 518642 79134
rect 518878 78898 522836 79134
rect 517800 78856 522836 78898
rect 1104 66454 2200 66496
rect 1104 66218 1706 66454
rect 1942 66218 2200 66454
rect 1104 66134 2200 66218
rect 1104 65898 1706 66134
rect 1942 65898 2200 66134
rect 1104 65856 2200 65898
rect 109800 66454 120200 66496
rect 109800 66218 109998 66454
rect 110234 66218 119706 66454
rect 119942 66218 120200 66454
rect 109800 66134 120200 66218
rect 109800 65898 109998 66134
rect 110234 65898 119706 66134
rect 119942 65898 120200 66134
rect 109800 65856 120200 65898
rect 517800 66454 522836 66496
rect 517800 66218 517982 66454
rect 518218 66218 522836 66454
rect 517800 66134 522836 66218
rect 517800 65898 517982 66134
rect 518218 65898 522836 66134
rect 517800 65856 522836 65898
rect 1072 53454 2200 53496
rect 1072 53218 1096 53454
rect 1332 53218 2200 53454
rect 1072 53134 2200 53218
rect 1072 52898 1096 53134
rect 1332 52898 2200 53134
rect 1072 52856 2200 52898
rect 109800 53454 120200 53496
rect 109800 53218 110658 53454
rect 110894 53218 119046 53454
rect 119282 53218 120200 53454
rect 109800 53134 120200 53218
rect 109800 52898 110658 53134
rect 110894 52898 119046 53134
rect 119282 52898 120200 53134
rect 109800 52856 120200 52898
rect 517800 53454 522836 53496
rect 517800 53218 518642 53454
rect 518878 53218 522836 53454
rect 517800 53134 522836 53218
rect 517800 52898 518642 53134
rect 518878 52898 522836 53134
rect 517800 52856 522836 52898
rect 1104 40454 2200 40496
rect 1104 40218 1706 40454
rect 1942 40218 2200 40454
rect 1104 40134 2200 40218
rect 1104 39898 1706 40134
rect 1942 39898 2200 40134
rect 1104 39856 2200 39898
rect 109800 40454 120200 40496
rect 109800 40218 109998 40454
rect 110234 40218 119706 40454
rect 119942 40218 120200 40454
rect 109800 40134 120200 40218
rect 109800 39898 109998 40134
rect 110234 39898 119706 40134
rect 119942 39898 120200 40134
rect 109800 39856 120200 39898
rect 517800 40454 522836 40496
rect 517800 40218 517982 40454
rect 518218 40218 522836 40454
rect 517800 40134 522836 40218
rect 517800 39898 517982 40134
rect 518218 39898 522836 40134
rect 517800 39856 522836 39898
rect 1072 27454 2200 27496
rect 1072 27218 1096 27454
rect 1332 27218 2200 27454
rect 1072 27134 2200 27218
rect 1072 26898 1096 27134
rect 1332 26898 2200 27134
rect 1072 26856 2200 26898
rect 109800 27454 120200 27496
rect 109800 27218 110658 27454
rect 110894 27218 119046 27454
rect 119282 27218 120200 27454
rect 109800 27134 120200 27218
rect 109800 26898 110658 27134
rect 110894 26898 119046 27134
rect 119282 26898 120200 27134
rect 109800 26856 120200 26898
rect 517800 27454 522836 27496
rect 517800 27218 518642 27454
rect 518878 27218 522836 27454
rect 517800 27134 522836 27218
rect 517800 26898 518642 27134
rect 518878 26898 522836 27134
rect 517800 26856 522836 26898
rect 1104 14454 2200 14496
rect 1104 14218 1706 14454
rect 1942 14218 2200 14454
rect 1104 14134 2200 14218
rect 1104 13898 1706 14134
rect 1942 13898 2200 14134
rect 1104 13856 2200 13898
rect 109800 14454 120200 14496
rect 109800 14218 109998 14454
rect 110234 14218 119706 14454
rect 119942 14218 120200 14454
rect 109800 14134 120200 14218
rect 109800 13898 109998 14134
rect 110234 13898 119706 14134
rect 119942 13898 120200 14134
rect 109800 13856 120200 13898
rect 517800 14454 522836 14496
rect 517800 14218 517982 14454
rect 518218 14218 522836 14454
rect 517800 14134 522836 14218
rect 517800 13898 517982 14134
rect 518218 13898 522836 14134
rect 517800 13856 522836 13898
use mgmt_core  core
timestamp 1637416515
transform 1 0 119000 0 1 2000
box 0 0 400000 148000
use DFFRAM  DFFRAM
timestamp 1637416515
transform 1 0 1000 0 1 2000
box 4 0 110000 148000
<< labels >>
rlabel metal5 s 1104 26856 2200 27496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 26856 120200 27496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 26856 522836 27496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 52856 2200 53496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 52856 120200 53496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 52856 522836 53496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 78856 2200 79496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 78856 120200 79496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 78856 522836 79496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 104856 2200 105496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 104856 120200 105496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 104856 522836 105496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 130856 2200 131496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 130856 120200 131496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 130856 522836 131496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 156856 522836 157496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 13856 2200 14496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 13856 120200 14496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 13856 522836 14496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 39856 2200 40496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 39856 120200 40496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 39856 522836 40496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 65856 2200 66496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 65856 120200 66496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 65856 522836 66496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 91856 2200 92496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 91856 120200 92496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 91856 522836 92496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 117856 2200 118496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 117856 120200 118496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 117856 522836 118496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 143856 2200 144496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 143856 120200 144496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 143856 522836 144496 6 VPWR
port 1 nsew power input
rlabel metal2 s 294786 -400 294842 800 6 core_clk
port 2 nsew signal input
rlabel metal2 s 98274 -400 98330 800 6 core_rstn
port 3 nsew signal input
rlabel metal3 s 523200 64472 524400 64592 6 debug_in
port 4 nsew signal input
rlabel metal3 s 523200 65968 524400 66088 6 debug_mode
port 5 nsew signal tristate
rlabel metal3 s 523200 67464 524400 67584 6 debug_oeb
port 6 nsew signal tristate
rlabel metal3 s 523200 68960 524400 69080 6 debug_out
port 7 nsew signal tristate
rlabel metal3 s 523200 144848 524400 144968 6 flash_clk
port 8 nsew signal tristate
rlabel metal3 s 523200 143352 524400 143472 6 flash_csb
port 9 nsew signal tristate
rlabel metal3 s 523200 146480 524400 146600 6 flash_io0_di
port 10 nsew signal input
rlabel metal3 s 523200 147976 524400 148096 6 flash_io0_do
port 11 nsew signal tristate
rlabel metal3 s 523200 149472 524400 149592 6 flash_io0_oeb
port 12 nsew signal tristate
rlabel metal3 s 523200 150968 524400 151088 6 flash_io1_di
port 13 nsew signal input
rlabel metal3 s 523200 152464 524400 152584 6 flash_io1_do
port 14 nsew signal tristate
rlabel metal3 s 523200 153960 524400 154080 6 flash_io1_oeb
port 15 nsew signal tristate
rlabel metal3 s 523200 155592 524400 155712 6 flash_io2_di
port 16 nsew signal input
rlabel metal3 s 523200 157088 524400 157208 6 flash_io2_do
port 17 nsew signal tristate
rlabel metal3 s 523200 158584 524400 158704 6 flash_io2_oeb
port 18 nsew signal tristate
rlabel metal3 s 523200 160080 524400 160200 6 flash_io3_di
port 19 nsew signal input
rlabel metal3 s 523200 161576 524400 161696 6 flash_io3_do
port 20 nsew signal tristate
rlabel metal3 s 523200 163072 524400 163192 6 flash_io3_oeb
port 21 nsew signal tristate
rlabel metal2 s 32770 -400 32826 800 6 gpio_in_pad
port 22 nsew signal input
rlabel metal2 s 163778 -400 163834 800 6 gpio_inenb_pad
port 23 nsew signal tristate
rlabel metal2 s 229282 -400 229338 800 6 gpio_mode0_pad
port 24 nsew signal tristate
rlabel metal2 s 360290 -400 360346 800 6 gpio_mode1_pad
port 25 nsew signal tristate
rlabel metal2 s 425794 -400 425850 800 6 gpio_out_pad
port 26 nsew signal tristate
rlabel metal2 s 491298 -400 491354 800 6 gpio_outenb_pad
port 27 nsew signal tristate
rlabel metal3 s 523200 91808 524400 91928 6 hk_ack_i
port 28 nsew signal input
rlabel metal3 s 523200 94800 524400 94920 6 hk_dat_i[0]
port 29 nsew signal input
rlabel metal3 s 523200 110032 524400 110152 6 hk_dat_i[10]
port 30 nsew signal input
rlabel metal3 s 523200 111528 524400 111648 6 hk_dat_i[11]
port 31 nsew signal input
rlabel metal3 s 523200 113024 524400 113144 6 hk_dat_i[12]
port 32 nsew signal input
rlabel metal3 s 523200 114520 524400 114640 6 hk_dat_i[13]
port 33 nsew signal input
rlabel metal3 s 523200 116016 524400 116136 6 hk_dat_i[14]
port 34 nsew signal input
rlabel metal3 s 523200 117512 524400 117632 6 hk_dat_i[15]
port 35 nsew signal input
rlabel metal3 s 523200 119144 524400 119264 6 hk_dat_i[16]
port 36 nsew signal input
rlabel metal3 s 523200 120640 524400 120760 6 hk_dat_i[17]
port 37 nsew signal input
rlabel metal3 s 523200 122136 524400 122256 6 hk_dat_i[18]
port 38 nsew signal input
rlabel metal3 s 523200 123632 524400 123752 6 hk_dat_i[19]
port 39 nsew signal input
rlabel metal3 s 523200 96296 524400 96416 6 hk_dat_i[1]
port 40 nsew signal input
rlabel metal3 s 523200 125128 524400 125248 6 hk_dat_i[20]
port 41 nsew signal input
rlabel metal3 s 523200 126624 524400 126744 6 hk_dat_i[21]
port 42 nsew signal input
rlabel metal3 s 523200 128256 524400 128376 6 hk_dat_i[22]
port 43 nsew signal input
rlabel metal3 s 523200 129752 524400 129872 6 hk_dat_i[23]
port 44 nsew signal input
rlabel metal3 s 523200 131248 524400 131368 6 hk_dat_i[24]
port 45 nsew signal input
rlabel metal3 s 523200 132744 524400 132864 6 hk_dat_i[25]
port 46 nsew signal input
rlabel metal3 s 523200 134240 524400 134360 6 hk_dat_i[26]
port 47 nsew signal input
rlabel metal3 s 523200 135736 524400 135856 6 hk_dat_i[27]
port 48 nsew signal input
rlabel metal3 s 523200 137368 524400 137488 6 hk_dat_i[28]
port 49 nsew signal input
rlabel metal3 s 523200 138864 524400 138984 6 hk_dat_i[29]
port 50 nsew signal input
rlabel metal3 s 523200 97792 524400 97912 6 hk_dat_i[2]
port 51 nsew signal input
rlabel metal3 s 523200 140360 524400 140480 6 hk_dat_i[30]
port 52 nsew signal input
rlabel metal3 s 523200 141856 524400 141976 6 hk_dat_i[31]
port 53 nsew signal input
rlabel metal3 s 523200 99288 524400 99408 6 hk_dat_i[3]
port 54 nsew signal input
rlabel metal3 s 523200 100920 524400 101040 6 hk_dat_i[4]
port 55 nsew signal input
rlabel metal3 s 523200 102416 524400 102536 6 hk_dat_i[5]
port 56 nsew signal input
rlabel metal3 s 523200 103912 524400 104032 6 hk_dat_i[6]
port 57 nsew signal input
rlabel metal3 s 523200 105408 524400 105528 6 hk_dat_i[7]
port 58 nsew signal input
rlabel metal3 s 523200 106904 524400 107024 6 hk_dat_i[8]
port 59 nsew signal input
rlabel metal3 s 523200 108400 524400 108520 6 hk_dat_i[9]
port 60 nsew signal input
rlabel metal3 s 523200 93304 524400 93424 6 hk_stb_o
port 61 nsew signal tristate
rlabel metal2 s 521842 163200 521898 164400 6 irq[0]
port 62 nsew signal input
rlabel metal2 s 522670 163200 522726 164400 6 irq[1]
port 63 nsew signal input
rlabel metal2 s 523498 163200 523554 164400 6 irq[2]
port 64 nsew signal input
rlabel metal3 s 523200 75080 524400 75200 6 irq[3]
port 65 nsew signal input
rlabel metal3 s 523200 73584 524400 73704 6 irq[4]
port 66 nsew signal input
rlabel metal3 s 523200 71952 524400 72072 6 irq[5]
port 67 nsew signal input
rlabel metal2 s 386 163200 442 164400 6 la_iena[0]
port 68 nsew signal tristate
rlabel metal2 s 336830 163200 336886 164400 6 la_iena[100]
port 69 nsew signal tristate
rlabel metal2 s 340142 163200 340198 164400 6 la_iena[101]
port 70 nsew signal tristate
rlabel metal2 s 343546 163200 343602 164400 6 la_iena[102]
port 71 nsew signal tristate
rlabel metal2 s 346858 163200 346914 164400 6 la_iena[103]
port 72 nsew signal tristate
rlabel metal2 s 350262 163200 350318 164400 6 la_iena[104]
port 73 nsew signal tristate
rlabel metal2 s 353666 163200 353722 164400 6 la_iena[105]
port 74 nsew signal tristate
rlabel metal2 s 356978 163200 357034 164400 6 la_iena[106]
port 75 nsew signal tristate
rlabel metal2 s 360382 163200 360438 164400 6 la_iena[107]
port 76 nsew signal tristate
rlabel metal2 s 363694 163200 363750 164400 6 la_iena[108]
port 77 nsew signal tristate
rlabel metal2 s 367098 163200 367154 164400 6 la_iena[109]
port 78 nsew signal tristate
rlabel metal2 s 33966 163200 34022 164400 6 la_iena[10]
port 79 nsew signal tristate
rlabel metal2 s 370410 163200 370466 164400 6 la_iena[110]
port 80 nsew signal tristate
rlabel metal2 s 373814 163200 373870 164400 6 la_iena[111]
port 81 nsew signal tristate
rlabel metal2 s 377218 163200 377274 164400 6 la_iena[112]
port 82 nsew signal tristate
rlabel metal2 s 380530 163200 380586 164400 6 la_iena[113]
port 83 nsew signal tristate
rlabel metal2 s 383934 163200 383990 164400 6 la_iena[114]
port 84 nsew signal tristate
rlabel metal2 s 387246 163200 387302 164400 6 la_iena[115]
port 85 nsew signal tristate
rlabel metal2 s 390650 163200 390706 164400 6 la_iena[116]
port 86 nsew signal tristate
rlabel metal2 s 393962 163200 394018 164400 6 la_iena[117]
port 87 nsew signal tristate
rlabel metal2 s 397366 163200 397422 164400 6 la_iena[118]
port 88 nsew signal tristate
rlabel metal2 s 400770 163200 400826 164400 6 la_iena[119]
port 89 nsew signal tristate
rlabel metal2 s 37370 163200 37426 164400 6 la_iena[11]
port 90 nsew signal tristate
rlabel metal2 s 404082 163200 404138 164400 6 la_iena[120]
port 91 nsew signal tristate
rlabel metal2 s 407486 163200 407542 164400 6 la_iena[121]
port 92 nsew signal tristate
rlabel metal2 s 410798 163200 410854 164400 6 la_iena[122]
port 93 nsew signal tristate
rlabel metal2 s 414202 163200 414258 164400 6 la_iena[123]
port 94 nsew signal tristate
rlabel metal2 s 417514 163200 417570 164400 6 la_iena[124]
port 95 nsew signal tristate
rlabel metal2 s 420918 163200 420974 164400 6 la_iena[125]
port 96 nsew signal tristate
rlabel metal2 s 424322 163200 424378 164400 6 la_iena[126]
port 97 nsew signal tristate
rlabel metal2 s 427634 163200 427690 164400 6 la_iena[127]
port 98 nsew signal tristate
rlabel metal2 s 40682 163200 40738 164400 6 la_iena[12]
port 99 nsew signal tristate
rlabel metal2 s 44086 163200 44142 164400 6 la_iena[13]
port 100 nsew signal tristate
rlabel metal2 s 47490 163200 47546 164400 6 la_iena[14]
port 101 nsew signal tristate
rlabel metal2 s 50802 163200 50858 164400 6 la_iena[15]
port 102 nsew signal tristate
rlabel metal2 s 54206 163200 54262 164400 6 la_iena[16]
port 103 nsew signal tristate
rlabel metal2 s 57518 163200 57574 164400 6 la_iena[17]
port 104 nsew signal tristate
rlabel metal2 s 60922 163200 60978 164400 6 la_iena[18]
port 105 nsew signal tristate
rlabel metal2 s 64234 163200 64290 164400 6 la_iena[19]
port 106 nsew signal tristate
rlabel metal2 s 3698 163200 3754 164400 6 la_iena[1]
port 107 nsew signal tristate
rlabel metal2 s 67638 163200 67694 164400 6 la_iena[20]
port 108 nsew signal tristate
rlabel metal2 s 71042 163200 71098 164400 6 la_iena[21]
port 109 nsew signal tristate
rlabel metal2 s 74354 163200 74410 164400 6 la_iena[22]
port 110 nsew signal tristate
rlabel metal2 s 77758 163200 77814 164400 6 la_iena[23]
port 111 nsew signal tristate
rlabel metal2 s 81070 163200 81126 164400 6 la_iena[24]
port 112 nsew signal tristate
rlabel metal2 s 84474 163200 84530 164400 6 la_iena[25]
port 113 nsew signal tristate
rlabel metal2 s 87786 163200 87842 164400 6 la_iena[26]
port 114 nsew signal tristate
rlabel metal2 s 91190 163200 91246 164400 6 la_iena[27]
port 115 nsew signal tristate
rlabel metal2 s 94594 163200 94650 164400 6 la_iena[28]
port 116 nsew signal tristate
rlabel metal2 s 97906 163200 97962 164400 6 la_iena[29]
port 117 nsew signal tristate
rlabel metal2 s 7102 163200 7158 164400 6 la_iena[2]
port 118 nsew signal tristate
rlabel metal2 s 101310 163200 101366 164400 6 la_iena[30]
port 119 nsew signal tristate
rlabel metal2 s 104622 163200 104678 164400 6 la_iena[31]
port 120 nsew signal tristate
rlabel metal2 s 108026 163200 108082 164400 6 la_iena[32]
port 121 nsew signal tristate
rlabel metal2 s 111338 163200 111394 164400 6 la_iena[33]
port 122 nsew signal tristate
rlabel metal2 s 114742 163200 114798 164400 6 la_iena[34]
port 123 nsew signal tristate
rlabel metal2 s 118146 163200 118202 164400 6 la_iena[35]
port 124 nsew signal tristate
rlabel metal2 s 121458 163200 121514 164400 6 la_iena[36]
port 125 nsew signal tristate
rlabel metal2 s 124862 163200 124918 164400 6 la_iena[37]
port 126 nsew signal tristate
rlabel metal2 s 128174 163200 128230 164400 6 la_iena[38]
port 127 nsew signal tristate
rlabel metal2 s 131578 163200 131634 164400 6 la_iena[39]
port 128 nsew signal tristate
rlabel metal2 s 10414 163200 10470 164400 6 la_iena[3]
port 129 nsew signal tristate
rlabel metal2 s 134890 163200 134946 164400 6 la_iena[40]
port 130 nsew signal tristate
rlabel metal2 s 138294 163200 138350 164400 6 la_iena[41]
port 131 nsew signal tristate
rlabel metal2 s 141698 163200 141754 164400 6 la_iena[42]
port 132 nsew signal tristate
rlabel metal2 s 145010 163200 145066 164400 6 la_iena[43]
port 133 nsew signal tristate
rlabel metal2 s 148414 163200 148470 164400 6 la_iena[44]
port 134 nsew signal tristate
rlabel metal2 s 151726 163200 151782 164400 6 la_iena[45]
port 135 nsew signal tristate
rlabel metal2 s 155130 163200 155186 164400 6 la_iena[46]
port 136 nsew signal tristate
rlabel metal2 s 158442 163200 158498 164400 6 la_iena[47]
port 137 nsew signal tristate
rlabel metal2 s 161846 163200 161902 164400 6 la_iena[48]
port 138 nsew signal tristate
rlabel metal2 s 165250 163200 165306 164400 6 la_iena[49]
port 139 nsew signal tristate
rlabel metal2 s 13818 163200 13874 164400 6 la_iena[4]
port 140 nsew signal tristate
rlabel metal2 s 168562 163200 168618 164400 6 la_iena[50]
port 141 nsew signal tristate
rlabel metal2 s 171966 163200 172022 164400 6 la_iena[51]
port 142 nsew signal tristate
rlabel metal2 s 175278 163200 175334 164400 6 la_iena[52]
port 143 nsew signal tristate
rlabel metal2 s 178682 163200 178738 164400 6 la_iena[53]
port 144 nsew signal tristate
rlabel metal2 s 181994 163200 182050 164400 6 la_iena[54]
port 145 nsew signal tristate
rlabel metal2 s 185398 163200 185454 164400 6 la_iena[55]
port 146 nsew signal tristate
rlabel metal2 s 188802 163200 188858 164400 6 la_iena[56]
port 147 nsew signal tristate
rlabel metal2 s 192114 163200 192170 164400 6 la_iena[57]
port 148 nsew signal tristate
rlabel metal2 s 195518 163200 195574 164400 6 la_iena[58]
port 149 nsew signal tristate
rlabel metal2 s 198830 163200 198886 164400 6 la_iena[59]
port 150 nsew signal tristate
rlabel metal2 s 17130 163200 17186 164400 6 la_iena[5]
port 151 nsew signal tristate
rlabel metal2 s 202234 163200 202290 164400 6 la_iena[60]
port 152 nsew signal tristate
rlabel metal2 s 205546 163200 205602 164400 6 la_iena[61]
port 153 nsew signal tristate
rlabel metal2 s 208950 163200 209006 164400 6 la_iena[62]
port 154 nsew signal tristate
rlabel metal2 s 212354 163200 212410 164400 6 la_iena[63]
port 155 nsew signal tristate
rlabel metal2 s 215666 163200 215722 164400 6 la_iena[64]
port 156 nsew signal tristate
rlabel metal2 s 219070 163200 219126 164400 6 la_iena[65]
port 157 nsew signal tristate
rlabel metal2 s 222382 163200 222438 164400 6 la_iena[66]
port 158 nsew signal tristate
rlabel metal2 s 225786 163200 225842 164400 6 la_iena[67]
port 159 nsew signal tristate
rlabel metal2 s 229098 163200 229154 164400 6 la_iena[68]
port 160 nsew signal tristate
rlabel metal2 s 232502 163200 232558 164400 6 la_iena[69]
port 161 nsew signal tristate
rlabel metal2 s 20534 163200 20590 164400 6 la_iena[6]
port 162 nsew signal tristate
rlabel metal2 s 235906 163200 235962 164400 6 la_iena[70]
port 163 nsew signal tristate
rlabel metal2 s 239218 163200 239274 164400 6 la_iena[71]
port 164 nsew signal tristate
rlabel metal2 s 242622 163200 242678 164400 6 la_iena[72]
port 165 nsew signal tristate
rlabel metal2 s 245934 163200 245990 164400 6 la_iena[73]
port 166 nsew signal tristate
rlabel metal2 s 249338 163200 249394 164400 6 la_iena[74]
port 167 nsew signal tristate
rlabel metal2 s 252650 163200 252706 164400 6 la_iena[75]
port 168 nsew signal tristate
rlabel metal2 s 256054 163200 256110 164400 6 la_iena[76]
port 169 nsew signal tristate
rlabel metal2 s 259458 163200 259514 164400 6 la_iena[77]
port 170 nsew signal tristate
rlabel metal2 s 262770 163200 262826 164400 6 la_iena[78]
port 171 nsew signal tristate
rlabel metal2 s 266174 163200 266230 164400 6 la_iena[79]
port 172 nsew signal tristate
rlabel metal2 s 23938 163200 23994 164400 6 la_iena[7]
port 173 nsew signal tristate
rlabel metal2 s 269486 163200 269542 164400 6 la_iena[80]
port 174 nsew signal tristate
rlabel metal2 s 272890 163200 272946 164400 6 la_iena[81]
port 175 nsew signal tristate
rlabel metal2 s 276202 163200 276258 164400 6 la_iena[82]
port 176 nsew signal tristate
rlabel metal2 s 279606 163200 279662 164400 6 la_iena[83]
port 177 nsew signal tristate
rlabel metal2 s 283010 163200 283066 164400 6 la_iena[84]
port 178 nsew signal tristate
rlabel metal2 s 286322 163200 286378 164400 6 la_iena[85]
port 179 nsew signal tristate
rlabel metal2 s 289726 163200 289782 164400 6 la_iena[86]
port 180 nsew signal tristate
rlabel metal2 s 293038 163200 293094 164400 6 la_iena[87]
port 181 nsew signal tristate
rlabel metal2 s 296442 163200 296498 164400 6 la_iena[88]
port 182 nsew signal tristate
rlabel metal2 s 299754 163200 299810 164400 6 la_iena[89]
port 183 nsew signal tristate
rlabel metal2 s 27250 163200 27306 164400 6 la_iena[8]
port 184 nsew signal tristate
rlabel metal2 s 303158 163200 303214 164400 6 la_iena[90]
port 185 nsew signal tristate
rlabel metal2 s 306562 163200 306618 164400 6 la_iena[91]
port 186 nsew signal tristate
rlabel metal2 s 309874 163200 309930 164400 6 la_iena[92]
port 187 nsew signal tristate
rlabel metal2 s 313278 163200 313334 164400 6 la_iena[93]
port 188 nsew signal tristate
rlabel metal2 s 316590 163200 316646 164400 6 la_iena[94]
port 189 nsew signal tristate
rlabel metal2 s 319994 163200 320050 164400 6 la_iena[95]
port 190 nsew signal tristate
rlabel metal2 s 323306 163200 323362 164400 6 la_iena[96]
port 191 nsew signal tristate
rlabel metal2 s 326710 163200 326766 164400 6 la_iena[97]
port 192 nsew signal tristate
rlabel metal2 s 330114 163200 330170 164400 6 la_iena[98]
port 193 nsew signal tristate
rlabel metal2 s 333426 163200 333482 164400 6 la_iena[99]
port 194 nsew signal tristate
rlabel metal2 s 30654 163200 30710 164400 6 la_iena[9]
port 195 nsew signal tristate
rlabel metal2 s 1214 163200 1270 164400 6 la_input[0]
port 196 nsew signal input
rlabel metal2 s 337658 163200 337714 164400 6 la_input[100]
port 197 nsew signal input
rlabel metal2 s 340970 163200 341026 164400 6 la_input[101]
port 198 nsew signal input
rlabel metal2 s 344374 163200 344430 164400 6 la_input[102]
port 199 nsew signal input
rlabel metal2 s 347778 163200 347834 164400 6 la_input[103]
port 200 nsew signal input
rlabel metal2 s 351090 163200 351146 164400 6 la_input[104]
port 201 nsew signal input
rlabel metal2 s 354494 163200 354550 164400 6 la_input[105]
port 202 nsew signal input
rlabel metal2 s 357806 163200 357862 164400 6 la_input[106]
port 203 nsew signal input
rlabel metal2 s 361210 163200 361266 164400 6 la_input[107]
port 204 nsew signal input
rlabel metal2 s 364522 163200 364578 164400 6 la_input[108]
port 205 nsew signal input
rlabel metal2 s 367926 163200 367982 164400 6 la_input[109]
port 206 nsew signal input
rlabel metal2 s 34794 163200 34850 164400 6 la_input[10]
port 207 nsew signal input
rlabel metal2 s 371330 163200 371386 164400 6 la_input[110]
port 208 nsew signal input
rlabel metal2 s 374642 163200 374698 164400 6 la_input[111]
port 209 nsew signal input
rlabel metal2 s 378046 163200 378102 164400 6 la_input[112]
port 210 nsew signal input
rlabel metal2 s 381358 163200 381414 164400 6 la_input[113]
port 211 nsew signal input
rlabel metal2 s 384762 163200 384818 164400 6 la_input[114]
port 212 nsew signal input
rlabel metal2 s 388074 163200 388130 164400 6 la_input[115]
port 213 nsew signal input
rlabel metal2 s 391478 163200 391534 164400 6 la_input[116]
port 214 nsew signal input
rlabel metal2 s 394882 163200 394938 164400 6 la_input[117]
port 215 nsew signal input
rlabel metal2 s 398194 163200 398250 164400 6 la_input[118]
port 216 nsew signal input
rlabel metal2 s 401598 163200 401654 164400 6 la_input[119]
port 217 nsew signal input
rlabel metal2 s 38198 163200 38254 164400 6 la_input[11]
port 218 nsew signal input
rlabel metal2 s 404910 163200 404966 164400 6 la_input[120]
port 219 nsew signal input
rlabel metal2 s 408314 163200 408370 164400 6 la_input[121]
port 220 nsew signal input
rlabel metal2 s 411626 163200 411682 164400 6 la_input[122]
port 221 nsew signal input
rlabel metal2 s 415030 163200 415086 164400 6 la_input[123]
port 222 nsew signal input
rlabel metal2 s 418434 163200 418490 164400 6 la_input[124]
port 223 nsew signal input
rlabel metal2 s 421746 163200 421802 164400 6 la_input[125]
port 224 nsew signal input
rlabel metal2 s 425150 163200 425206 164400 6 la_input[126]
port 225 nsew signal input
rlabel metal2 s 428462 163200 428518 164400 6 la_input[127]
port 226 nsew signal input
rlabel metal2 s 41602 163200 41658 164400 6 la_input[12]
port 227 nsew signal input
rlabel metal2 s 44914 163200 44970 164400 6 la_input[13]
port 228 nsew signal input
rlabel metal2 s 48318 163200 48374 164400 6 la_input[14]
port 229 nsew signal input
rlabel metal2 s 51630 163200 51686 164400 6 la_input[15]
port 230 nsew signal input
rlabel metal2 s 55034 163200 55090 164400 6 la_input[16]
port 231 nsew signal input
rlabel metal2 s 58346 163200 58402 164400 6 la_input[17]
port 232 nsew signal input
rlabel metal2 s 61750 163200 61806 164400 6 la_input[18]
port 233 nsew signal input
rlabel metal2 s 65154 163200 65210 164400 6 la_input[19]
port 234 nsew signal input
rlabel metal2 s 4526 163200 4582 164400 6 la_input[1]
port 235 nsew signal input
rlabel metal2 s 68466 163200 68522 164400 6 la_input[20]
port 236 nsew signal input
rlabel metal2 s 71870 163200 71926 164400 6 la_input[21]
port 237 nsew signal input
rlabel metal2 s 75182 163200 75238 164400 6 la_input[22]
port 238 nsew signal input
rlabel metal2 s 78586 163200 78642 164400 6 la_input[23]
port 239 nsew signal input
rlabel metal2 s 81898 163200 81954 164400 6 la_input[24]
port 240 nsew signal input
rlabel metal2 s 85302 163200 85358 164400 6 la_input[25]
port 241 nsew signal input
rlabel metal2 s 88706 163200 88762 164400 6 la_input[26]
port 242 nsew signal input
rlabel metal2 s 92018 163200 92074 164400 6 la_input[27]
port 243 nsew signal input
rlabel metal2 s 95422 163200 95478 164400 6 la_input[28]
port 244 nsew signal input
rlabel metal2 s 98734 163200 98790 164400 6 la_input[29]
port 245 nsew signal input
rlabel metal2 s 7930 163200 7986 164400 6 la_input[2]
port 246 nsew signal input
rlabel metal2 s 102138 163200 102194 164400 6 la_input[30]
port 247 nsew signal input
rlabel metal2 s 105450 163200 105506 164400 6 la_input[31]
port 248 nsew signal input
rlabel metal2 s 108854 163200 108910 164400 6 la_input[32]
port 249 nsew signal input
rlabel metal2 s 112258 163200 112314 164400 6 la_input[33]
port 250 nsew signal input
rlabel metal2 s 115570 163200 115626 164400 6 la_input[34]
port 251 nsew signal input
rlabel metal2 s 118974 163200 119030 164400 6 la_input[35]
port 252 nsew signal input
rlabel metal2 s 122286 163200 122342 164400 6 la_input[36]
port 253 nsew signal input
rlabel metal2 s 125690 163200 125746 164400 6 la_input[37]
port 254 nsew signal input
rlabel metal2 s 129002 163200 129058 164400 6 la_input[38]
port 255 nsew signal input
rlabel metal2 s 132406 163200 132462 164400 6 la_input[39]
port 256 nsew signal input
rlabel metal2 s 11242 163200 11298 164400 6 la_input[3]
port 257 nsew signal input
rlabel metal2 s 135810 163200 135866 164400 6 la_input[40]
port 258 nsew signal input
rlabel metal2 s 139122 163200 139178 164400 6 la_input[41]
port 259 nsew signal input
rlabel metal2 s 142526 163200 142582 164400 6 la_input[42]
port 260 nsew signal input
rlabel metal2 s 145838 163200 145894 164400 6 la_input[43]
port 261 nsew signal input
rlabel metal2 s 149242 163200 149298 164400 6 la_input[44]
port 262 nsew signal input
rlabel metal2 s 152554 163200 152610 164400 6 la_input[45]
port 263 nsew signal input
rlabel metal2 s 155958 163200 156014 164400 6 la_input[46]
port 264 nsew signal input
rlabel metal2 s 159362 163200 159418 164400 6 la_input[47]
port 265 nsew signal input
rlabel metal2 s 162674 163200 162730 164400 6 la_input[48]
port 266 nsew signal input
rlabel metal2 s 166078 163200 166134 164400 6 la_input[49]
port 267 nsew signal input
rlabel metal2 s 14646 163200 14702 164400 6 la_input[4]
port 268 nsew signal input
rlabel metal2 s 169390 163200 169446 164400 6 la_input[50]
port 269 nsew signal input
rlabel metal2 s 172794 163200 172850 164400 6 la_input[51]
port 270 nsew signal input
rlabel metal2 s 176106 163200 176162 164400 6 la_input[52]
port 271 nsew signal input
rlabel metal2 s 179510 163200 179566 164400 6 la_input[53]
port 272 nsew signal input
rlabel metal2 s 182914 163200 182970 164400 6 la_input[54]
port 273 nsew signal input
rlabel metal2 s 186226 163200 186282 164400 6 la_input[55]
port 274 nsew signal input
rlabel metal2 s 189630 163200 189686 164400 6 la_input[56]
port 275 nsew signal input
rlabel metal2 s 192942 163200 192998 164400 6 la_input[57]
port 276 nsew signal input
rlabel metal2 s 196346 163200 196402 164400 6 la_input[58]
port 277 nsew signal input
rlabel metal2 s 199658 163200 199714 164400 6 la_input[59]
port 278 nsew signal input
rlabel metal2 s 18050 163200 18106 164400 6 la_input[5]
port 279 nsew signal input
rlabel metal2 s 203062 163200 203118 164400 6 la_input[60]
port 280 nsew signal input
rlabel metal2 s 206466 163200 206522 164400 6 la_input[61]
port 281 nsew signal input
rlabel metal2 s 209778 163200 209834 164400 6 la_input[62]
port 282 nsew signal input
rlabel metal2 s 213182 163200 213238 164400 6 la_input[63]
port 283 nsew signal input
rlabel metal2 s 216494 163200 216550 164400 6 la_input[64]
port 284 nsew signal input
rlabel metal2 s 219898 163200 219954 164400 6 la_input[65]
port 285 nsew signal input
rlabel metal2 s 223210 163200 223266 164400 6 la_input[66]
port 286 nsew signal input
rlabel metal2 s 226614 163200 226670 164400 6 la_input[67]
port 287 nsew signal input
rlabel metal2 s 230018 163200 230074 164400 6 la_input[68]
port 288 nsew signal input
rlabel metal2 s 233330 163200 233386 164400 6 la_input[69]
port 289 nsew signal input
rlabel metal2 s 21362 163200 21418 164400 6 la_input[6]
port 290 nsew signal input
rlabel metal2 s 236734 163200 236790 164400 6 la_input[70]
port 291 nsew signal input
rlabel metal2 s 240046 163200 240102 164400 6 la_input[71]
port 292 nsew signal input
rlabel metal2 s 243450 163200 243506 164400 6 la_input[72]
port 293 nsew signal input
rlabel metal2 s 246762 163200 246818 164400 6 la_input[73]
port 294 nsew signal input
rlabel metal2 s 250166 163200 250222 164400 6 la_input[74]
port 295 nsew signal input
rlabel metal2 s 253570 163200 253626 164400 6 la_input[75]
port 296 nsew signal input
rlabel metal2 s 256882 163200 256938 164400 6 la_input[76]
port 297 nsew signal input
rlabel metal2 s 260286 163200 260342 164400 6 la_input[77]
port 298 nsew signal input
rlabel metal2 s 263598 163200 263654 164400 6 la_input[78]
port 299 nsew signal input
rlabel metal2 s 267002 163200 267058 164400 6 la_input[79]
port 300 nsew signal input
rlabel metal2 s 24766 163200 24822 164400 6 la_input[7]
port 301 nsew signal input
rlabel metal2 s 270314 163200 270370 164400 6 la_input[80]
port 302 nsew signal input
rlabel metal2 s 273718 163200 273774 164400 6 la_input[81]
port 303 nsew signal input
rlabel metal2 s 277122 163200 277178 164400 6 la_input[82]
port 304 nsew signal input
rlabel metal2 s 280434 163200 280490 164400 6 la_input[83]
port 305 nsew signal input
rlabel metal2 s 283838 163200 283894 164400 6 la_input[84]
port 306 nsew signal input
rlabel metal2 s 287150 163200 287206 164400 6 la_input[85]
port 307 nsew signal input
rlabel metal2 s 290554 163200 290610 164400 6 la_input[86]
port 308 nsew signal input
rlabel metal2 s 293866 163200 293922 164400 6 la_input[87]
port 309 nsew signal input
rlabel metal2 s 297270 163200 297326 164400 6 la_input[88]
port 310 nsew signal input
rlabel metal2 s 300674 163200 300730 164400 6 la_input[89]
port 311 nsew signal input
rlabel metal2 s 28078 163200 28134 164400 6 la_input[8]
port 312 nsew signal input
rlabel metal2 s 303986 163200 304042 164400 6 la_input[90]
port 313 nsew signal input
rlabel metal2 s 307390 163200 307446 164400 6 la_input[91]
port 314 nsew signal input
rlabel metal2 s 310702 163200 310758 164400 6 la_input[92]
port 315 nsew signal input
rlabel metal2 s 314106 163200 314162 164400 6 la_input[93]
port 316 nsew signal input
rlabel metal2 s 317418 163200 317474 164400 6 la_input[94]
port 317 nsew signal input
rlabel metal2 s 320822 163200 320878 164400 6 la_input[95]
port 318 nsew signal input
rlabel metal2 s 324226 163200 324282 164400 6 la_input[96]
port 319 nsew signal input
rlabel metal2 s 327538 163200 327594 164400 6 la_input[97]
port 320 nsew signal input
rlabel metal2 s 330942 163200 330998 164400 6 la_input[98]
port 321 nsew signal input
rlabel metal2 s 334254 163200 334310 164400 6 la_input[99]
port 322 nsew signal input
rlabel metal2 s 31482 163200 31538 164400 6 la_input[9]
port 323 nsew signal input
rlabel metal2 s 2042 163200 2098 164400 6 la_oenb[0]
port 324 nsew signal tristate
rlabel metal2 s 338486 163200 338542 164400 6 la_oenb[100]
port 325 nsew signal tristate
rlabel metal2 s 341890 163200 341946 164400 6 la_oenb[101]
port 326 nsew signal tristate
rlabel metal2 s 345202 163200 345258 164400 6 la_oenb[102]
port 327 nsew signal tristate
rlabel metal2 s 348606 163200 348662 164400 6 la_oenb[103]
port 328 nsew signal tristate
rlabel metal2 s 351918 163200 351974 164400 6 la_oenb[104]
port 329 nsew signal tristate
rlabel metal2 s 355322 163200 355378 164400 6 la_oenb[105]
port 330 nsew signal tristate
rlabel metal2 s 358634 163200 358690 164400 6 la_oenb[106]
port 331 nsew signal tristate
rlabel metal2 s 362038 163200 362094 164400 6 la_oenb[107]
port 332 nsew signal tristate
rlabel metal2 s 365442 163200 365498 164400 6 la_oenb[108]
port 333 nsew signal tristate
rlabel metal2 s 368754 163200 368810 164400 6 la_oenb[109]
port 334 nsew signal tristate
rlabel metal2 s 35714 163200 35770 164400 6 la_oenb[10]
port 335 nsew signal tristate
rlabel metal2 s 372158 163200 372214 164400 6 la_oenb[110]
port 336 nsew signal tristate
rlabel metal2 s 375470 163200 375526 164400 6 la_oenb[111]
port 337 nsew signal tristate
rlabel metal2 s 378874 163200 378930 164400 6 la_oenb[112]
port 338 nsew signal tristate
rlabel metal2 s 382186 163200 382242 164400 6 la_oenb[113]
port 339 nsew signal tristate
rlabel metal2 s 385590 163200 385646 164400 6 la_oenb[114]
port 340 nsew signal tristate
rlabel metal2 s 388994 163200 389050 164400 6 la_oenb[115]
port 341 nsew signal tristate
rlabel metal2 s 392306 163200 392362 164400 6 la_oenb[116]
port 342 nsew signal tristate
rlabel metal2 s 395710 163200 395766 164400 6 la_oenb[117]
port 343 nsew signal tristate
rlabel metal2 s 399022 163200 399078 164400 6 la_oenb[118]
port 344 nsew signal tristate
rlabel metal2 s 402426 163200 402482 164400 6 la_oenb[119]
port 345 nsew signal tristate
rlabel metal2 s 39026 163200 39082 164400 6 la_oenb[11]
port 346 nsew signal tristate
rlabel metal2 s 405738 163200 405794 164400 6 la_oenb[120]
port 347 nsew signal tristate
rlabel metal2 s 409142 163200 409198 164400 6 la_oenb[121]
port 348 nsew signal tristate
rlabel metal2 s 412546 163200 412602 164400 6 la_oenb[122]
port 349 nsew signal tristate
rlabel metal2 s 415858 163200 415914 164400 6 la_oenb[123]
port 350 nsew signal tristate
rlabel metal2 s 419262 163200 419318 164400 6 la_oenb[124]
port 351 nsew signal tristate
rlabel metal2 s 422574 163200 422630 164400 6 la_oenb[125]
port 352 nsew signal tristate
rlabel metal2 s 425978 163200 426034 164400 6 la_oenb[126]
port 353 nsew signal tristate
rlabel metal2 s 429290 163200 429346 164400 6 la_oenb[127]
port 354 nsew signal tristate
rlabel metal2 s 42430 163200 42486 164400 6 la_oenb[12]
port 355 nsew signal tristate
rlabel metal2 s 45742 163200 45798 164400 6 la_oenb[13]
port 356 nsew signal tristate
rlabel metal2 s 49146 163200 49202 164400 6 la_oenb[14]
port 357 nsew signal tristate
rlabel metal2 s 52458 163200 52514 164400 6 la_oenb[15]
port 358 nsew signal tristate
rlabel metal2 s 55862 163200 55918 164400 6 la_oenb[16]
port 359 nsew signal tristate
rlabel metal2 s 59266 163200 59322 164400 6 la_oenb[17]
port 360 nsew signal tristate
rlabel metal2 s 62578 163200 62634 164400 6 la_oenb[18]
port 361 nsew signal tristate
rlabel metal2 s 65982 163200 66038 164400 6 la_oenb[19]
port 362 nsew signal tristate
rlabel metal2 s 5354 163200 5410 164400 6 la_oenb[1]
port 363 nsew signal tristate
rlabel metal2 s 69294 163200 69350 164400 6 la_oenb[20]
port 364 nsew signal tristate
rlabel metal2 s 72698 163200 72754 164400 6 la_oenb[21]
port 365 nsew signal tristate
rlabel metal2 s 76010 163200 76066 164400 6 la_oenb[22]
port 366 nsew signal tristate
rlabel metal2 s 79414 163200 79470 164400 6 la_oenb[23]
port 367 nsew signal tristate
rlabel metal2 s 82818 163200 82874 164400 6 la_oenb[24]
port 368 nsew signal tristate
rlabel metal2 s 86130 163200 86186 164400 6 la_oenb[25]
port 369 nsew signal tristate
rlabel metal2 s 89534 163200 89590 164400 6 la_oenb[26]
port 370 nsew signal tristate
rlabel metal2 s 92846 163200 92902 164400 6 la_oenb[27]
port 371 nsew signal tristate
rlabel metal2 s 96250 163200 96306 164400 6 la_oenb[28]
port 372 nsew signal tristate
rlabel metal2 s 99562 163200 99618 164400 6 la_oenb[29]
port 373 nsew signal tristate
rlabel metal2 s 8758 163200 8814 164400 6 la_oenb[2]
port 374 nsew signal tristate
rlabel metal2 s 102966 163200 103022 164400 6 la_oenb[30]
port 375 nsew signal tristate
rlabel metal2 s 106370 163200 106426 164400 6 la_oenb[31]
port 376 nsew signal tristate
rlabel metal2 s 109682 163200 109738 164400 6 la_oenb[32]
port 377 nsew signal tristate
rlabel metal2 s 113086 163200 113142 164400 6 la_oenb[33]
port 378 nsew signal tristate
rlabel metal2 s 116398 163200 116454 164400 6 la_oenb[34]
port 379 nsew signal tristate
rlabel metal2 s 119802 163200 119858 164400 6 la_oenb[35]
port 380 nsew signal tristate
rlabel metal2 s 123114 163200 123170 164400 6 la_oenb[36]
port 381 nsew signal tristate
rlabel metal2 s 126518 163200 126574 164400 6 la_oenb[37]
port 382 nsew signal tristate
rlabel metal2 s 129922 163200 129978 164400 6 la_oenb[38]
port 383 nsew signal tristate
rlabel metal2 s 133234 163200 133290 164400 6 la_oenb[39]
port 384 nsew signal tristate
rlabel metal2 s 12162 163200 12218 164400 6 la_oenb[3]
port 385 nsew signal tristate
rlabel metal2 s 136638 163200 136694 164400 6 la_oenb[40]
port 386 nsew signal tristate
rlabel metal2 s 139950 163200 140006 164400 6 la_oenb[41]
port 387 nsew signal tristate
rlabel metal2 s 143354 163200 143410 164400 6 la_oenb[42]
port 388 nsew signal tristate
rlabel metal2 s 146666 163200 146722 164400 6 la_oenb[43]
port 389 nsew signal tristate
rlabel metal2 s 150070 163200 150126 164400 6 la_oenb[44]
port 390 nsew signal tristate
rlabel metal2 s 153474 163200 153530 164400 6 la_oenb[45]
port 391 nsew signal tristate
rlabel metal2 s 156786 163200 156842 164400 6 la_oenb[46]
port 392 nsew signal tristate
rlabel metal2 s 160190 163200 160246 164400 6 la_oenb[47]
port 393 nsew signal tristate
rlabel metal2 s 163502 163200 163558 164400 6 la_oenb[48]
port 394 nsew signal tristate
rlabel metal2 s 166906 163200 166962 164400 6 la_oenb[49]
port 395 nsew signal tristate
rlabel metal2 s 15474 163200 15530 164400 6 la_oenb[4]
port 396 nsew signal tristate
rlabel metal2 s 170218 163200 170274 164400 6 la_oenb[50]
port 397 nsew signal tristate
rlabel metal2 s 173622 163200 173678 164400 6 la_oenb[51]
port 398 nsew signal tristate
rlabel metal2 s 177026 163200 177082 164400 6 la_oenb[52]
port 399 nsew signal tristate
rlabel metal2 s 180338 163200 180394 164400 6 la_oenb[53]
port 400 nsew signal tristate
rlabel metal2 s 183742 163200 183798 164400 6 la_oenb[54]
port 401 nsew signal tristate
rlabel metal2 s 187054 163200 187110 164400 6 la_oenb[55]
port 402 nsew signal tristate
rlabel metal2 s 190458 163200 190514 164400 6 la_oenb[56]
port 403 nsew signal tristate
rlabel metal2 s 193770 163200 193826 164400 6 la_oenb[57]
port 404 nsew signal tristate
rlabel metal2 s 197174 163200 197230 164400 6 la_oenb[58]
port 405 nsew signal tristate
rlabel metal2 s 200578 163200 200634 164400 6 la_oenb[59]
port 406 nsew signal tristate
rlabel metal2 s 18878 163200 18934 164400 6 la_oenb[5]
port 407 nsew signal tristate
rlabel metal2 s 203890 163200 203946 164400 6 la_oenb[60]
port 408 nsew signal tristate
rlabel metal2 s 207294 163200 207350 164400 6 la_oenb[61]
port 409 nsew signal tristate
rlabel metal2 s 210606 163200 210662 164400 6 la_oenb[62]
port 410 nsew signal tristate
rlabel metal2 s 214010 163200 214066 164400 6 la_oenb[63]
port 411 nsew signal tristate
rlabel metal2 s 217322 163200 217378 164400 6 la_oenb[64]
port 412 nsew signal tristate
rlabel metal2 s 220726 163200 220782 164400 6 la_oenb[65]
port 413 nsew signal tristate
rlabel metal2 s 224130 163200 224186 164400 6 la_oenb[66]
port 414 nsew signal tristate
rlabel metal2 s 227442 163200 227498 164400 6 la_oenb[67]
port 415 nsew signal tristate
rlabel metal2 s 230846 163200 230902 164400 6 la_oenb[68]
port 416 nsew signal tristate
rlabel metal2 s 234158 163200 234214 164400 6 la_oenb[69]
port 417 nsew signal tristate
rlabel metal2 s 22190 163200 22246 164400 6 la_oenb[6]
port 418 nsew signal tristate
rlabel metal2 s 237562 163200 237618 164400 6 la_oenb[70]
port 419 nsew signal tristate
rlabel metal2 s 240874 163200 240930 164400 6 la_oenb[71]
port 420 nsew signal tristate
rlabel metal2 s 244278 163200 244334 164400 6 la_oenb[72]
port 421 nsew signal tristate
rlabel metal2 s 247682 163200 247738 164400 6 la_oenb[73]
port 422 nsew signal tristate
rlabel metal2 s 250994 163200 251050 164400 6 la_oenb[74]
port 423 nsew signal tristate
rlabel metal2 s 254398 163200 254454 164400 6 la_oenb[75]
port 424 nsew signal tristate
rlabel metal2 s 257710 163200 257766 164400 6 la_oenb[76]
port 425 nsew signal tristate
rlabel metal2 s 261114 163200 261170 164400 6 la_oenb[77]
port 426 nsew signal tristate
rlabel metal2 s 264426 163200 264482 164400 6 la_oenb[78]
port 427 nsew signal tristate
rlabel metal2 s 267830 163200 267886 164400 6 la_oenb[79]
port 428 nsew signal tristate
rlabel metal2 s 25594 163200 25650 164400 6 la_oenb[7]
port 429 nsew signal tristate
rlabel metal2 s 271234 163200 271290 164400 6 la_oenb[80]
port 430 nsew signal tristate
rlabel metal2 s 274546 163200 274602 164400 6 la_oenb[81]
port 431 nsew signal tristate
rlabel metal2 s 277950 163200 278006 164400 6 la_oenb[82]
port 432 nsew signal tristate
rlabel metal2 s 281262 163200 281318 164400 6 la_oenb[83]
port 433 nsew signal tristate
rlabel metal2 s 284666 163200 284722 164400 6 la_oenb[84]
port 434 nsew signal tristate
rlabel metal2 s 287978 163200 288034 164400 6 la_oenb[85]
port 435 nsew signal tristate
rlabel metal2 s 291382 163200 291438 164400 6 la_oenb[86]
port 436 nsew signal tristate
rlabel metal2 s 294786 163200 294842 164400 6 la_oenb[87]
port 437 nsew signal tristate
rlabel metal2 s 298098 163200 298154 164400 6 la_oenb[88]
port 438 nsew signal tristate
rlabel metal2 s 301502 163200 301558 164400 6 la_oenb[89]
port 439 nsew signal tristate
rlabel metal2 s 28906 163200 28962 164400 6 la_oenb[8]
port 440 nsew signal tristate
rlabel metal2 s 304814 163200 304870 164400 6 la_oenb[90]
port 441 nsew signal tristate
rlabel metal2 s 308218 163200 308274 164400 6 la_oenb[91]
port 442 nsew signal tristate
rlabel metal2 s 311530 163200 311586 164400 6 la_oenb[92]
port 443 nsew signal tristate
rlabel metal2 s 314934 163200 314990 164400 6 la_oenb[93]
port 444 nsew signal tristate
rlabel metal2 s 318338 163200 318394 164400 6 la_oenb[94]
port 445 nsew signal tristate
rlabel metal2 s 321650 163200 321706 164400 6 la_oenb[95]
port 446 nsew signal tristate
rlabel metal2 s 325054 163200 325110 164400 6 la_oenb[96]
port 447 nsew signal tristate
rlabel metal2 s 328366 163200 328422 164400 6 la_oenb[97]
port 448 nsew signal tristate
rlabel metal2 s 331770 163200 331826 164400 6 la_oenb[98]
port 449 nsew signal tristate
rlabel metal2 s 335082 163200 335138 164400 6 la_oenb[99]
port 450 nsew signal tristate
rlabel metal2 s 32310 163200 32366 164400 6 la_oenb[9]
port 451 nsew signal tristate
rlabel metal2 s 2870 163200 2926 164400 6 la_output[0]
port 452 nsew signal tristate
rlabel metal2 s 339314 163200 339370 164400 6 la_output[100]
port 453 nsew signal tristate
rlabel metal2 s 342718 163200 342774 164400 6 la_output[101]
port 454 nsew signal tristate
rlabel metal2 s 346030 163200 346086 164400 6 la_output[102]
port 455 nsew signal tristate
rlabel metal2 s 349434 163200 349490 164400 6 la_output[103]
port 456 nsew signal tristate
rlabel metal2 s 352746 163200 352802 164400 6 la_output[104]
port 457 nsew signal tristate
rlabel metal2 s 356150 163200 356206 164400 6 la_output[105]
port 458 nsew signal tristate
rlabel metal2 s 359554 163200 359610 164400 6 la_output[106]
port 459 nsew signal tristate
rlabel metal2 s 362866 163200 362922 164400 6 la_output[107]
port 460 nsew signal tristate
rlabel metal2 s 366270 163200 366326 164400 6 la_output[108]
port 461 nsew signal tristate
rlabel metal2 s 369582 163200 369638 164400 6 la_output[109]
port 462 nsew signal tristate
rlabel metal2 s 36542 163200 36598 164400 6 la_output[10]
port 463 nsew signal tristate
rlabel metal2 s 372986 163200 373042 164400 6 la_output[110]
port 464 nsew signal tristate
rlabel metal2 s 376298 163200 376354 164400 6 la_output[111]
port 465 nsew signal tristate
rlabel metal2 s 379702 163200 379758 164400 6 la_output[112]
port 466 nsew signal tristate
rlabel metal2 s 383106 163200 383162 164400 6 la_output[113]
port 467 nsew signal tristate
rlabel metal2 s 386418 163200 386474 164400 6 la_output[114]
port 468 nsew signal tristate
rlabel metal2 s 389822 163200 389878 164400 6 la_output[115]
port 469 nsew signal tristate
rlabel metal2 s 393134 163200 393190 164400 6 la_output[116]
port 470 nsew signal tristate
rlabel metal2 s 396538 163200 396594 164400 6 la_output[117]
port 471 nsew signal tristate
rlabel metal2 s 399850 163200 399906 164400 6 la_output[118]
port 472 nsew signal tristate
rlabel metal2 s 403254 163200 403310 164400 6 la_output[119]
port 473 nsew signal tristate
rlabel metal2 s 39854 163200 39910 164400 6 la_output[11]
port 474 nsew signal tristate
rlabel metal2 s 406658 163200 406714 164400 6 la_output[120]
port 475 nsew signal tristate
rlabel metal2 s 409970 163200 410026 164400 6 la_output[121]
port 476 nsew signal tristate
rlabel metal2 s 413374 163200 413430 164400 6 la_output[122]
port 477 nsew signal tristate
rlabel metal2 s 416686 163200 416742 164400 6 la_output[123]
port 478 nsew signal tristate
rlabel metal2 s 420090 163200 420146 164400 6 la_output[124]
port 479 nsew signal tristate
rlabel metal2 s 423402 163200 423458 164400 6 la_output[125]
port 480 nsew signal tristate
rlabel metal2 s 426806 163200 426862 164400 6 la_output[126]
port 481 nsew signal tristate
rlabel metal2 s 430210 163200 430266 164400 6 la_output[127]
port 482 nsew signal tristate
rlabel metal2 s 43258 163200 43314 164400 6 la_output[12]
port 483 nsew signal tristate
rlabel metal2 s 46570 163200 46626 164400 6 la_output[13]
port 484 nsew signal tristate
rlabel metal2 s 49974 163200 50030 164400 6 la_output[14]
port 485 nsew signal tristate
rlabel metal2 s 53378 163200 53434 164400 6 la_output[15]
port 486 nsew signal tristate
rlabel metal2 s 56690 163200 56746 164400 6 la_output[16]
port 487 nsew signal tristate
rlabel metal2 s 60094 163200 60150 164400 6 la_output[17]
port 488 nsew signal tristate
rlabel metal2 s 63406 163200 63462 164400 6 la_output[18]
port 489 nsew signal tristate
rlabel metal2 s 66810 163200 66866 164400 6 la_output[19]
port 490 nsew signal tristate
rlabel metal2 s 6274 163200 6330 164400 6 la_output[1]
port 491 nsew signal tristate
rlabel metal2 s 70122 163200 70178 164400 6 la_output[20]
port 492 nsew signal tristate
rlabel metal2 s 73526 163200 73582 164400 6 la_output[21]
port 493 nsew signal tristate
rlabel metal2 s 76930 163200 76986 164400 6 la_output[22]
port 494 nsew signal tristate
rlabel metal2 s 80242 163200 80298 164400 6 la_output[23]
port 495 nsew signal tristate
rlabel metal2 s 83646 163200 83702 164400 6 la_output[24]
port 496 nsew signal tristate
rlabel metal2 s 86958 163200 87014 164400 6 la_output[25]
port 497 nsew signal tristate
rlabel metal2 s 90362 163200 90418 164400 6 la_output[26]
port 498 nsew signal tristate
rlabel metal2 s 93674 163200 93730 164400 6 la_output[27]
port 499 nsew signal tristate
rlabel metal2 s 97078 163200 97134 164400 6 la_output[28]
port 500 nsew signal tristate
rlabel metal2 s 100482 163200 100538 164400 6 la_output[29]
port 501 nsew signal tristate
rlabel metal2 s 9586 163200 9642 164400 6 la_output[2]
port 502 nsew signal tristate
rlabel metal2 s 103794 163200 103850 164400 6 la_output[30]
port 503 nsew signal tristate
rlabel metal2 s 107198 163200 107254 164400 6 la_output[31]
port 504 nsew signal tristate
rlabel metal2 s 110510 163200 110566 164400 6 la_output[32]
port 505 nsew signal tristate
rlabel metal2 s 113914 163200 113970 164400 6 la_output[33]
port 506 nsew signal tristate
rlabel metal2 s 117226 163200 117282 164400 6 la_output[34]
port 507 nsew signal tristate
rlabel metal2 s 120630 163200 120686 164400 6 la_output[35]
port 508 nsew signal tristate
rlabel metal2 s 124034 163200 124090 164400 6 la_output[36]
port 509 nsew signal tristate
rlabel metal2 s 127346 163200 127402 164400 6 la_output[37]
port 510 nsew signal tristate
rlabel metal2 s 130750 163200 130806 164400 6 la_output[38]
port 511 nsew signal tristate
rlabel metal2 s 134062 163200 134118 164400 6 la_output[39]
port 512 nsew signal tristate
rlabel metal2 s 12990 163200 13046 164400 6 la_output[3]
port 513 nsew signal tristate
rlabel metal2 s 137466 163200 137522 164400 6 la_output[40]
port 514 nsew signal tristate
rlabel metal2 s 140778 163200 140834 164400 6 la_output[41]
port 515 nsew signal tristate
rlabel metal2 s 144182 163200 144238 164400 6 la_output[42]
port 516 nsew signal tristate
rlabel metal2 s 147586 163200 147642 164400 6 la_output[43]
port 517 nsew signal tristate
rlabel metal2 s 150898 163200 150954 164400 6 la_output[44]
port 518 nsew signal tristate
rlabel metal2 s 154302 163200 154358 164400 6 la_output[45]
port 519 nsew signal tristate
rlabel metal2 s 157614 163200 157670 164400 6 la_output[46]
port 520 nsew signal tristate
rlabel metal2 s 161018 163200 161074 164400 6 la_output[47]
port 521 nsew signal tristate
rlabel metal2 s 164330 163200 164386 164400 6 la_output[48]
port 522 nsew signal tristate
rlabel metal2 s 167734 163200 167790 164400 6 la_output[49]
port 523 nsew signal tristate
rlabel metal2 s 16302 163200 16358 164400 6 la_output[4]
port 524 nsew signal tristate
rlabel metal2 s 171138 163200 171194 164400 6 la_output[50]
port 525 nsew signal tristate
rlabel metal2 s 174450 163200 174506 164400 6 la_output[51]
port 526 nsew signal tristate
rlabel metal2 s 177854 163200 177910 164400 6 la_output[52]
port 527 nsew signal tristate
rlabel metal2 s 181166 163200 181222 164400 6 la_output[53]
port 528 nsew signal tristate
rlabel metal2 s 184570 163200 184626 164400 6 la_output[54]
port 529 nsew signal tristate
rlabel metal2 s 187882 163200 187938 164400 6 la_output[55]
port 530 nsew signal tristate
rlabel metal2 s 191286 163200 191342 164400 6 la_output[56]
port 531 nsew signal tristate
rlabel metal2 s 194690 163200 194746 164400 6 la_output[57]
port 532 nsew signal tristate
rlabel metal2 s 198002 163200 198058 164400 6 la_output[58]
port 533 nsew signal tristate
rlabel metal2 s 201406 163200 201462 164400 6 la_output[59]
port 534 nsew signal tristate
rlabel metal2 s 19706 163200 19762 164400 6 la_output[5]
port 535 nsew signal tristate
rlabel metal2 s 204718 163200 204774 164400 6 la_output[60]
port 536 nsew signal tristate
rlabel metal2 s 208122 163200 208178 164400 6 la_output[61]
port 537 nsew signal tristate
rlabel metal2 s 211434 163200 211490 164400 6 la_output[62]
port 538 nsew signal tristate
rlabel metal2 s 214838 163200 214894 164400 6 la_output[63]
port 539 nsew signal tristate
rlabel metal2 s 218242 163200 218298 164400 6 la_output[64]
port 540 nsew signal tristate
rlabel metal2 s 221554 163200 221610 164400 6 la_output[65]
port 541 nsew signal tristate
rlabel metal2 s 224958 163200 225014 164400 6 la_output[66]
port 542 nsew signal tristate
rlabel metal2 s 228270 163200 228326 164400 6 la_output[67]
port 543 nsew signal tristate
rlabel metal2 s 231674 163200 231730 164400 6 la_output[68]
port 544 nsew signal tristate
rlabel metal2 s 234986 163200 235042 164400 6 la_output[69]
port 545 nsew signal tristate
rlabel metal2 s 23018 163200 23074 164400 6 la_output[6]
port 546 nsew signal tristate
rlabel metal2 s 238390 163200 238446 164400 6 la_output[70]
port 547 nsew signal tristate
rlabel metal2 s 241794 163200 241850 164400 6 la_output[71]
port 548 nsew signal tristate
rlabel metal2 s 245106 163200 245162 164400 6 la_output[72]
port 549 nsew signal tristate
rlabel metal2 s 248510 163200 248566 164400 6 la_output[73]
port 550 nsew signal tristate
rlabel metal2 s 251822 163200 251878 164400 6 la_output[74]
port 551 nsew signal tristate
rlabel metal2 s 255226 163200 255282 164400 6 la_output[75]
port 552 nsew signal tristate
rlabel metal2 s 258538 163200 258594 164400 6 la_output[76]
port 553 nsew signal tristate
rlabel metal2 s 261942 163200 261998 164400 6 la_output[77]
port 554 nsew signal tristate
rlabel metal2 s 265346 163200 265402 164400 6 la_output[78]
port 555 nsew signal tristate
rlabel metal2 s 268658 163200 268714 164400 6 la_output[79]
port 556 nsew signal tristate
rlabel metal2 s 26422 163200 26478 164400 6 la_output[7]
port 557 nsew signal tristate
rlabel metal2 s 272062 163200 272118 164400 6 la_output[80]
port 558 nsew signal tristate
rlabel metal2 s 275374 163200 275430 164400 6 la_output[81]
port 559 nsew signal tristate
rlabel metal2 s 278778 163200 278834 164400 6 la_output[82]
port 560 nsew signal tristate
rlabel metal2 s 282090 163200 282146 164400 6 la_output[83]
port 561 nsew signal tristate
rlabel metal2 s 285494 163200 285550 164400 6 la_output[84]
port 562 nsew signal tristate
rlabel metal2 s 288898 163200 288954 164400 6 la_output[85]
port 563 nsew signal tristate
rlabel metal2 s 292210 163200 292266 164400 6 la_output[86]
port 564 nsew signal tristate
rlabel metal2 s 295614 163200 295670 164400 6 la_output[87]
port 565 nsew signal tristate
rlabel metal2 s 298926 163200 298982 164400 6 la_output[88]
port 566 nsew signal tristate
rlabel metal2 s 302330 163200 302386 164400 6 la_output[89]
port 567 nsew signal tristate
rlabel metal2 s 29826 163200 29882 164400 6 la_output[8]
port 568 nsew signal tristate
rlabel metal2 s 305642 163200 305698 164400 6 la_output[90]
port 569 nsew signal tristate
rlabel metal2 s 309046 163200 309102 164400 6 la_output[91]
port 570 nsew signal tristate
rlabel metal2 s 312450 163200 312506 164400 6 la_output[92]
port 571 nsew signal tristate
rlabel metal2 s 315762 163200 315818 164400 6 la_output[93]
port 572 nsew signal tristate
rlabel metal2 s 319166 163200 319222 164400 6 la_output[94]
port 573 nsew signal tristate
rlabel metal2 s 322478 163200 322534 164400 6 la_output[95]
port 574 nsew signal tristate
rlabel metal2 s 325882 163200 325938 164400 6 la_output[96]
port 575 nsew signal tristate
rlabel metal2 s 329194 163200 329250 164400 6 la_output[97]
port 576 nsew signal tristate
rlabel metal2 s 332598 163200 332654 164400 6 la_output[98]
port 577 nsew signal tristate
rlabel metal2 s 336002 163200 336058 164400 6 la_output[99]
port 578 nsew signal tristate
rlabel metal2 s 33138 163200 33194 164400 6 la_output[9]
port 579 nsew signal tristate
rlabel metal2 s 431038 163200 431094 164400 6 mprj_ack_i
port 580 nsew signal input
rlabel metal2 s 435178 163200 435234 164400 6 mprj_adr_o[0]
port 581 nsew signal tristate
rlabel metal2 s 463790 163200 463846 164400 6 mprj_adr_o[10]
port 582 nsew signal tristate
rlabel metal2 s 466366 163200 466422 164400 6 mprj_adr_o[11]
port 583 nsew signal tristate
rlabel metal2 s 468850 163200 468906 164400 6 mprj_adr_o[12]
port 584 nsew signal tristate
rlabel metal2 s 471426 163200 471482 164400 6 mprj_adr_o[13]
port 585 nsew signal tristate
rlabel metal2 s 473910 163200 473966 164400 6 mprj_adr_o[14]
port 586 nsew signal tristate
rlabel metal2 s 476394 163200 476450 164400 6 mprj_adr_o[15]
port 587 nsew signal tristate
rlabel metal2 s 478970 163200 479026 164400 6 mprj_adr_o[16]
port 588 nsew signal tristate
rlabel metal2 s 481454 163200 481510 164400 6 mprj_adr_o[17]
port 589 nsew signal tristate
rlabel metal2 s 484030 163200 484086 164400 6 mprj_adr_o[18]
port 590 nsew signal tristate
rlabel metal2 s 486514 163200 486570 164400 6 mprj_adr_o[19]
port 591 nsew signal tristate
rlabel metal2 s 438582 163200 438638 164400 6 mprj_adr_o[1]
port 592 nsew signal tristate
rlabel metal2 s 489090 163200 489146 164400 6 mprj_adr_o[20]
port 593 nsew signal tristate
rlabel metal2 s 491574 163200 491630 164400 6 mprj_adr_o[21]
port 594 nsew signal tristate
rlabel metal2 s 494058 163200 494114 164400 6 mprj_adr_o[22]
port 595 nsew signal tristate
rlabel metal2 s 496634 163200 496690 164400 6 mprj_adr_o[23]
port 596 nsew signal tristate
rlabel metal2 s 499118 163200 499174 164400 6 mprj_adr_o[24]
port 597 nsew signal tristate
rlabel metal2 s 501694 163200 501750 164400 6 mprj_adr_o[25]
port 598 nsew signal tristate
rlabel metal2 s 504178 163200 504234 164400 6 mprj_adr_o[26]
port 599 nsew signal tristate
rlabel metal2 s 506754 163200 506810 164400 6 mprj_adr_o[27]
port 600 nsew signal tristate
rlabel metal2 s 509238 163200 509294 164400 6 mprj_adr_o[28]
port 601 nsew signal tristate
rlabel metal2 s 511722 163200 511778 164400 6 mprj_adr_o[29]
port 602 nsew signal tristate
rlabel metal2 s 441986 163200 442042 164400 6 mprj_adr_o[2]
port 603 nsew signal tristate
rlabel metal2 s 514298 163200 514354 164400 6 mprj_adr_o[30]
port 604 nsew signal tristate
rlabel metal2 s 516782 163200 516838 164400 6 mprj_adr_o[31]
port 605 nsew signal tristate
rlabel metal2 s 445298 163200 445354 164400 6 mprj_adr_o[3]
port 606 nsew signal tristate
rlabel metal2 s 448702 163200 448758 164400 6 mprj_adr_o[4]
port 607 nsew signal tristate
rlabel metal2 s 451186 163200 451242 164400 6 mprj_adr_o[5]
port 608 nsew signal tristate
rlabel metal2 s 453762 163200 453818 164400 6 mprj_adr_o[6]
port 609 nsew signal tristate
rlabel metal2 s 456246 163200 456302 164400 6 mprj_adr_o[7]
port 610 nsew signal tristate
rlabel metal2 s 458730 163200 458786 164400 6 mprj_adr_o[8]
port 611 nsew signal tristate
rlabel metal2 s 461306 163200 461362 164400 6 mprj_adr_o[9]
port 612 nsew signal tristate
rlabel metal2 s 431866 163200 431922 164400 6 mprj_cyc_o
port 613 nsew signal tristate
rlabel metal2 s 436098 163200 436154 164400 6 mprj_dat_i[0]
port 614 nsew signal input
rlabel metal2 s 464618 163200 464674 164400 6 mprj_dat_i[10]
port 615 nsew signal input
rlabel metal2 s 467194 163200 467250 164400 6 mprj_dat_i[11]
port 616 nsew signal input
rlabel metal2 s 469678 163200 469734 164400 6 mprj_dat_i[12]
port 617 nsew signal input
rlabel metal2 s 472254 163200 472310 164400 6 mprj_dat_i[13]
port 618 nsew signal input
rlabel metal2 s 474738 163200 474794 164400 6 mprj_dat_i[14]
port 619 nsew signal input
rlabel metal2 s 477314 163200 477370 164400 6 mprj_dat_i[15]
port 620 nsew signal input
rlabel metal2 s 479798 163200 479854 164400 6 mprj_dat_i[16]
port 621 nsew signal input
rlabel metal2 s 482282 163200 482338 164400 6 mprj_dat_i[17]
port 622 nsew signal input
rlabel metal2 s 484858 163200 484914 164400 6 mprj_dat_i[18]
port 623 nsew signal input
rlabel metal2 s 487342 163200 487398 164400 6 mprj_dat_i[19]
port 624 nsew signal input
rlabel metal2 s 439410 163200 439466 164400 6 mprj_dat_i[1]
port 625 nsew signal input
rlabel metal2 s 489918 163200 489974 164400 6 mprj_dat_i[20]
port 626 nsew signal input
rlabel metal2 s 492402 163200 492458 164400 6 mprj_dat_i[21]
port 627 nsew signal input
rlabel metal2 s 494978 163200 495034 164400 6 mprj_dat_i[22]
port 628 nsew signal input
rlabel metal2 s 497462 163200 497518 164400 6 mprj_dat_i[23]
port 629 nsew signal input
rlabel metal2 s 499946 163200 500002 164400 6 mprj_dat_i[24]
port 630 nsew signal input
rlabel metal2 s 502522 163200 502578 164400 6 mprj_dat_i[25]
port 631 nsew signal input
rlabel metal2 s 505006 163200 505062 164400 6 mprj_dat_i[26]
port 632 nsew signal input
rlabel metal2 s 507582 163200 507638 164400 6 mprj_dat_i[27]
port 633 nsew signal input
rlabel metal2 s 510066 163200 510122 164400 6 mprj_dat_i[28]
port 634 nsew signal input
rlabel metal2 s 512642 163200 512698 164400 6 mprj_dat_i[29]
port 635 nsew signal input
rlabel metal2 s 442814 163200 442870 164400 6 mprj_dat_i[2]
port 636 nsew signal input
rlabel metal2 s 515126 163200 515182 164400 6 mprj_dat_i[30]
port 637 nsew signal input
rlabel metal2 s 517610 163200 517666 164400 6 mprj_dat_i[31]
port 638 nsew signal input
rlabel metal2 s 446126 163200 446182 164400 6 mprj_dat_i[3]
port 639 nsew signal input
rlabel metal2 s 449530 163200 449586 164400 6 mprj_dat_i[4]
port 640 nsew signal input
rlabel metal2 s 452014 163200 452070 164400 6 mprj_dat_i[5]
port 641 nsew signal input
rlabel metal2 s 454590 163200 454646 164400 6 mprj_dat_i[6]
port 642 nsew signal input
rlabel metal2 s 457074 163200 457130 164400 6 mprj_dat_i[7]
port 643 nsew signal input
rlabel metal2 s 459650 163200 459706 164400 6 mprj_dat_i[8]
port 644 nsew signal input
rlabel metal2 s 462134 163200 462190 164400 6 mprj_dat_i[9]
port 645 nsew signal input
rlabel metal2 s 436926 163200 436982 164400 6 mprj_dat_o[0]
port 646 nsew signal tristate
rlabel metal2 s 465538 163200 465594 164400 6 mprj_dat_o[10]
port 647 nsew signal tristate
rlabel metal2 s 468022 163200 468078 164400 6 mprj_dat_o[11]
port 648 nsew signal tristate
rlabel metal2 s 470506 163200 470562 164400 6 mprj_dat_o[12]
port 649 nsew signal tristate
rlabel metal2 s 473082 163200 473138 164400 6 mprj_dat_o[13]
port 650 nsew signal tristate
rlabel metal2 s 475566 163200 475622 164400 6 mprj_dat_o[14]
port 651 nsew signal tristate
rlabel metal2 s 478142 163200 478198 164400 6 mprj_dat_o[15]
port 652 nsew signal tristate
rlabel metal2 s 480626 163200 480682 164400 6 mprj_dat_o[16]
port 653 nsew signal tristate
rlabel metal2 s 483202 163200 483258 164400 6 mprj_dat_o[17]
port 654 nsew signal tristate
rlabel metal2 s 485686 163200 485742 164400 6 mprj_dat_o[18]
port 655 nsew signal tristate
rlabel metal2 s 488170 163200 488226 164400 6 mprj_dat_o[19]
port 656 nsew signal tristate
rlabel metal2 s 440238 163200 440294 164400 6 mprj_dat_o[1]
port 657 nsew signal tristate
rlabel metal2 s 490746 163200 490802 164400 6 mprj_dat_o[20]
port 658 nsew signal tristate
rlabel metal2 s 493230 163200 493286 164400 6 mprj_dat_o[21]
port 659 nsew signal tristate
rlabel metal2 s 495806 163200 495862 164400 6 mprj_dat_o[22]
port 660 nsew signal tristate
rlabel metal2 s 498290 163200 498346 164400 6 mprj_dat_o[23]
port 661 nsew signal tristate
rlabel metal2 s 500866 163200 500922 164400 6 mprj_dat_o[24]
port 662 nsew signal tristate
rlabel metal2 s 503350 163200 503406 164400 6 mprj_dat_o[25]
port 663 nsew signal tristate
rlabel metal2 s 505834 163200 505890 164400 6 mprj_dat_o[26]
port 664 nsew signal tristate
rlabel metal2 s 508410 163200 508466 164400 6 mprj_dat_o[27]
port 665 nsew signal tristate
rlabel metal2 s 510894 163200 510950 164400 6 mprj_dat_o[28]
port 666 nsew signal tristate
rlabel metal2 s 513470 163200 513526 164400 6 mprj_dat_o[29]
port 667 nsew signal tristate
rlabel metal2 s 443642 163200 443698 164400 6 mprj_dat_o[2]
port 668 nsew signal tristate
rlabel metal2 s 515954 163200 516010 164400 6 mprj_dat_o[30]
port 669 nsew signal tristate
rlabel metal2 s 518530 163200 518586 164400 6 mprj_dat_o[31]
port 670 nsew signal tristate
rlabel metal2 s 446954 163200 447010 164400 6 mprj_dat_o[3]
port 671 nsew signal tristate
rlabel metal2 s 450358 163200 450414 164400 6 mprj_dat_o[4]
port 672 nsew signal tristate
rlabel metal2 s 452842 163200 452898 164400 6 mprj_dat_o[5]
port 673 nsew signal tristate
rlabel metal2 s 455418 163200 455474 164400 6 mprj_dat_o[6]
port 674 nsew signal tristate
rlabel metal2 s 457902 163200 457958 164400 6 mprj_dat_o[7]
port 675 nsew signal tristate
rlabel metal2 s 460478 163200 460534 164400 6 mprj_dat_o[8]
port 676 nsew signal tristate
rlabel metal2 s 462962 163200 463018 164400 6 mprj_dat_o[9]
port 677 nsew signal tristate
rlabel metal2 s 437754 163200 437810 164400 6 mprj_sel_o[0]
port 678 nsew signal tristate
rlabel metal2 s 441066 163200 441122 164400 6 mprj_sel_o[1]
port 679 nsew signal tristate
rlabel metal2 s 444470 163200 444526 164400 6 mprj_sel_o[2]
port 680 nsew signal tristate
rlabel metal2 s 447874 163200 447930 164400 6 mprj_sel_o[3]
port 681 nsew signal tristate
rlabel metal2 s 432694 163200 432750 164400 6 mprj_stb_o
port 682 nsew signal tristate
rlabel metal2 s 433522 163200 433578 164400 6 mprj_wb_iena
port 683 nsew signal tristate
rlabel metal2 s 434350 163200 434406 164400 6 mprj_we_o
port 684 nsew signal tristate
rlabel metal3 s 523200 90176 524400 90296 6 qspi_enabled
port 685 nsew signal tristate
rlabel metal3 s 523200 84192 524400 84312 6 ser_rx
port 686 nsew signal input
rlabel metal3 s 523200 85688 524400 85808 6 ser_tx
port 687 nsew signal tristate
rlabel metal3 s 523200 81064 524400 81184 6 spi_csb
port 688 nsew signal tristate
rlabel metal3 s 523200 87184 524400 87304 6 spi_enabled
port 689 nsew signal tristate
rlabel metal3 s 523200 79568 524400 79688 6 spi_sck
port 690 nsew signal tristate
rlabel metal3 s 523200 82696 524400 82816 6 spi_sdi
port 691 nsew signal input
rlabel metal3 s 523200 78072 524400 78192 6 spi_sdo
port 692 nsew signal tristate
rlabel metal3 s 523200 76576 524400 76696 6 spi_sdoenb
port 693 nsew signal tristate
rlabel metal3 s 523200 2184 524400 2304 6 sram_ro_addr[0]
port 694 nsew signal input
rlabel metal3 s 523200 3680 524400 3800 6 sram_ro_addr[1]
port 695 nsew signal input
rlabel metal3 s 523200 5176 524400 5296 6 sram_ro_addr[2]
port 696 nsew signal input
rlabel metal3 s 523200 6672 524400 6792 6 sram_ro_addr[3]
port 697 nsew signal input
rlabel metal3 s 523200 8168 524400 8288 6 sram_ro_addr[4]
port 698 nsew signal input
rlabel metal3 s 523200 9800 524400 9920 6 sram_ro_addr[5]
port 699 nsew signal input
rlabel metal3 s 523200 11296 524400 11416 6 sram_ro_addr[6]
port 700 nsew signal input
rlabel metal3 s 523200 12792 524400 12912 6 sram_ro_addr[7]
port 701 nsew signal input
rlabel metal3 s 523200 14288 524400 14408 6 sram_ro_clk
port 702 nsew signal input
rlabel metal3 s 523200 688 524400 808 6 sram_ro_csb
port 703 nsew signal input
rlabel metal3 s 523200 15784 524400 15904 6 sram_ro_data[0]
port 704 nsew signal tristate
rlabel metal3 s 523200 31016 524400 31136 6 sram_ro_data[10]
port 705 nsew signal tristate
rlabel metal3 s 523200 32512 524400 32632 6 sram_ro_data[11]
port 706 nsew signal tristate
rlabel metal3 s 523200 34008 524400 34128 6 sram_ro_data[12]
port 707 nsew signal tristate
rlabel metal3 s 523200 35504 524400 35624 6 sram_ro_data[13]
port 708 nsew signal tristate
rlabel metal3 s 523200 37136 524400 37256 6 sram_ro_data[14]
port 709 nsew signal tristate
rlabel metal3 s 523200 38632 524400 38752 6 sram_ro_data[15]
port 710 nsew signal tristate
rlabel metal3 s 523200 40128 524400 40248 6 sram_ro_data[16]
port 711 nsew signal tristate
rlabel metal3 s 523200 41624 524400 41744 6 sram_ro_data[17]
port 712 nsew signal tristate
rlabel metal3 s 523200 43120 524400 43240 6 sram_ro_data[18]
port 713 nsew signal tristate
rlabel metal3 s 523200 44616 524400 44736 6 sram_ro_data[19]
port 714 nsew signal tristate
rlabel metal3 s 523200 17280 524400 17400 6 sram_ro_data[1]
port 715 nsew signal tristate
rlabel metal3 s 523200 46248 524400 46368 6 sram_ro_data[20]
port 716 nsew signal tristate
rlabel metal3 s 523200 47744 524400 47864 6 sram_ro_data[21]
port 717 nsew signal tristate
rlabel metal3 s 523200 49240 524400 49360 6 sram_ro_data[22]
port 718 nsew signal tristate
rlabel metal3 s 523200 50736 524400 50856 6 sram_ro_data[23]
port 719 nsew signal tristate
rlabel metal3 s 523200 52232 524400 52352 6 sram_ro_data[24]
port 720 nsew signal tristate
rlabel metal3 s 523200 53728 524400 53848 6 sram_ro_data[25]
port 721 nsew signal tristate
rlabel metal3 s 523200 55360 524400 55480 6 sram_ro_data[26]
port 722 nsew signal tristate
rlabel metal3 s 523200 56856 524400 56976 6 sram_ro_data[27]
port 723 nsew signal tristate
rlabel metal3 s 523200 58352 524400 58472 6 sram_ro_data[28]
port 724 nsew signal tristate
rlabel metal3 s 523200 59848 524400 59968 6 sram_ro_data[29]
port 725 nsew signal tristate
rlabel metal3 s 523200 18912 524400 19032 6 sram_ro_data[2]
port 726 nsew signal tristate
rlabel metal3 s 523200 61344 524400 61464 6 sram_ro_data[30]
port 727 nsew signal tristate
rlabel metal3 s 523200 62840 524400 62960 6 sram_ro_data[31]
port 728 nsew signal tristate
rlabel metal3 s 523200 20408 524400 20528 6 sram_ro_data[3]
port 729 nsew signal tristate
rlabel metal3 s 523200 21904 524400 22024 6 sram_ro_data[4]
port 730 nsew signal tristate
rlabel metal3 s 523200 23400 524400 23520 6 sram_ro_data[5]
port 731 nsew signal tristate
rlabel metal3 s 523200 24896 524400 25016 6 sram_ro_data[6]
port 732 nsew signal tristate
rlabel metal3 s 523200 26392 524400 26512 6 sram_ro_data[7]
port 733 nsew signal tristate
rlabel metal3 s 523200 28024 524400 28144 6 sram_ro_data[8]
port 734 nsew signal tristate
rlabel metal3 s 523200 29520 524400 29640 6 sram_ro_data[9]
port 735 nsew signal tristate
rlabel metal3 s 523200 70456 524400 70576 6 trap
port 736 nsew signal tristate
rlabel metal3 s 523200 88680 524400 88800 6 uart_enabled
port 737 nsew signal tristate
rlabel metal2 s 519358 163200 519414 164400 6 user_irq_ena[0]
port 738 nsew signal tristate
rlabel metal2 s 520186 163200 520242 164400 6 user_irq_ena[1]
port 739 nsew signal tristate
rlabel metal2 s 521014 163200 521070 164400 6 user_irq_ena[2]
port 740 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 524000 164000
<< end >>
