magic
tech sky130A
magscale 1 2
timestamp 1636710816
<< locali >>
rect 63635 163897 63969 163931
rect 232513 160531 232547 160769
rect 471713 159715 471747 159817
rect 194609 156451 194643 156553
rect 205557 156451 205591 157165
rect 233433 156451 233467 156689
rect 340797 156451 340831 156893
rect 415501 155363 415535 155737
rect 301513 153663 301547 154445
rect 437397 154003 437431 154241
rect 538689 153935 538723 158729
rect 539517 154003 539551 158729
rect 250729 152371 250763 153017
rect 272257 152439 272291 153085
rect 60841 150535 60875 151385
rect 64429 150603 64463 151385
rect 67649 150739 67683 151317
rect 71329 150807 71363 151317
rect 74549 150875 74583 151317
rect 78137 150943 78171 151317
rect 81449 151011 81483 151317
rect 85037 151079 85071 151317
rect 88349 151147 88383 151317
rect 98837 150467 98871 151317
rect 52653 4675 52687 4845
rect 55965 4675 55999 4913
rect 62681 4675 62715 4981
rect 65993 4675 66027 5049
rect 75837 4675 75871 5117
rect 79333 4675 79367 5185
rect 82645 4675 82679 5253
rect 95985 4675 96019 5321
<< viali >>
rect 63601 163897 63635 163931
rect 63969 163897 64003 163931
rect 232513 160769 232547 160803
rect 232513 160497 232547 160531
rect 471713 159817 471747 159851
rect 471713 159681 471747 159715
rect 538689 158729 538723 158763
rect 205557 157165 205591 157199
rect 194609 156553 194643 156587
rect 194609 156417 194643 156451
rect 340797 156893 340831 156927
rect 205557 156417 205591 156451
rect 233433 156689 233467 156723
rect 233433 156417 233467 156451
rect 340797 156417 340831 156451
rect 415501 155737 415535 155771
rect 415501 155329 415535 155363
rect 301513 154445 301547 154479
rect 437397 154241 437431 154275
rect 437397 153969 437431 154003
rect 539517 158729 539551 158763
rect 539517 153969 539551 154003
rect 538689 153901 538723 153935
rect 301513 153629 301547 153663
rect 272257 153085 272291 153119
rect 250729 153017 250763 153051
rect 272257 152405 272291 152439
rect 250729 152337 250763 152371
rect 60841 151385 60875 151419
rect 64429 151385 64463 151419
rect 67649 151317 67683 151351
rect 71329 151317 71363 151351
rect 74549 151317 74583 151351
rect 78137 151317 78171 151351
rect 81449 151317 81483 151351
rect 85037 151317 85071 151351
rect 88349 151317 88383 151351
rect 88349 151113 88383 151147
rect 98837 151317 98871 151351
rect 85037 151045 85071 151079
rect 81449 150977 81483 151011
rect 78137 150909 78171 150943
rect 74549 150841 74583 150875
rect 71329 150773 71363 150807
rect 67649 150705 67683 150739
rect 64429 150569 64463 150603
rect 60841 150501 60875 150535
rect 98837 150433 98871 150467
rect 95985 5321 96019 5355
rect 82645 5253 82679 5287
rect 79333 5185 79367 5219
rect 75837 5117 75871 5151
rect 65993 5049 66027 5083
rect 62681 4981 62715 5015
rect 55965 4913 55999 4947
rect 52653 4845 52687 4879
rect 52653 4641 52687 4675
rect 55965 4641 55999 4675
rect 62681 4641 62715 4675
rect 65993 4641 66027 4675
rect 75837 4641 75871 4675
rect 79333 4641 79367 4675
rect 82645 4641 82679 4675
rect 95985 4641 96019 4675
<< metal1 >>
rect 60476 163968 60734 163996
rect 60476 163940 60504 163968
rect 60458 163888 60464 163940
rect 60516 163888 60522 163940
rect 60706 163928 60734 163968
rect 63880 163968 177160 163996
rect 63880 163940 63908 163968
rect 177132 163940 177160 163968
rect 63589 163931 63647 163937
rect 63589 163928 63601 163931
rect 60706 163900 63601 163928
rect 63589 163897 63601 163900
rect 63635 163897 63647 163931
rect 63589 163891 63647 163897
rect 63862 163888 63868 163940
rect 63920 163888 63926 163940
rect 63957 163931 64015 163937
rect 63957 163897 63969 163931
rect 64003 163928 64015 163931
rect 174446 163928 174452 163940
rect 64003 163900 174452 163928
rect 64003 163897 64015 163900
rect 63957 163891 64015 163897
rect 174446 163888 174452 163900
rect 174504 163888 174510 163940
rect 177114 163888 177120 163940
rect 177172 163888 177178 163940
rect 56778 163820 56784 163872
rect 56836 163860 56842 163872
rect 171870 163860 171876 163872
rect 56836 163832 171876 163860
rect 56836 163820 56842 163832
rect 171870 163820 171876 163832
rect 171928 163820 171934 163872
rect 53282 163752 53288 163804
rect 53340 163792 53346 163804
rect 169294 163792 169300 163804
rect 53340 163764 169300 163792
rect 53340 163752 53346 163764
rect 169294 163752 169300 163764
rect 169352 163752 169358 163804
rect 49878 163684 49884 163736
rect 49936 163724 49942 163736
rect 165614 163724 165620 163736
rect 49936 163696 165620 163724
rect 49936 163684 49942 163696
rect 165614 163684 165620 163696
rect 165672 163684 165678 163736
rect 42886 163616 42892 163668
rect 42944 163656 42950 163668
rect 161658 163656 161664 163668
rect 42944 163628 161664 163656
rect 42944 163616 42950 163628
rect 161658 163616 161664 163628
rect 161716 163616 161722 163668
rect 46382 163548 46388 163600
rect 46440 163588 46446 163600
rect 164234 163588 164240 163600
rect 46440 163560 164240 163588
rect 46440 163548 46446 163560
rect 164234 163548 164240 163560
rect 164292 163548 164298 163600
rect 35986 163480 35992 163532
rect 36044 163520 36050 163532
rect 156230 163520 156236 163532
rect 36044 163492 156236 163520
rect 36044 163480 36050 163492
rect 156230 163480 156236 163492
rect 156288 163480 156294 163532
rect 39390 163412 39396 163464
rect 39448 163452 39454 163464
rect 159174 163452 159180 163464
rect 39448 163424 159180 163452
rect 39448 163412 39454 163424
rect 159174 163412 159180 163424
rect 159232 163412 159238 163464
rect 167730 163412 167736 163464
rect 167788 163452 167794 163464
rect 254118 163452 254124 163464
rect 167788 163424 254124 163452
rect 167788 163412 167794 163424
rect 254118 163412 254124 163424
rect 254176 163412 254182 163464
rect 114830 163344 114836 163396
rect 114888 163384 114894 163396
rect 214374 163384 214380 163396
rect 114888 163356 214380 163384
rect 114888 163344 114894 163356
rect 214374 163344 214380 163356
rect 214432 163344 214438 163396
rect 112254 163276 112260 163328
rect 112312 163316 112318 163328
rect 212626 163316 212632 163328
rect 112312 163288 212632 163316
rect 112312 163276 112318 163288
rect 212626 163276 212632 163288
rect 212684 163276 212690 163328
rect 110506 163208 110512 163260
rect 110564 163248 110570 163260
rect 211798 163248 211804 163260
rect 110564 163220 211804 163248
rect 110564 163208 110570 163220
rect 211798 163208 211804 163220
rect 211856 163208 211862 163260
rect 98362 163140 98368 163192
rect 98420 163180 98426 163192
rect 202230 163180 202236 163192
rect 98420 163152 202236 163180
rect 98420 163140 98426 163152
rect 202230 163140 202236 163152
rect 202288 163140 202294 163192
rect 87874 163072 87880 163124
rect 87932 163112 87938 163124
rect 195054 163112 195060 163124
rect 87932 163084 195060 163112
rect 87932 163072 87938 163084
rect 195054 163072 195060 163084
rect 195112 163072 195118 163124
rect 84378 163004 84384 163056
rect 84436 163044 84442 163056
rect 192478 163044 192484 163056
rect 84436 163016 192484 163044
rect 84436 163004 84442 163016
rect 192478 163004 192484 163016
rect 192536 163004 192542 163056
rect 88794 162936 88800 162988
rect 88852 162976 88858 162988
rect 194686 162976 194692 162988
rect 88852 162948 194692 162976
rect 88852 162936 88858 162948
rect 194686 162936 194692 162948
rect 194744 162936 194750 162988
rect 80974 162868 80980 162920
rect 81032 162908 81038 162920
rect 189258 162908 189264 162920
rect 81032 162880 189264 162908
rect 81032 162868 81038 162880
rect 189258 162868 189264 162880
rect 189316 162868 189322 162920
rect 77478 162800 77484 162852
rect 77536 162840 77542 162852
rect 186590 162840 186596 162852
rect 77536 162812 186596 162840
rect 77536 162800 77542 162812
rect 186590 162800 186596 162812
rect 186648 162800 186654 162852
rect 79226 162732 79232 162784
rect 79284 162772 79290 162784
rect 188338 162772 188344 162784
rect 79284 162744 188344 162772
rect 79284 162732 79290 162744
rect 188338 162732 188344 162744
rect 188396 162732 188402 162784
rect 73982 162664 73988 162716
rect 74040 162704 74046 162716
rect 183554 162704 183560 162716
rect 74040 162676 183560 162704
rect 74040 162664 74046 162676
rect 183554 162664 183560 162676
rect 183612 162664 183618 162716
rect 70578 162596 70584 162648
rect 70636 162636 70642 162648
rect 182266 162636 182272 162648
rect 70636 162608 182272 162636
rect 70636 162596 70642 162608
rect 182266 162596 182272 162608
rect 182324 162596 182330 162648
rect 184934 162596 184940 162648
rect 184992 162636 184998 162648
rect 266998 162636 267004 162648
rect 184992 162608 267004 162636
rect 184992 162596 184998 162608
rect 266998 162596 267004 162608
rect 267056 162596 267062 162648
rect 165890 162528 165896 162580
rect 165948 162568 165954 162580
rect 252922 162568 252928 162580
rect 165948 162540 252928 162568
rect 165948 162528 165954 162540
rect 252922 162528 252928 162540
rect 252980 162528 252986 162580
rect 67082 162460 67088 162512
rect 67140 162500 67146 162512
rect 179690 162500 179696 162512
rect 67140 162472 179696 162500
rect 67140 162460 67146 162472
rect 179690 162460 179696 162472
rect 179748 162460 179754 162512
rect 58434 162392 58440 162444
rect 58492 162432 58498 162444
rect 172790 162432 172796 162444
rect 58492 162404 172796 162432
rect 58492 162392 58498 162404
rect 172790 162392 172796 162404
rect 172848 162392 172854 162444
rect 174538 162392 174544 162444
rect 174596 162432 174602 162444
rect 258074 162432 258080 162444
rect 174596 162404 258080 162432
rect 174596 162392 174602 162404
rect 258074 162392 258080 162404
rect 258132 162392 258138 162444
rect 160738 162324 160744 162376
rect 160796 162364 160802 162376
rect 249058 162364 249064 162376
rect 160796 162336 249064 162364
rect 160796 162324 160802 162336
rect 249058 162324 249064 162336
rect 249116 162324 249122 162376
rect 164142 162256 164148 162308
rect 164200 162296 164206 162308
rect 251634 162296 251640 162308
rect 164200 162268 251640 162296
rect 164200 162256 164206 162268
rect 251634 162256 251640 162268
rect 251692 162256 251698 162308
rect 149422 162188 149428 162240
rect 149480 162228 149486 162240
rect 240318 162228 240324 162240
rect 149480 162200 240324 162228
rect 149480 162188 149486 162200
rect 240318 162188 240324 162200
rect 240376 162188 240382 162240
rect 153746 162120 153752 162172
rect 153804 162160 153810 162172
rect 243814 162160 243820 162172
rect 153804 162132 243820 162160
rect 153804 162120 153810 162132
rect 243814 162120 243820 162132
rect 243872 162120 243878 162172
rect 141602 162052 141608 162104
rect 141660 162092 141666 162104
rect 234890 162092 234896 162104
rect 141660 162064 234896 162092
rect 141660 162052 141666 162064
rect 234890 162052 234896 162064
rect 234948 162052 234954 162104
rect 139854 161984 139860 162036
rect 139912 162024 139918 162036
rect 233418 162024 233424 162036
rect 139912 161996 233424 162024
rect 139912 161984 139918 161996
rect 233418 161984 233424 161996
rect 233476 161984 233482 162036
rect 124306 161916 124312 161968
rect 124364 161956 124370 161968
rect 221274 161956 221280 161968
rect 124364 161928 221280 161956
rect 124364 161916 124370 161928
rect 221274 161916 221280 161928
rect 221332 161916 221338 161968
rect 126054 161848 126060 161900
rect 126112 161888 126118 161900
rect 223022 161888 223028 161900
rect 126112 161860 223028 161888
rect 126112 161848 126118 161860
rect 223022 161848 223028 161860
rect 223080 161848 223086 161900
rect 31570 161780 31576 161832
rect 31628 161820 31634 161832
rect 153378 161820 153384 161832
rect 31628 161792 153384 161820
rect 31628 161780 31634 161792
rect 153378 161780 153384 161792
rect 153436 161780 153442 161832
rect 182358 161780 182364 161832
rect 182416 161820 182422 161832
rect 265066 161820 265072 161832
rect 182416 161792 265072 161820
rect 182416 161780 182422 161792
rect 265066 161780 265072 161792
rect 265124 161780 265130 161832
rect 28074 161712 28080 161764
rect 28132 161752 28138 161764
rect 150802 161752 150808 161764
rect 28132 161724 150808 161752
rect 28132 161712 28138 161724
rect 150802 161712 150808 161724
rect 150860 161712 150866 161764
rect 178034 161712 178040 161764
rect 178092 161752 178098 161764
rect 261202 161752 261208 161764
rect 178092 161724 261208 161752
rect 178092 161712 178098 161724
rect 261202 161712 261208 161724
rect 261260 161712 261266 161764
rect 24578 161644 24584 161696
rect 24636 161684 24642 161696
rect 148226 161684 148232 161696
rect 24636 161656 148232 161684
rect 24636 161644 24642 161656
rect 148226 161644 148232 161656
rect 148284 161644 148290 161696
rect 161566 161644 161572 161696
rect 161624 161684 161630 161696
rect 248506 161684 248512 161696
rect 161624 161656 248512 161684
rect 161624 161644 161630 161656
rect 248506 161644 248512 161656
rect 248564 161644 248570 161696
rect 21174 161576 21180 161628
rect 21232 161616 21238 161628
rect 145650 161616 145656 161628
rect 21232 161588 145656 161616
rect 21232 161576 21238 161588
rect 145650 161576 145656 161588
rect 145708 161576 145714 161628
rect 158990 161576 158996 161628
rect 159048 161616 159054 161628
rect 247310 161616 247316 161628
rect 159048 161588 247316 161616
rect 159048 161576 159054 161588
rect 247310 161576 247316 161588
rect 247368 161576 247374 161628
rect 17678 161508 17684 161560
rect 17736 161548 17742 161560
rect 142430 161548 142436 161560
rect 17736 161520 142436 161548
rect 17736 161508 17742 161520
rect 142430 161508 142436 161520
rect 142488 161508 142494 161560
rect 157242 161508 157248 161560
rect 157300 161548 157306 161560
rect 246390 161548 246396 161560
rect 157300 161520 246396 161548
rect 157300 161508 157306 161520
rect 246390 161508 246396 161520
rect 246448 161508 246454 161560
rect 14182 161440 14188 161492
rect 14240 161480 14246 161492
rect 140498 161480 140504 161492
rect 14240 161452 140504 161480
rect 14240 161440 14246 161452
rect 140498 161440 140504 161452
rect 140556 161440 140562 161492
rect 146846 161440 146852 161492
rect 146904 161480 146910 161492
rect 238846 161480 238852 161492
rect 146904 161452 238852 161480
rect 146904 161440 146910 161452
rect 238846 161440 238852 161452
rect 238904 161440 238910 161492
rect 243078 161440 243084 161492
rect 243136 161480 243142 161492
rect 309686 161480 309692 161492
rect 243136 161452 309692 161480
rect 243136 161440 243142 161452
rect 309686 161440 309692 161452
rect 309744 161440 309750 161492
rect 163314 161372 163320 161424
rect 163372 161412 163378 161424
rect 250990 161412 250996 161424
rect 163372 161384 250996 161412
rect 163372 161372 163378 161384
rect 250990 161372 250996 161384
rect 251048 161372 251054 161424
rect 253474 161372 253480 161424
rect 253532 161412 253538 161424
rect 317690 161412 317696 161424
rect 253532 161384 317696 161412
rect 253532 161372 253538 161384
rect 317690 161372 317696 161384
rect 317748 161372 317754 161424
rect 121730 161304 121736 161356
rect 121788 161344 121794 161356
rect 220170 161344 220176 161356
rect 121788 161316 220176 161344
rect 121788 161304 121794 161316
rect 220170 161304 220176 161316
rect 220228 161304 220234 161356
rect 225690 161304 225696 161356
rect 225748 161344 225754 161356
rect 297174 161344 297180 161356
rect 225748 161316 297180 161344
rect 225748 161304 225754 161316
rect 297174 161304 297180 161316
rect 297232 161304 297238 161356
rect 105262 161236 105268 161288
rect 105320 161276 105326 161288
rect 207934 161276 207940 161288
rect 105320 161248 207940 161276
rect 105320 161236 105326 161248
rect 207934 161236 207940 161248
rect 207992 161236 207998 161288
rect 211890 161236 211896 161288
rect 211948 161276 211954 161288
rect 286870 161276 286876 161288
rect 211948 161248 286876 161276
rect 211948 161236 211954 161248
rect 286870 161236 286876 161248
rect 286928 161236 286934 161288
rect 90450 161168 90456 161220
rect 90508 161208 90514 161220
rect 196986 161208 196992 161220
rect 90508 161180 196992 161208
rect 90508 161168 90514 161180
rect 196986 161168 196992 161180
rect 197044 161168 197050 161220
rect 199746 161168 199752 161220
rect 199804 161208 199810 161220
rect 277946 161208 277952 161220
rect 199804 161180 277952 161208
rect 199804 161168 199810 161180
rect 277946 161168 277952 161180
rect 278004 161168 278010 161220
rect 80054 161100 80060 161152
rect 80112 161140 80118 161152
rect 189166 161140 189172 161152
rect 80112 161112 189172 161140
rect 80112 161100 80118 161112
rect 189166 161100 189172 161112
rect 189224 161100 189230 161152
rect 191006 161100 191012 161152
rect 191064 161140 191070 161152
rect 271506 161140 271512 161152
rect 191064 161112 271512 161140
rect 191064 161100 191070 161112
rect 271506 161100 271512 161112
rect 271564 161100 271570 161152
rect 66254 161032 66260 161084
rect 66312 161072 66318 161084
rect 179046 161072 179052 161084
rect 66312 161044 179052 161072
rect 66312 161032 66318 161044
rect 179046 161032 179052 161044
rect 179104 161032 179110 161084
rect 180610 161032 180616 161084
rect 180668 161072 180674 161084
rect 263778 161072 263784 161084
rect 180668 161044 263784 161072
rect 180668 161032 180674 161044
rect 263778 161032 263784 161044
rect 263836 161032 263842 161084
rect 265618 161032 265624 161084
rect 265676 161072 265682 161084
rect 326706 161072 326712 161084
rect 265676 161044 326712 161072
rect 265676 161032 265682 161044
rect 326706 161032 326712 161044
rect 326764 161032 326770 161084
rect 37642 160964 37648 161016
rect 37700 161004 37706 161016
rect 157886 161004 157892 161016
rect 37700 160976 157892 161004
rect 37700 160964 37706 160976
rect 157886 160964 157892 160976
rect 157944 160964 157950 161016
rect 166810 160964 166816 161016
rect 166868 161004 166874 161016
rect 253474 161004 253480 161016
rect 166868 160976 253480 161004
rect 166868 160964 166874 160976
rect 253474 160964 253480 160976
rect 253532 160964 253538 161016
rect 255222 160964 255228 161016
rect 255280 161004 255286 161016
rect 318978 161004 318984 161016
rect 255280 160976 318984 161004
rect 255280 160964 255286 160976
rect 318978 160964 318984 160976
rect 319036 160964 319042 161016
rect 26326 160896 26332 160948
rect 26384 160936 26390 160948
rect 149514 160936 149520 160948
rect 26384 160908 149520 160936
rect 26384 160896 26390 160908
rect 149514 160896 149520 160908
rect 149572 160896 149578 160948
rect 159818 160896 159824 160948
rect 159876 160936 159882 160948
rect 248414 160936 248420 160948
rect 159876 160908 248420 160936
rect 159876 160896 159882 160908
rect 248414 160896 248420 160908
rect 248472 160896 248478 160948
rect 249978 160896 249984 160948
rect 250036 160936 250042 160948
rect 315114 160936 315120 160948
rect 250036 160908 315120 160936
rect 250036 160896 250042 160908
rect 315114 160896 315120 160908
rect 315172 160896 315178 160948
rect 18506 160828 18512 160880
rect 18564 160868 18570 160880
rect 143718 160868 143724 160880
rect 18564 160840 143724 160868
rect 18564 160828 18570 160840
rect 143718 160828 143724 160840
rect 143776 160828 143782 160880
rect 152918 160828 152924 160880
rect 152976 160868 152982 160880
rect 243262 160868 243268 160880
rect 152976 160840 243268 160868
rect 152976 160828 152982 160840
rect 243262 160828 243268 160840
rect 243320 160828 243326 160880
rect 246482 160828 246488 160880
rect 246540 160868 246546 160880
rect 312630 160868 312636 160880
rect 246540 160840 312636 160868
rect 246540 160828 246546 160840
rect 312630 160828 312636 160840
rect 312688 160828 312694 160880
rect 11606 160760 11612 160812
rect 11664 160800 11670 160812
rect 138566 160800 138572 160812
rect 11664 160772 138572 160800
rect 11664 160760 11670 160772
rect 138566 160760 138572 160772
rect 138624 160760 138630 160812
rect 145926 160760 145932 160812
rect 145984 160800 145990 160812
rect 232501 160803 232559 160809
rect 232501 160800 232513 160803
rect 145984 160772 232513 160800
rect 145984 160760 145990 160772
rect 232501 160769 232513 160772
rect 232547 160769 232559 160803
rect 232958 160800 232964 160812
rect 232501 160763 232559 160769
rect 232608 160772 232964 160800
rect 4706 160692 4712 160744
rect 4764 160732 4770 160744
rect 133414 160732 133420 160744
rect 4764 160704 133420 160732
rect 4764 160692 4770 160704
rect 133414 160692 133420 160704
rect 133472 160692 133478 160744
rect 139026 160692 139032 160744
rect 139084 160732 139090 160744
rect 232608 160732 232636 160772
rect 232958 160760 232964 160772
rect 233016 160760 233022 160812
rect 239582 160760 239588 160812
rect 239640 160800 239646 160812
rect 307478 160800 307484 160812
rect 239640 160772 307484 160800
rect 239640 160760 239646 160772
rect 307478 160760 307484 160772
rect 307536 160760 307542 160812
rect 139084 160704 232636 160732
rect 139084 160692 139090 160704
rect 232682 160692 232688 160744
rect 232740 160732 232746 160744
rect 302326 160732 302332 160744
rect 232740 160704 302332 160732
rect 232740 160692 232746 160704
rect 302326 160692 302332 160704
rect 302384 160692 302390 160744
rect 170214 160624 170220 160676
rect 170272 160664 170278 160676
rect 255958 160664 255964 160676
rect 170272 160636 255964 160664
rect 170272 160624 170278 160636
rect 255958 160624 255964 160636
rect 256016 160624 256022 160676
rect 256878 160624 256884 160676
rect 256936 160664 256942 160676
rect 320266 160664 320272 160676
rect 256936 160636 320272 160664
rect 256936 160624 256942 160636
rect 320266 160624 320272 160636
rect 320324 160624 320330 160676
rect 173710 160556 173716 160608
rect 173768 160596 173774 160608
rect 258534 160596 258540 160608
rect 173768 160568 258540 160596
rect 173768 160556 173774 160568
rect 258534 160556 258540 160568
rect 258592 160556 258598 160608
rect 263870 160556 263876 160608
rect 263928 160596 263934 160608
rect 325326 160596 325332 160608
rect 263928 160568 325332 160596
rect 263928 160556 263934 160568
rect 325326 160556 325332 160568
rect 325384 160556 325390 160608
rect 232501 160531 232559 160537
rect 232501 160497 232513 160531
rect 232547 160528 232559 160531
rect 238110 160528 238116 160540
rect 232547 160500 238116 160528
rect 232547 160497 232559 160500
rect 232501 160491 232559 160497
rect 238110 160488 238116 160500
rect 238168 160488 238174 160540
rect 100938 160216 100944 160268
rect 100996 160256 101002 160268
rect 165522 160256 165528 160268
rect 100996 160228 165528 160256
rect 100996 160216 101002 160228
rect 165522 160216 165528 160228
rect 165580 160216 165586 160268
rect 50614 160148 50620 160200
rect 50672 160188 50678 160200
rect 167454 160188 167460 160200
rect 50672 160160 167460 160188
rect 50672 160148 50678 160160
rect 167454 160148 167460 160160
rect 167512 160148 167518 160200
rect 28902 160080 28908 160132
rect 28960 160120 28966 160132
rect 151446 160120 151452 160132
rect 28960 160092 151452 160120
rect 28960 160080 28966 160092
rect 151446 160080 151452 160092
rect 151504 160080 151510 160132
rect 138198 160012 138204 160064
rect 138256 160052 138262 160064
rect 232314 160052 232320 160064
rect 138256 160024 232320 160052
rect 138256 160012 138262 160024
rect 232314 160012 232320 160024
rect 232372 160012 232378 160064
rect 259546 160012 259552 160064
rect 259604 160052 259610 160064
rect 311894 160052 311900 160064
rect 259604 160024 311900 160052
rect 259604 160012 259610 160024
rect 311894 160012 311900 160024
rect 311952 160012 311958 160064
rect 338390 160012 338396 160064
rect 338448 160052 338454 160064
rect 376662 160052 376668 160064
rect 338448 160024 376668 160052
rect 338448 160012 338454 160024
rect 376662 160012 376668 160024
rect 376720 160012 376726 160064
rect 418154 160012 418160 160064
rect 418212 160052 418218 160064
rect 439682 160052 439688 160064
rect 418212 160024 439688 160052
rect 418212 160012 418218 160024
rect 439682 160012 439688 160024
rect 439740 160012 439746 160064
rect 452838 160012 452844 160064
rect 452896 160052 452902 160064
rect 463786 160052 463792 160064
rect 452896 160024 463792 160052
rect 452896 160012 452902 160024
rect 463786 160012 463792 160024
rect 463844 160012 463850 160064
rect 484026 160012 484032 160064
rect 484084 160012 484090 160064
rect 486602 160012 486608 160064
rect 486660 160052 486666 160064
rect 488258 160052 488264 160064
rect 486660 160024 488264 160052
rect 486660 160012 486666 160024
rect 488258 160012 488264 160024
rect 488316 160012 488322 160064
rect 61838 159944 61844 159996
rect 61896 159984 61902 159996
rect 118694 159984 118700 159996
rect 61896 159956 118700 159984
rect 61896 159944 61902 159956
rect 118694 159944 118700 159956
rect 118752 159944 118758 159996
rect 131206 159944 131212 159996
rect 131264 159984 131270 159996
rect 225046 159984 225052 159996
rect 131264 159956 225052 159984
rect 131264 159944 131270 159956
rect 225046 159944 225052 159956
rect 225104 159944 225110 159996
rect 245654 159944 245660 159996
rect 245712 159984 245718 159996
rect 301774 159984 301780 159996
rect 245712 159956 301780 159984
rect 245712 159944 245718 159956
rect 301774 159944 301780 159956
rect 301832 159944 301838 159996
rect 331490 159944 331496 159996
rect 331548 159984 331554 159996
rect 372706 159984 372712 159996
rect 331548 159956 372712 159984
rect 331548 159944 331554 159956
rect 372706 159944 372712 159956
rect 372764 159944 372770 159996
rect 408586 159944 408592 159996
rect 408644 159984 408650 159996
rect 432690 159984 432696 159996
rect 408644 159956 432696 159984
rect 408644 159944 408650 159956
rect 432690 159944 432696 159956
rect 432748 159944 432754 159996
rect 445846 159944 445852 159996
rect 445904 159984 445910 159996
rect 456886 159984 456892 159996
rect 445904 159956 456892 159984
rect 445904 159944 445910 159956
rect 456886 159944 456892 159956
rect 456944 159944 456950 159996
rect 458910 159944 458916 159996
rect 458968 159984 458974 159996
rect 469858 159984 469864 159996
rect 458968 159956 469864 159984
rect 458968 159944 458974 159956
rect 469858 159944 469864 159956
rect 469916 159944 469922 159996
rect 475378 159944 475384 159996
rect 475436 159984 475442 159996
rect 481082 159984 481088 159996
rect 475436 159956 481088 159984
rect 475436 159944 475442 159956
rect 481082 159944 481088 159956
rect 481140 159944 481146 159996
rect 484044 159984 484072 160012
rect 488718 159984 488724 159996
rect 484044 159956 488724 159984
rect 488718 159944 488724 159956
rect 488776 159944 488782 159996
rect 41046 159876 41052 159928
rect 41104 159916 41110 159928
rect 56502 159916 56508 159928
rect 41104 159888 56508 159916
rect 41104 159876 41110 159888
rect 56502 159876 56508 159888
rect 56560 159876 56566 159928
rect 89622 159876 89628 159928
rect 89680 159916 89686 159928
rect 186222 159916 186228 159928
rect 89680 159888 186228 159916
rect 89680 159876 89686 159888
rect 186222 159876 186228 159888
rect 186280 159876 186286 159928
rect 196250 159876 196256 159928
rect 196308 159916 196314 159928
rect 260558 159916 260564 159928
rect 196308 159888 260564 159916
rect 196308 159876 196314 159888
rect 260558 159876 260564 159888
rect 260616 159876 260622 159928
rect 266446 159876 266452 159928
rect 266504 159916 266510 159928
rect 316218 159916 316224 159928
rect 266504 159888 316224 159916
rect 266504 159876 266510 159888
rect 316218 159876 316224 159888
rect 316276 159876 316282 159928
rect 339310 159876 339316 159928
rect 339368 159916 339374 159928
rect 381262 159916 381268 159928
rect 339368 159888 381268 159916
rect 339368 159876 339374 159888
rect 381262 159876 381268 159888
rect 381320 159876 381326 159928
rect 394786 159876 394792 159928
rect 394844 159916 394850 159928
rect 420914 159916 420920 159928
rect 394844 159888 420920 159916
rect 394844 159876 394850 159888
rect 420914 159876 420920 159888
rect 420972 159876 420978 159928
rect 451090 159876 451096 159928
rect 451148 159916 451154 159928
rect 462130 159916 462136 159928
rect 451148 159888 462136 159916
rect 451148 159876 451154 159888
rect 462130 159876 462136 159888
rect 462188 159876 462194 159928
rect 468386 159876 468392 159928
rect 468444 159916 468450 159928
rect 468444 159888 471836 159916
rect 468444 159876 468450 159888
rect 33318 159808 33324 159860
rect 33376 159848 33382 159860
rect 49602 159848 49608 159860
rect 33376 159820 49608 159848
rect 33376 159808 33382 159820
rect 49602 159808 49608 159820
rect 49660 159808 49666 159860
rect 71406 159808 71412 159860
rect 71464 159848 71470 159860
rect 114646 159848 114652 159860
rect 71464 159820 114652 159848
rect 71464 159808 71470 159820
rect 114646 159808 114652 159820
rect 114704 159808 114710 159860
rect 119062 159808 119068 159860
rect 119120 159848 119126 159860
rect 218238 159848 218244 159860
rect 119120 159820 218244 159848
rect 119120 159808 119126 159820
rect 218238 159808 218244 159820
rect 218296 159808 218302 159860
rect 235258 159808 235264 159860
rect 235316 159848 235322 159860
rect 291838 159848 291844 159860
rect 235316 159820 291844 159848
rect 235316 159808 235322 159820
rect 291838 159808 291844 159820
rect 291896 159808 291902 159860
rect 321922 159808 321928 159860
rect 321980 159848 321986 159860
rect 366910 159848 366916 159860
rect 321980 159820 366916 159848
rect 321980 159808 321986 159820
rect 366910 159808 366916 159820
rect 366968 159808 366974 159860
rect 376570 159808 376576 159860
rect 376628 159848 376634 159860
rect 391934 159848 391940 159860
rect 376628 159820 391940 159848
rect 376628 159808 376634 159820
rect 391934 159808 391940 159820
rect 391992 159808 391998 159860
rect 393866 159808 393872 159860
rect 393924 159848 393930 159860
rect 421742 159848 421748 159860
rect 393924 159820 421748 159848
rect 393924 159808 393930 159820
rect 421742 159808 421748 159820
rect 421800 159808 421806 159860
rect 432046 159808 432052 159860
rect 432104 159848 432110 159860
rect 436002 159848 436008 159860
rect 432104 159820 436008 159848
rect 432104 159808 432110 159820
rect 436002 159808 436008 159820
rect 436060 159808 436066 159860
rect 450262 159808 450268 159860
rect 450320 159848 450326 159860
rect 462222 159848 462228 159860
rect 450320 159820 462228 159848
rect 450320 159808 450326 159820
rect 462222 159808 462228 159820
rect 462280 159808 462286 159860
rect 470134 159808 470140 159860
rect 470192 159848 470198 159860
rect 471701 159851 471759 159857
rect 471701 159848 471713 159851
rect 470192 159820 471713 159848
rect 470192 159808 470198 159820
rect 471701 159817 471713 159820
rect 471747 159817 471759 159851
rect 471808 159848 471836 159888
rect 471882 159876 471888 159928
rect 471940 159916 471946 159928
rect 476114 159916 476120 159928
rect 471940 159888 476120 159916
rect 471940 159876 471946 159888
rect 476114 159876 476120 159888
rect 476172 159876 476178 159928
rect 477954 159876 477960 159928
rect 478012 159916 478018 159928
rect 484026 159916 484032 159928
rect 478012 159888 484032 159916
rect 478012 159876 478018 159888
rect 484026 159876 484032 159888
rect 484084 159876 484090 159928
rect 473722 159848 473728 159860
rect 471808 159820 473728 159848
rect 471701 159811 471759 159817
rect 473722 159808 473728 159820
rect 473780 159808 473786 159860
rect 19426 159740 19432 159792
rect 19484 159780 19490 159792
rect 41414 159780 41420 159792
rect 19484 159752 41420 159780
rect 19484 159740 19490 159752
rect 41414 159740 41420 159752
rect 41472 159740 41478 159792
rect 47118 159740 47124 159792
rect 47176 159780 47182 159792
rect 100754 159780 100760 159792
rect 47176 159752 100760 159780
rect 47176 159740 47182 159752
rect 100754 159740 100760 159752
rect 100812 159740 100818 159792
rect 113910 159740 113916 159792
rect 113968 159780 113974 159792
rect 214282 159780 214288 159792
rect 113968 159752 214288 159780
rect 113968 159740 113974 159752
rect 214282 159740 214288 159752
rect 214340 159740 214346 159792
rect 238754 159740 238760 159792
rect 238812 159780 238818 159792
rect 296622 159780 296628 159792
rect 238812 159752 296628 159780
rect 238812 159740 238818 159752
rect 296622 159740 296628 159752
rect 296680 159740 296686 159792
rect 324498 159740 324504 159792
rect 324556 159780 324562 159792
rect 370406 159780 370412 159792
rect 324556 159752 370412 159780
rect 324556 159740 324562 159752
rect 370406 159740 370412 159752
rect 370464 159740 370470 159792
rect 380894 159740 380900 159792
rect 380952 159780 380958 159792
rect 411990 159780 411996 159792
rect 380952 159752 411996 159780
rect 380952 159740 380958 159752
rect 411990 159740 411996 159752
rect 412048 159740 412054 159792
rect 425974 159740 425980 159792
rect 426032 159780 426038 159792
rect 445478 159780 445484 159792
rect 426032 159752 445484 159780
rect 426032 159740 426038 159752
rect 445478 159740 445484 159752
rect 445536 159740 445542 159792
rect 451918 159740 451924 159792
rect 451976 159780 451982 159792
rect 462866 159780 462872 159792
rect 451976 159752 462872 159780
rect 451976 159740 451982 159752
rect 462866 159740 462872 159752
rect 462924 159740 462930 159792
rect 465810 159740 465816 159792
rect 465868 159780 465874 159792
rect 471882 159780 471888 159792
rect 465868 159752 471888 159780
rect 465868 159740 465874 159752
rect 471882 159740 471888 159752
rect 471940 159740 471946 159792
rect 478874 159740 478880 159792
rect 478932 159780 478938 159792
rect 484670 159780 484676 159792
rect 478932 159752 484676 159780
rect 478932 159740 478938 159752
rect 484670 159740 484676 159752
rect 484728 159740 484734 159792
rect 32398 159672 32404 159724
rect 32456 159712 32462 159724
rect 69658 159712 69664 159724
rect 32456 159684 69664 159712
rect 32456 159672 32462 159684
rect 69658 159672 69664 159684
rect 69716 159672 69722 159724
rect 82722 159672 82728 159724
rect 82780 159712 82786 159724
rect 183462 159712 183468 159724
rect 82780 159684 183468 159712
rect 82780 159672 82786 159684
rect 183462 159672 183468 159684
rect 183520 159672 183526 159724
rect 185854 159672 185860 159724
rect 185912 159712 185918 159724
rect 264974 159712 264980 159724
rect 185912 159684 264980 159712
rect 185912 159672 185918 159684
rect 264974 159672 264980 159684
rect 265032 159672 265038 159724
rect 273346 159672 273352 159724
rect 273404 159712 273410 159724
rect 328362 159712 328368 159724
rect 273404 159684 328368 159712
rect 273404 159672 273410 159684
rect 328362 159672 328368 159684
rect 328420 159672 328426 159724
rect 328822 159672 328828 159724
rect 328880 159712 328886 159724
rect 373626 159712 373632 159724
rect 328880 159684 373632 159712
rect 328880 159672 328886 159684
rect 373626 159672 373632 159684
rect 373684 159672 373690 159724
rect 379974 159672 379980 159724
rect 380032 159712 380038 159724
rect 411162 159712 411168 159724
rect 380032 159684 411168 159712
rect 380032 159672 380038 159684
rect 411162 159672 411168 159684
rect 411220 159672 411226 159724
rect 412082 159672 412088 159724
rect 412140 159712 412146 159724
rect 435266 159712 435272 159724
rect 412140 159684 435272 159712
rect 412140 159672 412146 159684
rect 435266 159672 435272 159684
rect 435324 159672 435330 159724
rect 448514 159672 448520 159724
rect 448572 159712 448578 159724
rect 459830 159712 459836 159724
rect 448572 159684 459836 159712
rect 448572 159672 448578 159684
rect 459830 159672 459836 159684
rect 459888 159672 459894 159724
rect 471701 159715 471759 159721
rect 471701 159681 471713 159715
rect 471747 159712 471759 159715
rect 475746 159712 475752 159724
rect 471747 159684 475752 159712
rect 471747 159681 471759 159684
rect 471701 159675 471759 159681
rect 475746 159672 475752 159684
rect 475804 159672 475810 159724
rect 22002 159604 22008 159656
rect 22060 159644 22066 159656
rect 62114 159644 62120 159656
rect 22060 159616 62120 159644
rect 22060 159604 22066 159616
rect 62114 159604 62120 159616
rect 62172 159604 62178 159656
rect 101766 159604 101772 159656
rect 101824 159644 101830 159656
rect 205358 159644 205364 159656
rect 101824 159616 205364 159644
rect 101824 159604 101830 159616
rect 205358 159604 205364 159616
rect 205416 159604 205422 159656
rect 221366 159604 221372 159656
rect 221424 159644 221430 159656
rect 280982 159644 280988 159656
rect 221424 159616 280988 159644
rect 221424 159604 221430 159616
rect 280982 159604 280988 159616
rect 281040 159604 281046 159656
rect 308030 159604 308036 159656
rect 308088 159644 308094 159656
rect 356422 159644 356428 159656
rect 308088 159616 356428 159644
rect 308088 159604 308094 159616
rect 356422 159604 356428 159616
rect 356480 159604 356486 159656
rect 367002 159604 367008 159656
rect 367060 159644 367066 159656
rect 397270 159644 397276 159656
rect 367060 159616 397276 159644
rect 367060 159604 367066 159616
rect 397270 159604 397276 159616
rect 397328 159604 397334 159656
rect 401686 159604 401692 159656
rect 401744 159644 401750 159656
rect 427538 159644 427544 159656
rect 401744 159616 427544 159644
rect 401744 159604 401750 159616
rect 427538 159604 427544 159616
rect 427596 159604 427602 159656
rect 431126 159604 431132 159656
rect 431184 159644 431190 159656
rect 437474 159644 437480 159656
rect 431184 159616 437480 159644
rect 431184 159604 431190 159616
rect 437474 159604 437480 159616
rect 437532 159604 437538 159656
rect 442442 159604 442448 159656
rect 442500 159644 442506 159656
rect 445662 159644 445668 159656
rect 442500 159616 445668 159644
rect 442500 159604 442506 159616
rect 445662 159604 445668 159616
rect 445720 159604 445726 159656
rect 447594 159604 447600 159656
rect 447652 159644 447658 159656
rect 458174 159644 458180 159656
rect 447652 159616 458180 159644
rect 447652 159604 447658 159616
rect 458174 159604 458180 159616
rect 458232 159604 458238 159656
rect 460658 159604 460664 159656
rect 460716 159644 460722 159656
rect 471146 159644 471152 159656
rect 460716 159616 471152 159644
rect 460716 159604 460722 159616
rect 471146 159604 471152 159616
rect 471204 159604 471210 159656
rect 5534 159536 5540 159588
rect 5592 159576 5598 159588
rect 28902 159576 28908 159588
rect 5592 159548 28908 159576
rect 5592 159536 5598 159548
rect 28902 159536 28908 159548
rect 28960 159536 28966 159588
rect 34974 159536 34980 159588
rect 35032 159576 35038 159588
rect 80054 159576 80060 159588
rect 35032 159548 80060 159576
rect 35032 159536 35038 159548
rect 80054 159536 80060 159548
rect 80112 159536 80118 159588
rect 100846 159536 100852 159588
rect 100904 159576 100910 159588
rect 204714 159576 204720 159588
rect 100904 159548 204720 159576
rect 100904 159536 100910 159548
rect 204714 159536 204720 159548
rect 204772 159536 204778 159588
rect 213546 159536 213552 159588
rect 213604 159576 213610 159588
rect 224954 159576 224960 159588
rect 213604 159548 224960 159576
rect 213604 159536 213610 159548
rect 224954 159536 224960 159548
rect 225012 159536 225018 159588
rect 228358 159536 228364 159588
rect 228416 159576 228422 159588
rect 289722 159576 289728 159588
rect 228416 159548 289728 159576
rect 228416 159536 228422 159548
rect 289722 159536 289728 159548
rect 289780 159536 289786 159588
rect 301130 159536 301136 159588
rect 301188 159576 301194 159588
rect 350166 159576 350172 159588
rect 301188 159548 350172 159576
rect 301188 159536 301194 159548
rect 350166 159536 350172 159548
rect 350224 159536 350230 159588
rect 353110 159536 353116 159588
rect 353168 159576 353174 159588
rect 385954 159576 385960 159588
rect 353168 159548 385960 159576
rect 353168 159536 353174 159548
rect 385954 159536 385960 159548
rect 386012 159536 386018 159588
rect 386966 159536 386972 159588
rect 387024 159576 387030 159588
rect 415210 159576 415216 159588
rect 387024 159548 415216 159576
rect 387024 159536 387030 159548
rect 415210 159536 415216 159548
rect 415268 159536 415274 159588
rect 421650 159536 421656 159588
rect 421708 159576 421714 159588
rect 442258 159576 442264 159588
rect 421708 159548 442264 159576
rect 421708 159536 421714 159548
rect 442258 159536 442264 159548
rect 442316 159536 442322 159588
rect 449342 159536 449348 159588
rect 449400 159576 449406 159588
rect 449400 159548 451274 159576
rect 449400 159536 449406 159548
rect 1210 159468 1216 159520
rect 1268 159508 1274 159520
rect 89714 159508 89720 159520
rect 1268 159480 89720 159508
rect 1268 159468 1274 159480
rect 89714 159468 89720 159480
rect 89772 159468 89778 159520
rect 91370 159468 91376 159520
rect 91428 159508 91434 159520
rect 99374 159508 99380 159520
rect 91428 159480 99380 159508
rect 91428 159468 91434 159480
rect 99374 159468 99380 159480
rect 99432 159468 99438 159520
rect 104342 159468 104348 159520
rect 104400 159508 104406 159520
rect 207290 159508 207296 159520
rect 104400 159480 207296 159508
rect 104400 159468 104406 159480
rect 207290 159468 207296 159480
rect 207348 159468 207354 159520
rect 210142 159468 210148 159520
rect 210200 159508 210206 159520
rect 276106 159508 276112 159520
rect 210200 159480 276112 159508
rect 210200 159468 210206 159480
rect 276106 159468 276112 159480
rect 276164 159468 276170 159520
rect 294230 159468 294236 159520
rect 294288 159508 294294 159520
rect 347682 159508 347688 159520
rect 294288 159480 347688 159508
rect 294288 159468 294294 159480
rect 347682 159468 347688 159480
rect 347740 159468 347746 159520
rect 360102 159468 360108 159520
rect 360160 159508 360166 159520
rect 396718 159508 396724 159520
rect 360160 159480 396724 159508
rect 360160 159468 360166 159480
rect 396718 159468 396724 159480
rect 396776 159468 396782 159520
rect 400858 159468 400864 159520
rect 400916 159508 400922 159520
rect 426894 159508 426900 159520
rect 400916 159480 426900 159508
rect 400916 159468 400922 159480
rect 426894 159468 426900 159480
rect 426952 159468 426958 159520
rect 429378 159468 429384 159520
rect 429436 159508 429442 159520
rect 446858 159508 446864 159520
rect 429436 159480 446864 159508
rect 429436 159468 429442 159480
rect 446858 159468 446864 159480
rect 446916 159468 446922 159520
rect 451246 159508 451274 159548
rect 457990 159536 457996 159588
rect 458048 159576 458054 159588
rect 469122 159576 469128 159588
rect 458048 159548 469128 159576
rect 458048 159536 458054 159548
rect 469122 159536 469128 159548
rect 469180 159536 469186 159588
rect 469306 159536 469312 159588
rect 469364 159576 469370 159588
rect 474734 159576 474740 159588
rect 469364 159548 474740 159576
rect 469364 159536 469370 159548
rect 474734 159536 474740 159548
rect 474792 159536 474798 159588
rect 459554 159508 459560 159520
rect 451246 159480 459560 159508
rect 459554 159468 459560 159480
rect 459612 159468 459618 159520
rect 462406 159468 462412 159520
rect 462464 159508 462470 159520
rect 468202 159508 468208 159520
rect 462464 159480 468208 159508
rect 462464 159468 462470 159480
rect 468202 159468 468208 159480
rect 468260 159468 468266 159520
rect 479702 159468 479708 159520
rect 479760 159508 479766 159520
rect 485314 159508 485320 159520
rect 479760 159480 485320 159508
rect 479760 159468 479766 159480
rect 485314 159468 485320 159480
rect 485372 159468 485378 159520
rect 382 159400 388 159452
rect 440 159440 446 159452
rect 39942 159440 39948 159452
rect 440 159412 39948 159440
rect 440 159400 446 159412
rect 39942 159400 39948 159412
rect 40000 159400 40006 159452
rect 45370 159400 45376 159452
rect 45428 159440 45434 159452
rect 154390 159440 154396 159452
rect 45428 159412 154396 159440
rect 45428 159400 45434 159412
rect 154390 159400 154396 159412
rect 154448 159400 154454 159452
rect 162394 159400 162400 159452
rect 162452 159440 162458 159452
rect 245654 159440 245660 159452
rect 162452 159412 245660 159440
rect 162452 159400 162458 159412
rect 245654 159400 245660 159412
rect 245712 159400 245718 159452
rect 258626 159400 258632 159452
rect 258684 159440 258690 159452
rect 282178 159440 282184 159452
rect 258684 159412 282184 159440
rect 258684 159400 258690 159412
rect 282178 159400 282184 159412
rect 282236 159400 282242 159452
rect 342714 159400 342720 159452
rect 342772 159440 342778 159452
rect 382274 159440 382280 159452
rect 342772 159412 382280 159440
rect 342772 159400 342778 159412
rect 382274 159400 382280 159412
rect 382332 159400 382338 159452
rect 387794 159400 387800 159452
rect 387852 159440 387858 159452
rect 417234 159440 417240 159452
rect 387852 159412 417240 159440
rect 387852 159400 387858 159412
rect 417234 159400 417240 159412
rect 417292 159400 417298 159452
rect 439866 159400 439872 159452
rect 439924 159440 439930 159452
rect 446398 159440 446404 159452
rect 439924 159412 446404 159440
rect 439924 159400 439930 159412
rect 446398 159400 446404 159412
rect 446456 159400 446462 159452
rect 454586 159400 454592 159452
rect 454644 159440 454650 159452
rect 466362 159440 466368 159452
rect 454644 159412 466368 159440
rect 454644 159400 454650 159412
rect 466362 159400 466368 159412
rect 466420 159400 466426 159452
rect 3786 159332 3792 159384
rect 3844 159372 3850 159384
rect 34514 159372 34520 159384
rect 3844 159344 34520 159372
rect 3844 159332 3850 159344
rect 34514 159332 34520 159344
rect 34572 159332 34578 159384
rect 38470 159332 38476 159384
rect 38528 159372 38534 159384
rect 154482 159372 154488 159384
rect 38528 159344 154488 159372
rect 38528 159332 38534 159344
rect 154482 159332 154488 159344
rect 154540 159332 154546 159384
rect 155494 159332 155500 159384
rect 155552 159372 155558 159384
rect 245194 159372 245200 159384
rect 155552 159344 245200 159372
rect 155552 159332 155558 159344
rect 245194 159332 245200 159344
rect 245252 159332 245258 159384
rect 252554 159332 252560 159384
rect 252612 159372 252618 159384
rect 310238 159372 310244 159384
rect 252612 159344 310244 159372
rect 252612 159332 252618 159344
rect 310238 159332 310244 159344
rect 310296 159332 310302 159384
rect 315022 159332 315028 159384
rect 315080 159372 315086 159384
rect 363322 159372 363328 159384
rect 315080 159344 363328 159372
rect 315080 159332 315086 159344
rect 363322 159332 363328 159344
rect 363380 159332 363386 159384
rect 373902 159332 373908 159384
rect 373960 159372 373966 159384
rect 406746 159372 406752 159384
rect 373960 159344 406752 159372
rect 373960 159332 373966 159344
rect 406746 159332 406752 159344
rect 406804 159332 406810 159384
rect 407758 159332 407764 159384
rect 407816 159372 407822 159384
rect 432046 159372 432052 159384
rect 407816 159344 432052 159372
rect 407816 159332 407822 159344
rect 432046 159332 432052 159344
rect 432104 159332 432110 159384
rect 453666 159332 453672 159384
rect 453724 159372 453730 159384
rect 463694 159372 463700 159384
rect 453724 159344 463700 159372
rect 453724 159332 453730 159344
rect 463694 159332 463700 159344
rect 463752 159332 463758 159384
rect 473630 159332 473636 159384
rect 473688 159372 473694 159384
rect 478966 159372 478972 159384
rect 473688 159344 478972 159372
rect 473688 159332 473694 159344
rect 478966 159332 478972 159344
rect 479024 159332 479030 159384
rect 48038 159264 48044 159316
rect 48096 159304 48102 159316
rect 100938 159304 100944 159316
rect 48096 159276 100944 159304
rect 48096 159264 48102 159276
rect 100938 159264 100944 159276
rect 100996 159264 101002 159316
rect 106918 159264 106924 159316
rect 106976 159304 106982 159316
rect 198734 159304 198740 159316
rect 106976 159276 198740 159304
rect 106976 159264 106982 159276
rect 198734 159264 198740 159276
rect 198792 159264 198798 159316
rect 244826 159264 244832 159316
rect 244884 159304 244890 159316
rect 272426 159304 272432 159316
rect 244884 159276 272432 159304
rect 244884 159264 244890 159276
rect 272426 159264 272432 159276
rect 272484 159264 272490 159316
rect 276014 159264 276020 159316
rect 276072 159304 276078 159316
rect 293954 159304 293960 159316
rect 276072 159276 293960 159304
rect 276072 159264 276078 159276
rect 293954 159264 293960 159276
rect 294012 159264 294018 159316
rect 296806 159264 296812 159316
rect 296864 159304 296870 159316
rect 332594 159304 332600 159316
rect 296864 159276 332600 159304
rect 296864 159264 296870 159276
rect 332594 159264 332600 159276
rect 332652 159264 332658 159316
rect 345382 159264 345388 159316
rect 345440 159304 345446 159316
rect 379514 159304 379520 159316
rect 345440 159276 379520 159304
rect 345440 159264 345446 159276
rect 379514 159264 379520 159276
rect 379572 159264 379578 159316
rect 456334 159264 456340 159316
rect 456392 159304 456398 159316
rect 467742 159304 467748 159316
rect 456392 159276 467748 159304
rect 456392 159264 456398 159276
rect 467742 159264 467748 159276
rect 467800 159264 467806 159316
rect 99190 159196 99196 159248
rect 99248 159236 99254 159248
rect 138014 159236 138020 159248
rect 99248 159208 138020 159236
rect 99248 159196 99254 159208
rect 138014 159196 138020 159208
rect 138072 159196 138078 159248
rect 148594 159196 148600 159248
rect 148652 159236 148658 159248
rect 238662 159236 238668 159248
rect 148652 159208 238668 159236
rect 148652 159196 148658 159208
rect 238662 159196 238668 159208
rect 238720 159196 238726 159248
rect 269022 159196 269028 159248
rect 269080 159236 269086 159248
rect 291102 159236 291108 159248
rect 269080 159208 291108 159236
rect 269080 159196 269086 159208
rect 291102 159196 291108 159208
rect 291160 159196 291166 159248
rect 303706 159196 303712 159248
rect 303764 159236 303770 159248
rect 339402 159236 339408 159248
rect 303764 159208 339408 159236
rect 303764 159196 303770 159208
rect 339402 159196 339408 159208
rect 339460 159196 339466 159248
rect 349706 159196 349712 159248
rect 349764 159236 349770 159248
rect 360194 159236 360200 159248
rect 349764 159208 360200 159236
rect 349764 159196 349770 159208
rect 360194 159196 360200 159208
rect 360252 159196 360258 159248
rect 373074 159196 373080 159248
rect 373132 159236 373138 159248
rect 388438 159236 388444 159248
rect 373132 159208 388444 159236
rect 373132 159196 373138 159208
rect 388438 159196 388444 159208
rect 388496 159196 388502 159248
rect 455414 159196 455420 159248
rect 455472 159236 455478 159248
rect 467374 159236 467380 159248
rect 455472 159208 467380 159236
rect 455472 159196 455478 159208
rect 467374 159196 467380 159208
rect 467432 159196 467438 159248
rect 12434 159128 12440 159180
rect 12492 159168 12498 159180
rect 13814 159168 13820 159180
rect 12492 159140 13820 159168
rect 12492 159128 12498 159140
rect 13814 159128 13820 159140
rect 13872 159128 13878 159180
rect 251726 159128 251732 159180
rect 251784 159168 251790 159180
rect 272058 159168 272064 159180
rect 251784 159140 272064 159168
rect 251784 159128 251790 159140
rect 272058 159128 272064 159140
rect 272116 159128 272122 159180
rect 289814 159128 289820 159180
rect 289872 159168 289878 159180
rect 308306 159168 308312 159180
rect 289872 159140 308312 159168
rect 289872 159128 289878 159140
rect 308306 159128 308312 159140
rect 308364 159128 308370 159180
rect 310698 159128 310704 159180
rect 310756 159168 310762 159180
rect 346302 159168 346308 159180
rect 310756 159140 346308 159168
rect 310756 159128 310762 159140
rect 346302 159128 346308 159140
rect 346360 159128 346366 159180
rect 366174 159128 366180 159180
rect 366232 159168 366238 159180
rect 378042 159168 378048 159180
rect 366232 159140 378048 159168
rect 366232 159128 366238 159140
rect 378042 159128 378048 159140
rect 378100 159128 378106 159180
rect 457162 159128 457168 159180
rect 457220 159168 457226 159180
rect 468662 159168 468668 159180
rect 457220 159140 468668 159168
rect 457220 159128 457226 159140
rect 468662 159128 468668 159140
rect 468720 159128 468726 159180
rect 234338 159060 234344 159112
rect 234396 159100 234402 159112
rect 253198 159100 253204 159112
rect 234396 159072 253204 159100
rect 234396 159060 234402 159072
rect 253198 159060 253204 159072
rect 253256 159060 253262 159112
rect 272518 159060 272524 159112
rect 272576 159100 272582 159112
rect 283006 159100 283012 159112
rect 272576 159072 283012 159100
rect 272576 159060 272582 159072
rect 283006 159060 283012 159072
rect 283064 159060 283070 159112
rect 293310 159060 293316 159112
rect 293368 159100 293374 159112
rect 322934 159100 322940 159112
rect 293368 159072 322940 159100
rect 293368 159060 293374 159072
rect 322934 159060 322940 159072
rect 322992 159060 322998 159112
rect 444190 159060 444196 159112
rect 444248 159100 444254 159112
rect 447226 159100 447232 159112
rect 444248 159072 447232 159100
rect 444248 159060 444254 159072
rect 447226 159060 447232 159072
rect 447284 159060 447290 159112
rect 464062 159060 464068 159112
rect 464120 159100 464126 159112
rect 469306 159100 469312 159112
rect 464120 159072 469312 159100
rect 464120 159060 464126 159072
rect 469306 159060 469312 159072
rect 469364 159060 469370 159112
rect 474458 159060 474464 159112
rect 474516 159100 474522 159112
rect 478874 159100 478880 159112
rect 474516 159072 478880 159100
rect 474516 159060 474522 159072
rect 478874 159060 478880 159072
rect 478932 159060 478938 159112
rect 223942 158992 223948 159044
rect 224000 159032 224006 159044
rect 231762 159032 231768 159044
rect 224000 159004 231768 159032
rect 224000 158992 224006 159004
rect 231762 158992 231768 159004
rect 231820 158992 231826 159044
rect 248230 158992 248236 159044
rect 248288 159032 248294 159044
rect 251082 159032 251088 159044
rect 248288 159004 251088 159032
rect 248288 158992 248294 159004
rect 251082 158992 251088 159004
rect 251140 158992 251146 159044
rect 282914 158992 282920 159044
rect 282972 159032 282978 159044
rect 311066 159032 311072 159044
rect 282972 159004 311072 159032
rect 282972 158992 282978 159004
rect 311066 158992 311072 159004
rect 311124 158992 311130 159044
rect 317598 158992 317604 159044
rect 317656 159032 317662 159044
rect 342254 159032 342260 159044
rect 317656 159004 342260 159032
rect 317656 158992 317662 159004
rect 342254 158992 342260 159004
rect 342312 158992 342318 159044
rect 384390 158992 384396 159044
rect 384448 159032 384454 159044
rect 390554 159032 390560 159044
rect 384448 159004 390560 159032
rect 384448 158992 384454 159004
rect 390554 158992 390560 159004
rect 390612 158992 390618 159044
rect 459738 158992 459744 159044
rect 459796 159032 459802 159044
rect 465626 159032 465632 159044
rect 459796 159004 465632 159032
rect 459796 158992 459802 159004
rect 465626 158992 465632 159004
rect 465684 158992 465690 159044
rect 471054 158992 471060 159044
rect 471112 159032 471118 159044
rect 476390 159032 476396 159044
rect 471112 159004 476396 159032
rect 471112 158992 471118 159004
rect 476390 158992 476396 159004
rect 476448 158992 476454 159044
rect 480530 158992 480536 159044
rect 480588 159032 480594 159044
rect 485958 159032 485964 159044
rect 480588 159004 485964 159032
rect 480588 158992 480594 159004
rect 485958 158992 485964 159004
rect 486016 158992 486022 159044
rect 287238 158924 287244 158976
rect 287296 158964 287302 158976
rect 342806 158964 342812 158976
rect 287296 158936 342812 158964
rect 287296 158924 287302 158936
rect 342806 158924 342812 158936
rect 342864 158924 342870 158976
rect 435450 158924 435456 158976
rect 435508 158964 435514 158976
rect 442810 158964 442816 158976
rect 435508 158936 442816 158964
rect 435508 158924 435514 158936
rect 442810 158924 442816 158936
rect 442868 158924 442874 158976
rect 466730 158924 466736 158976
rect 466788 158964 466794 158976
rect 473262 158964 473268 158976
rect 466788 158936 473268 158964
rect 466788 158924 466794 158936
rect 473262 158924 473268 158936
rect 473320 158924 473326 158976
rect 481450 158924 481456 158976
rect 481508 158964 481514 158976
rect 486602 158964 486608 158976
rect 481508 158936 486608 158964
rect 481508 158924 481514 158936
rect 486602 158924 486608 158936
rect 486660 158924 486666 158976
rect 487522 158924 487528 158976
rect 487580 158964 487586 158976
rect 488626 158964 488632 158976
rect 487580 158936 488632 158964
rect 487580 158924 487586 158936
rect 488626 158924 488632 158936
rect 488684 158924 488690 158976
rect 507118 158924 507124 158976
rect 507176 158964 507182 158976
rect 509142 158964 509148 158976
rect 507176 158936 509148 158964
rect 507176 158924 507182 158936
rect 509142 158924 509148 158936
rect 509200 158924 509206 158976
rect 509694 158924 509700 158976
rect 509752 158964 509758 158976
rect 512638 158964 512644 158976
rect 509752 158936 512644 158964
rect 509752 158924 509758 158936
rect 512638 158924 512644 158936
rect 512696 158924 512702 158976
rect 533154 158924 533160 158976
rect 533212 158964 533218 158976
rect 537754 158964 537760 158976
rect 533212 158936 537760 158964
rect 533212 158924 533218 158936
rect 537754 158924 537760 158936
rect 537812 158924 537818 158976
rect 237834 158856 237840 158908
rect 237892 158896 237898 158908
rect 240042 158896 240048 158908
rect 237892 158868 240048 158896
rect 237892 158856 237898 158868
rect 240042 158856 240048 158868
rect 240100 158856 240106 158908
rect 463234 158856 463240 158908
rect 463292 158896 463298 158908
rect 468110 158896 468116 158908
rect 463292 158868 468116 158896
rect 463292 158856 463298 158868
rect 468110 158856 468116 158868
rect 468168 158856 468174 158908
rect 472802 158856 472808 158908
rect 472860 158896 472866 158908
rect 477494 158896 477500 158908
rect 472860 158868 477500 158896
rect 472860 158856 472866 158868
rect 477494 158856 477500 158868
rect 477552 158856 477558 158908
rect 482278 158856 482284 158908
rect 482336 158896 482342 158908
rect 487246 158896 487252 158908
rect 482336 158868 487252 158896
rect 482336 158856 482342 158868
rect 487246 158856 487252 158868
rect 487304 158856 487310 158908
rect 489270 158856 489276 158908
rect 489328 158896 489334 158908
rect 491202 158896 491208 158908
rect 489328 158868 491208 158896
rect 489328 158856 489334 158868
rect 491202 158856 491208 158868
rect 491260 158856 491266 158908
rect 492674 158856 492680 158908
rect 492732 158896 492738 158908
rect 494974 158896 494980 158908
rect 492732 158868 494980 158896
rect 492732 158856 492738 158868
rect 494974 158856 494980 158868
rect 495032 158856 495038 158908
rect 506474 158856 506480 158908
rect 506532 158896 506538 158908
rect 508314 158896 508320 158908
rect 506532 158868 508320 158896
rect 506532 158856 506538 158868
rect 508314 158856 508320 158868
rect 508372 158856 508378 158908
rect 508406 158856 508412 158908
rect 508464 158896 508470 158908
rect 510890 158896 510896 158908
rect 508464 158868 510896 158896
rect 508464 158856 508470 158868
rect 510890 158856 510896 158868
rect 510948 158856 510954 158908
rect 532694 158856 532700 158908
rect 532752 158896 532758 158908
rect 535178 158896 535184 158908
rect 532752 158868 535184 158896
rect 532752 158856 532758 158868
rect 535178 158856 535184 158868
rect 535236 158856 535242 158908
rect 94866 158788 94872 158840
rect 94924 158828 94930 158840
rect 97810 158828 97816 158840
rect 94924 158800 97816 158828
rect 94924 158788 94930 158800
rect 97810 158788 97816 158800
rect 97868 158788 97874 158840
rect 318426 158788 318432 158840
rect 318484 158828 318490 158840
rect 324314 158828 324320 158840
rect 318484 158800 324320 158828
rect 318484 158788 318490 158800
rect 324314 158788 324320 158800
rect 324372 158788 324378 158840
rect 377398 158788 377404 158840
rect 377456 158828 377462 158840
rect 379422 158828 379428 158840
rect 377456 158800 379428 158828
rect 377456 158788 377462 158800
rect 379422 158788 379428 158800
rect 379480 158788 379486 158840
rect 398190 158788 398196 158840
rect 398248 158828 398254 158840
rect 399386 158828 399392 158840
rect 398248 158800 399392 158828
rect 398248 158788 398254 158800
rect 399386 158788 399392 158800
rect 399444 158788 399450 158840
rect 403434 158788 403440 158840
rect 403492 158828 403498 158840
rect 405642 158828 405648 158840
rect 403492 158800 405648 158828
rect 403492 158788 403498 158800
rect 405642 158788 405648 158800
rect 405700 158788 405706 158840
rect 426802 158788 426808 158840
rect 426860 158828 426866 158840
rect 429378 158828 429384 158840
rect 426860 158800 429384 158828
rect 426860 158788 426866 158800
rect 429378 158788 429384 158800
rect 429436 158788 429442 158840
rect 446766 158788 446772 158840
rect 446824 158828 446830 158840
rect 451734 158828 451740 158840
rect 446824 158800 451740 158828
rect 446824 158788 446830 158800
rect 451734 158788 451740 158800
rect 451792 158788 451798 158840
rect 461486 158788 461492 158840
rect 461544 158828 461550 158840
rect 466822 158828 466828 158840
rect 461544 158800 466828 158828
rect 461544 158788 461550 158800
rect 466822 158788 466828 158800
rect 466880 158788 466886 158840
rect 467558 158788 467564 158840
rect 467616 158828 467622 158840
rect 473170 158828 473176 158840
rect 467616 158800 473176 158828
rect 467616 158788 467622 158800
rect 473170 158788 473176 158800
rect 473228 158788 473234 158840
rect 477126 158788 477132 158840
rect 477184 158828 477190 158840
rect 482002 158828 482008 158840
rect 477184 158800 482008 158828
rect 477184 158788 477190 158800
rect 482002 158788 482008 158800
rect 482060 158788 482066 158840
rect 484854 158788 484860 158840
rect 484912 158828 484918 158840
rect 486970 158828 486976 158840
rect 484912 158800 486976 158828
rect 484912 158788 484918 158800
rect 486970 158788 486976 158800
rect 487028 158788 487034 158840
rect 491846 158788 491852 158840
rect 491904 158828 491910 158840
rect 493962 158828 493968 158840
rect 491904 158800 493968 158828
rect 491904 158788 491910 158800
rect 493962 158788 493968 158800
rect 494020 158788 494026 158840
rect 494422 158788 494428 158840
rect 494480 158828 494486 158840
rect 496262 158828 496268 158840
rect 494480 158800 496268 158828
rect 494480 158788 494486 158800
rect 496262 158788 496268 158800
rect 496320 158788 496326 158840
rect 496998 158788 497004 158840
rect 497056 158828 497062 158840
rect 498194 158828 498200 158840
rect 497056 158800 498200 158828
rect 497056 158788 497062 158800
rect 498194 158788 498200 158800
rect 498252 158788 498258 158840
rect 504542 158788 504548 158840
rect 504600 158828 504606 158840
rect 505738 158828 505744 158840
rect 504600 158800 505744 158828
rect 504600 158788 504606 158800
rect 505738 158788 505744 158800
rect 505796 158788 505802 158840
rect 505830 158788 505836 158840
rect 505888 158828 505894 158840
rect 507394 158828 507400 158840
rect 505888 158800 507400 158828
rect 505888 158788 505894 158800
rect 507394 158788 507400 158800
rect 507452 158788 507458 158840
rect 507762 158788 507768 158840
rect 507820 158828 507826 158840
rect 510062 158828 510068 158840
rect 507820 158800 510068 158828
rect 507820 158788 507826 158800
rect 510062 158788 510068 158800
rect 510120 158788 510126 158840
rect 510982 158788 510988 158840
rect 511040 158828 511046 158840
rect 514386 158828 514392 158840
rect 511040 158800 514392 158828
rect 511040 158788 511046 158800
rect 514386 158788 514392 158800
rect 514444 158788 514450 158840
rect 520550 158788 520556 158840
rect 520608 158828 520614 158840
rect 522206 158828 522212 158840
rect 520608 158800 522212 158828
rect 520608 158788 520614 158800
rect 522206 158788 522212 158800
rect 522264 158788 522270 158840
rect 523126 158788 523132 158840
rect 523184 158828 523190 158840
rect 525610 158828 525616 158840
rect 523184 158800 525616 158828
rect 523184 158788 523190 158800
rect 525610 158788 525616 158800
rect 525668 158788 525674 158840
rect 532786 158788 532792 158840
rect 532844 158828 532850 158840
rect 536926 158828 536932 158840
rect 532844 158800 536932 158828
rect 532844 158788 532850 158800
rect 536926 158788 536932 158800
rect 536984 158788 536990 158840
rect 41966 158720 41972 158772
rect 42024 158760 42030 158772
rect 46382 158760 46388 158772
rect 42024 158732 46388 158760
rect 42024 158720 42030 158732
rect 46382 158720 46388 158732
rect 46440 158720 46446 158772
rect 142522 158720 142528 158772
rect 142580 158760 142586 158772
rect 143258 158760 143264 158772
rect 142580 158732 143264 158760
rect 142580 158720 142586 158732
rect 143258 158720 143264 158732
rect 143316 158720 143322 158772
rect 172882 158720 172888 158772
rect 172940 158760 172946 158772
rect 173342 158760 173348 158772
rect 172940 158732 173348 158760
rect 172940 158720 172946 158732
rect 173342 158720 173348 158732
rect 173400 158720 173406 158772
rect 186682 158720 186688 158772
rect 186740 158760 186746 158772
rect 187602 158760 187608 158772
rect 186740 158732 187608 158760
rect 186740 158720 186746 158732
rect 187602 158720 187608 158732
rect 187660 158720 187666 158772
rect 212718 158720 212724 158772
rect 212776 158760 212782 158772
rect 213638 158760 213644 158772
rect 212776 158732 213644 158760
rect 212776 158720 212782 158732
rect 213638 158720 213644 158732
rect 213696 158720 213702 158772
rect 214466 158720 214472 158772
rect 214524 158760 214530 158772
rect 215110 158760 215116 158772
rect 214524 158732 215116 158760
rect 214524 158720 214530 158732
rect 215110 158720 215116 158732
rect 215168 158720 215174 158772
rect 230934 158720 230940 158772
rect 230992 158760 230998 158772
rect 230992 158732 234660 158760
rect 230992 158720 230998 158732
rect 127802 158652 127808 158704
rect 127860 158692 127866 158704
rect 224586 158692 224592 158704
rect 127860 158664 224592 158692
rect 127860 158652 127866 158664
rect 224586 158652 224592 158664
rect 224644 158652 224650 158704
rect 234632 158692 234660 158732
rect 247402 158720 247408 158772
rect 247460 158760 247466 158772
rect 247954 158760 247960 158772
rect 247460 158732 247960 158760
rect 247460 158720 247466 158732
rect 247954 158720 247960 158732
rect 248012 158720 248018 158772
rect 261294 158720 261300 158772
rect 261352 158760 261358 158772
rect 261938 158760 261944 158772
rect 261352 158732 261944 158760
rect 261352 158720 261358 158732
rect 261938 158720 261944 158732
rect 261996 158720 262002 158772
rect 290734 158720 290740 158772
rect 290792 158760 290798 158772
rect 292758 158760 292764 158772
rect 290792 158732 292764 158760
rect 290792 158720 290798 158732
rect 292758 158720 292764 158732
rect 292816 158720 292822 158772
rect 307202 158720 307208 158772
rect 307260 158760 307266 158772
rect 308858 158760 308864 158772
rect 307260 158732 308864 158760
rect 307260 158720 307266 158732
rect 308858 158720 308864 158732
rect 308916 158720 308922 158772
rect 311526 158720 311532 158772
rect 311584 158760 311590 158772
rect 313734 158760 313740 158772
rect 311584 158732 313740 158760
rect 311584 158720 311590 158732
rect 313734 158720 313740 158732
rect 313792 158720 313798 158772
rect 314102 158720 314108 158772
rect 314160 158760 314166 158772
rect 318702 158760 318708 158772
rect 314160 158732 318708 158760
rect 314160 158720 314166 158732
rect 318702 158720 318708 158732
rect 318760 158720 318766 158772
rect 321094 158720 321100 158772
rect 321152 158760 321158 158772
rect 321738 158760 321744 158772
rect 321152 158732 321744 158760
rect 321152 158720 321158 158732
rect 321738 158720 321744 158732
rect 321796 158720 321802 158772
rect 327994 158720 328000 158772
rect 328052 158760 328058 158772
rect 330754 158760 330760 158772
rect 328052 158732 330760 158760
rect 328052 158720 328058 158732
rect 330754 158720 330760 158732
rect 330812 158720 330818 158772
rect 346210 158720 346216 158772
rect 346268 158760 346274 158772
rect 352466 158760 352472 158772
rect 346268 158732 352472 158760
rect 346268 158720 346274 158732
rect 352466 158720 352472 158732
rect 352524 158720 352530 158772
rect 363506 158720 363512 158772
rect 363564 158760 363570 158772
rect 366266 158760 366272 158772
rect 363564 158732 366272 158760
rect 363564 158720 363570 158732
rect 366266 158720 366272 158732
rect 366324 158720 366330 158772
rect 382642 158720 382648 158772
rect 382700 158760 382706 158772
rect 384206 158760 384212 158772
rect 382700 158732 384212 158760
rect 382700 158720 382706 158732
rect 384206 158720 384212 158732
rect 384264 158720 384270 158772
rect 396442 158720 396448 158772
rect 396500 158760 396506 158772
rect 396500 158732 397500 158760
rect 396500 158720 396506 158732
rect 301038 158692 301044 158704
rect 234632 158664 301044 158692
rect 301038 158652 301044 158664
rect 301096 158652 301102 158704
rect 312354 158652 312360 158704
rect 312412 158692 312418 158704
rect 361390 158692 361396 158704
rect 312412 158664 361396 158692
rect 312412 158652 312418 158664
rect 361390 158652 361396 158664
rect 361448 158652 361454 158704
rect 397472 158692 397500 158732
rect 427722 158720 427728 158772
rect 427780 158760 427786 158772
rect 430574 158760 430580 158772
rect 427780 158732 430580 158760
rect 427780 158720 427786 158732
rect 430574 158720 430580 158732
rect 430632 158720 430638 158772
rect 445018 158720 445024 158772
rect 445076 158760 445082 158772
rect 447134 158760 447140 158772
rect 445076 158732 447140 158760
rect 445076 158720 445082 158732
rect 447134 158720 447140 158732
rect 447192 158720 447198 158772
rect 464982 158720 464988 158772
rect 465040 158760 465046 158772
rect 469214 158760 469220 158772
rect 465040 158732 469220 158760
rect 465040 158720 465046 158732
rect 469214 158720 469220 158732
rect 469272 158720 469278 158772
rect 476206 158720 476212 158772
rect 476264 158760 476270 158772
rect 482738 158760 482744 158772
rect 476264 158732 482744 158760
rect 476264 158720 476270 158732
rect 482738 158720 482744 158732
rect 482796 158720 482802 158772
rect 483198 158720 483204 158772
rect 483256 158760 483262 158772
rect 485498 158760 485504 158772
rect 483256 158732 485504 158760
rect 483256 158720 483262 158732
rect 485498 158720 485504 158732
rect 485556 158720 485562 158772
rect 485774 158720 485780 158772
rect 485832 158760 485838 158772
rect 487798 158760 487804 158772
rect 485832 158732 487804 158760
rect 485832 158720 485838 158732
rect 487798 158720 487804 158732
rect 487856 158720 487862 158772
rect 490098 158720 490104 158772
rect 490156 158760 490162 158772
rect 491570 158760 491576 158772
rect 490156 158732 491576 158760
rect 490156 158720 490162 158732
rect 491570 158720 491576 158732
rect 491628 158720 491634 158772
rect 493594 158720 493600 158772
rect 493652 158760 493658 158772
rect 495250 158760 495256 158772
rect 493652 158732 495256 158760
rect 493652 158720 493658 158732
rect 495250 158720 495256 158732
rect 495308 158720 495314 158772
rect 496170 158720 496176 158772
rect 496228 158760 496234 158772
rect 497550 158760 497556 158772
rect 496228 158732 497556 158760
rect 496228 158720 496234 158732
rect 497550 158720 497556 158732
rect 497608 158720 497614 158772
rect 497918 158720 497924 158772
rect 497976 158760 497982 158772
rect 498838 158760 498844 158772
rect 497976 158732 498844 158760
rect 497976 158720 497982 158732
rect 498838 158720 498844 158732
rect 498896 158720 498902 158772
rect 503254 158720 503260 158772
rect 503312 158760 503318 158772
rect 503714 158760 503720 158772
rect 503312 158732 503720 158760
rect 503312 158720 503318 158732
rect 503714 158720 503720 158732
rect 503772 158720 503778 158772
rect 503898 158720 503904 158772
rect 503956 158760 503962 158772
rect 504818 158760 504824 158772
rect 503956 158732 504824 158760
rect 503956 158720 503962 158732
rect 504818 158720 504824 158732
rect 504876 158720 504882 158772
rect 505186 158720 505192 158772
rect 505244 158760 505250 158772
rect 506566 158760 506572 158772
rect 505244 158732 506572 158760
rect 505244 158720 505250 158732
rect 506566 158720 506572 158732
rect 506624 158720 506630 158772
rect 509050 158720 509056 158772
rect 509108 158760 509114 158772
rect 511810 158760 511816 158772
rect 509108 158732 511816 158760
rect 509108 158720 509114 158732
rect 511810 158720 511816 158732
rect 511868 158720 511874 158772
rect 521654 158720 521660 158772
rect 521712 158760 521718 158772
rect 523862 158760 523868 158772
rect 521712 158732 523868 158760
rect 521712 158720 521718 158732
rect 523862 158720 523868 158732
rect 523920 158720 523926 158772
rect 527174 158720 527180 158772
rect 527232 158760 527238 158772
rect 530854 158760 530860 158772
rect 527232 158732 530860 158760
rect 527232 158720 527238 158732
rect 530854 158720 530860 158732
rect 530912 158720 530918 158772
rect 531406 158720 531412 158772
rect 531464 158760 531470 158772
rect 533430 158760 533436 158772
rect 531464 158732 533436 158760
rect 531464 158720 531470 158732
rect 533430 158720 533436 158732
rect 533488 158720 533494 158772
rect 538674 158760 538680 158772
rect 538635 158732 538680 158760
rect 538674 158720 538680 158732
rect 538732 158720 538738 158772
rect 539502 158760 539508 158772
rect 539463 158732 539508 158760
rect 539502 158720 539508 158732
rect 539560 158720 539566 158772
rect 397472 158664 402974 158692
rect 34514 158584 34520 158636
rect 34572 158624 34578 158636
rect 132770 158624 132776 158636
rect 34572 158596 132776 158624
rect 34572 158584 34578 158596
rect 132770 158584 132776 158596
rect 132828 158584 132834 158636
rect 133874 158584 133880 158636
rect 133932 158624 133938 158636
rect 229094 158624 229100 158636
rect 133932 158596 229100 158624
rect 133932 158584 133938 158596
rect 229094 158584 229100 158596
rect 229152 158584 229158 158636
rect 230014 158584 230020 158636
rect 230072 158624 230078 158636
rect 300394 158624 300400 158636
rect 230072 158596 300400 158624
rect 230072 158584 230078 158596
rect 300394 158584 300400 158596
rect 300452 158584 300458 158636
rect 305454 158584 305460 158636
rect 305512 158624 305518 158636
rect 356238 158624 356244 158636
rect 305512 158596 356244 158624
rect 305512 158584 305518 158596
rect 356238 158584 356244 158596
rect 356296 158584 356302 158636
rect 364426 158584 364432 158636
rect 364484 158624 364490 158636
rect 399938 158624 399944 158636
rect 364484 158596 399944 158624
rect 364484 158584 364490 158596
rect 399938 158584 399944 158596
rect 399996 158584 400002 158636
rect 119982 158516 119988 158568
rect 120040 158556 120046 158568
rect 218882 158556 218888 158568
rect 120040 158528 218888 158556
rect 120040 158516 120046 158528
rect 218882 158516 218888 158528
rect 218940 158516 218946 158568
rect 219618 158516 219624 158568
rect 219676 158556 219682 158568
rect 292666 158556 292672 158568
rect 219676 158528 292672 158556
rect 219676 158516 219682 158528
rect 292666 158516 292672 158528
rect 292724 158516 292730 158568
rect 301958 158516 301964 158568
rect 302016 158556 302022 158568
rect 353662 158556 353668 158568
rect 302016 158528 353668 158556
rect 302016 158516 302022 158528
rect 353662 158516 353668 158528
rect 353720 158516 353726 158568
rect 358354 158516 358360 158568
rect 358412 158556 358418 158568
rect 395430 158556 395436 158568
rect 358412 158528 395436 158556
rect 358412 158516 358418 158528
rect 395430 158516 395436 158528
rect 395488 158516 395494 158568
rect 102594 158448 102600 158500
rect 102652 158488 102658 158500
rect 206002 158488 206008 158500
rect 102652 158460 206008 158488
rect 102652 158448 102658 158460
rect 206002 158448 206008 158460
rect 206060 158448 206066 158500
rect 206646 158448 206652 158500
rect 206704 158488 206710 158500
rect 283098 158488 283104 158500
rect 206704 158460 283104 158488
rect 206704 158448 206710 158460
rect 283098 158448 283104 158460
rect 283156 158448 283162 158500
rect 295058 158448 295064 158500
rect 295116 158488 295122 158500
rect 348510 158488 348516 158500
rect 295116 158460 348516 158488
rect 295116 158448 295122 158460
rect 348510 158448 348516 158460
rect 348568 158448 348574 158500
rect 354030 158448 354036 158500
rect 354088 158488 354094 158500
rect 392210 158488 392216 158500
rect 354088 158460 392216 158488
rect 354088 158448 354094 158460
rect 392210 158448 392216 158460
rect 392268 158448 392274 158500
rect 76650 158380 76656 158432
rect 76708 158420 76714 158432
rect 186498 158420 186504 158432
rect 76708 158392 186504 158420
rect 76708 158380 76714 158392
rect 186498 158380 186504 158392
rect 186556 158380 186562 158432
rect 189350 158380 189356 158432
rect 189408 158420 189414 158432
rect 270218 158420 270224 158432
rect 189408 158392 270224 158420
rect 189408 158380 189414 158392
rect 270218 158380 270224 158392
rect 270276 158380 270282 158432
rect 276842 158380 276848 158432
rect 276900 158420 276906 158432
rect 281442 158420 281448 158432
rect 276900 158392 281448 158420
rect 276900 158380 276906 158392
rect 281442 158380 281448 158392
rect 281500 158380 281506 158432
rect 286410 158380 286416 158432
rect 286468 158420 286474 158432
rect 340782 158420 340788 158432
rect 286468 158392 340788 158420
rect 286468 158380 286474 158392
rect 340782 158380 340788 158392
rect 340840 158380 340846 158432
rect 350534 158380 350540 158432
rect 350592 158420 350598 158432
rect 389634 158420 389640 158432
rect 350592 158392 389640 158420
rect 350592 158380 350598 158392
rect 389634 158380 389640 158392
rect 389692 158380 389698 158432
rect 402946 158420 402974 158664
rect 423674 158420 423680 158432
rect 402946 158392 423680 158420
rect 423674 158380 423680 158392
rect 423732 158380 423738 158432
rect 59354 158312 59360 158364
rect 59412 158352 59418 158364
rect 173894 158352 173900 158364
rect 59412 158324 173900 158352
rect 59412 158312 59418 158324
rect 173894 158312 173900 158324
rect 173952 158312 173958 158364
rect 178862 158312 178868 158364
rect 178920 158352 178926 158364
rect 262490 158352 262496 158364
rect 178920 158324 262496 158352
rect 178920 158312 178926 158324
rect 262490 158312 262496 158324
rect 262548 158312 262554 158364
rect 270402 158312 270408 158364
rect 270460 158352 270466 158364
rect 279234 158352 279240 158364
rect 270460 158324 279240 158352
rect 270460 158312 270466 158324
rect 279234 158312 279240 158324
rect 279292 158312 279298 158364
rect 281166 158312 281172 158364
rect 281224 158352 281230 158364
rect 338298 158352 338304 158364
rect 281224 158324 338304 158352
rect 281224 158312 281230 158324
rect 338298 158312 338304 158324
rect 338356 158312 338362 158364
rect 344462 158312 344468 158364
rect 344520 158352 344526 158364
rect 384942 158352 384948 158364
rect 344520 158324 384948 158352
rect 344520 158312 344526 158324
rect 384942 158312 384948 158324
rect 385000 158312 385006 158364
rect 389542 158312 389548 158364
rect 389600 158352 389606 158364
rect 418522 158352 418528 158364
rect 389600 158324 418528 158352
rect 389600 158312 389606 158324
rect 418522 158312 418528 158324
rect 418580 158312 418586 158364
rect 51442 158244 51448 158296
rect 51500 158284 51506 158296
rect 168098 158284 168104 158296
rect 51500 158256 168104 158284
rect 51500 158244 51506 158256
rect 168098 158244 168104 158256
rect 168156 158244 168162 158296
rect 168742 158284 168748 158296
rect 168392 158256 168748 158284
rect 52454 158176 52460 158228
rect 52512 158216 52518 158228
rect 168392 158216 168420 158256
rect 168742 158244 168748 158256
rect 168800 158244 168806 158296
rect 175458 158244 175464 158296
rect 175516 158284 175522 158296
rect 259914 158284 259920 158296
rect 175516 158256 259920 158284
rect 175516 158244 175522 158256
rect 259914 158244 259920 158256
rect 259972 158244 259978 158296
rect 268194 158244 268200 158296
rect 268252 158284 268258 158296
rect 328638 158284 328644 158296
rect 268252 158256 328644 158284
rect 268252 158244 268258 158256
rect 328638 158244 328644 158256
rect 328696 158244 328702 158296
rect 334066 158244 334072 158296
rect 334124 158284 334130 158296
rect 377398 158284 377404 158296
rect 334124 158256 377404 158284
rect 334124 158244 334130 158256
rect 377398 158244 377404 158256
rect 377456 158244 377462 158296
rect 378318 158244 378324 158296
rect 378376 158284 378382 158296
rect 410150 158284 410156 158296
rect 378376 158256 410156 158284
rect 378376 158244 378382 158256
rect 410150 158244 410156 158256
rect 410208 158244 410214 158296
rect 52512 158188 168420 158216
rect 52512 158176 52518 158188
rect 168466 158176 168472 158228
rect 168524 158216 168530 158228
rect 254026 158216 254032 158228
rect 168524 158188 254032 158216
rect 168524 158176 168530 158188
rect 254026 158176 254032 158188
rect 254084 158176 254090 158228
rect 254302 158176 254308 158228
rect 254360 158216 254366 158228
rect 318334 158216 318340 158228
rect 254360 158188 318340 158216
rect 254360 158176 254366 158188
rect 318334 158176 318340 158188
rect 318392 158176 318398 158228
rect 322842 158176 322848 158228
rect 322900 158216 322906 158228
rect 369118 158216 369124 158228
rect 322900 158188 369124 158216
rect 322900 158176 322906 158188
rect 369118 158176 369124 158188
rect 369176 158176 369182 158228
rect 375650 158176 375656 158228
rect 375708 158216 375714 158228
rect 408218 158216 408224 158228
rect 375708 158188 408224 158216
rect 375708 158176 375714 158188
rect 408218 158176 408224 158188
rect 408276 158176 408282 158228
rect 15102 158108 15108 158160
rect 15160 158148 15166 158160
rect 141142 158148 141148 158160
rect 15160 158120 141148 158148
rect 15160 158108 15166 158120
rect 141142 158108 141148 158120
rect 141200 158108 141206 158160
rect 147674 158108 147680 158160
rect 147732 158148 147738 158160
rect 239398 158148 239404 158160
rect 147732 158120 239404 158148
rect 147732 158108 147738 158120
rect 239398 158108 239404 158120
rect 239456 158108 239462 158160
rect 250898 158108 250904 158160
rect 250956 158148 250962 158160
rect 315758 158148 315764 158160
rect 250956 158120 315764 158148
rect 250956 158108 250962 158120
rect 315758 158108 315764 158120
rect 315816 158108 315822 158160
rect 320174 158108 320180 158160
rect 320232 158148 320238 158160
rect 367186 158148 367192 158160
rect 320232 158120 367192 158148
rect 320232 158108 320238 158120
rect 367186 158108 367192 158120
rect 367244 158108 367250 158160
rect 368750 158108 368756 158160
rect 368808 158148 368814 158160
rect 403158 158148 403164 158160
rect 368808 158120 403164 158148
rect 368808 158108 368814 158120
rect 403158 158108 403164 158120
rect 403216 158108 403222 158160
rect 406010 158108 406016 158160
rect 406068 158148 406074 158160
rect 430758 158148 430764 158160
rect 406068 158120 430764 158148
rect 406068 158108 406074 158120
rect 430758 158108 430764 158120
rect 430816 158108 430822 158160
rect 10778 158040 10784 158092
rect 10836 158080 10842 158092
rect 137922 158080 137928 158092
rect 10836 158052 137928 158080
rect 10836 158040 10842 158052
rect 137922 158040 137928 158052
rect 137980 158040 137986 158092
rect 144270 158040 144276 158092
rect 144328 158080 144334 158092
rect 236822 158080 236828 158092
rect 144328 158052 236828 158080
rect 144328 158040 144334 158052
rect 236822 158040 236828 158052
rect 236880 158040 236886 158092
rect 240042 158040 240048 158092
rect 240100 158080 240106 158092
rect 306190 158080 306196 158092
rect 240100 158052 306196 158080
rect 240100 158040 240106 158052
rect 306190 158040 306196 158052
rect 306248 158040 306254 158092
rect 308950 158040 308956 158092
rect 309008 158080 309014 158092
rect 358814 158080 358820 158092
rect 309008 158052 358820 158080
rect 309008 158040 309014 158052
rect 358814 158040 358820 158052
rect 358872 158040 358878 158092
rect 359182 158040 359188 158092
rect 359240 158080 359246 158092
rect 394602 158080 394608 158092
rect 359240 158052 394608 158080
rect 359240 158040 359246 158052
rect 394602 158040 394608 158052
rect 394660 158040 394666 158092
rect 395614 158040 395620 158092
rect 395672 158080 395678 158092
rect 423030 158080 423036 158092
rect 395672 158052 423036 158080
rect 395672 158040 395678 158052
rect 423030 158040 423036 158052
rect 423088 158040 423094 158092
rect 423398 158040 423404 158092
rect 423456 158080 423462 158092
rect 443546 158080 443552 158092
rect 423456 158052 443552 158080
rect 423456 158040 423462 158052
rect 443546 158040 443552 158052
rect 443604 158040 443610 158092
rect 7282 157972 7288 158024
rect 7340 158012 7346 158024
rect 135346 158012 135352 158024
rect 7340 157984 135352 158012
rect 7340 157972 7346 157984
rect 135346 157972 135352 157984
rect 135404 157972 135410 158024
rect 140774 157972 140780 158024
rect 140832 158012 140838 158024
rect 234246 158012 234252 158024
rect 140832 157984 234252 158012
rect 140832 157972 140838 157984
rect 234246 157972 234252 157984
rect 234304 157972 234310 158024
rect 243906 157972 243912 158024
rect 243964 158012 243970 158024
rect 310698 158012 310704 158024
rect 243964 157984 310704 158012
rect 243964 157972 243970 157984
rect 310698 157972 310704 157984
rect 310756 157972 310762 158024
rect 315850 157972 315856 158024
rect 315908 158012 315914 158024
rect 363966 158012 363972 158024
rect 315908 157984 363972 158012
rect 315908 157972 315914 157984
rect 363966 157972 363972 157984
rect 364024 157972 364030 158024
rect 365254 157972 365260 158024
rect 365312 158012 365318 158024
rect 365312 157984 393314 158012
rect 365312 157972 365318 157984
rect 39942 157904 39948 157956
rect 40000 157944 40006 157956
rect 130286 157944 130292 157956
rect 40000 157916 130292 157944
rect 40000 157904 40006 157916
rect 130286 157904 130292 157916
rect 130344 157904 130350 157956
rect 130378 157904 130384 157956
rect 130436 157944 130442 157956
rect 226518 157944 226524 157956
rect 130436 157916 226524 157944
rect 130436 157904 130442 157916
rect 226518 157904 226524 157916
rect 226576 157904 226582 157956
rect 257798 157904 257804 157956
rect 257856 157944 257862 157956
rect 320910 157944 320916 157956
rect 257856 157916 320916 157944
rect 257856 157904 257862 157916
rect 320910 157904 320916 157916
rect 320968 157904 320974 157956
rect 347958 157904 347964 157956
rect 348016 157944 348022 157956
rect 387702 157944 387708 157956
rect 348016 157916 387708 157944
rect 348016 157904 348022 157916
rect 387702 157904 387708 157916
rect 387760 157904 387766 157956
rect 393286 157944 393314 157984
rect 400214 157972 400220 158024
rect 400272 158012 400278 158024
rect 426250 158012 426256 158024
rect 400272 157984 426256 158012
rect 400272 157972 400278 157984
rect 426250 157972 426256 157984
rect 426308 157972 426314 158024
rect 443270 157972 443276 158024
rect 443328 158012 443334 158024
rect 458358 158012 458364 158024
rect 443328 157984 458364 158012
rect 443328 157972 443334 157984
rect 458358 157972 458364 157984
rect 458416 157972 458422 158024
rect 400582 157944 400588 157956
rect 393286 157916 400588 157944
rect 400582 157904 400588 157916
rect 400640 157904 400646 157956
rect 80054 157836 80060 157888
rect 80112 157876 80118 157888
rect 155954 157876 155960 157888
rect 80112 157848 155960 157876
rect 80112 157836 80118 157848
rect 155954 157836 155960 157848
rect 156012 157836 156018 157888
rect 158070 157836 158076 157888
rect 158128 157876 158134 157888
rect 247126 157876 247132 157888
rect 158128 157848 247132 157876
rect 158128 157836 158134 157848
rect 247126 157836 247132 157848
rect 247184 157836 247190 157888
rect 260558 157836 260564 157888
rect 260616 157876 260622 157888
rect 275370 157876 275376 157888
rect 260616 157848 275376 157876
rect 260616 157836 260622 157848
rect 275370 157836 275376 157848
rect 275428 157836 275434 157888
rect 291562 157836 291568 157888
rect 291620 157876 291626 157888
rect 345934 157876 345940 157888
rect 291620 157848 345940 157876
rect 291620 157836 291626 157848
rect 345934 157836 345940 157848
rect 345992 157836 345998 157888
rect 356606 157836 356612 157888
rect 356664 157876 356670 157888
rect 357618 157876 357624 157888
rect 356664 157848 357624 157876
rect 356664 157836 356670 157848
rect 357618 157836 357624 157848
rect 357676 157836 357682 157888
rect 224954 157768 224960 157820
rect 225012 157808 225018 157820
rect 288158 157808 288164 157820
rect 225012 157780 288164 157808
rect 225012 157768 225018 157780
rect 288158 157768 288164 157780
rect 288216 157768 288222 157820
rect 318702 157768 318708 157820
rect 318760 157808 318766 157820
rect 362586 157808 362592 157820
rect 318760 157780 362592 157808
rect 318760 157768 318766 157780
rect 362586 157768 362592 157780
rect 362644 157768 362650 157820
rect 283834 157700 283840 157752
rect 283892 157740 283898 157752
rect 285674 157740 285680 157752
rect 283892 157712 285680 157740
rect 283892 157700 283898 157712
rect 285674 157700 285680 157712
rect 285732 157700 285738 157752
rect 339402 157700 339408 157752
rect 339460 157740 339466 157752
rect 354950 157740 354956 157752
rect 339460 157712 354956 157740
rect 339460 157700 339466 157712
rect 354950 157700 354956 157712
rect 355008 157700 355014 157752
rect 341886 157632 341892 157684
rect 341944 157672 341950 157684
rect 343542 157672 343548 157684
rect 341944 157644 343548 157672
rect 341944 157632 341950 157644
rect 343542 157632 343548 157644
rect 343600 157632 343606 157684
rect 254026 157360 254032 157412
rect 254084 157400 254090 157412
rect 254762 157400 254768 157412
rect 254084 157372 254768 157400
rect 254084 157360 254090 157372
rect 254762 157360 254768 157372
rect 254820 157360 254826 157412
rect 531958 157360 531964 157412
rect 532016 157400 532022 157412
rect 535454 157400 535460 157412
rect 532016 157372 535460 157400
rect 532016 157360 532022 157372
rect 535454 157360 535460 157372
rect 535512 157360 535518 157412
rect 108666 157292 108672 157344
rect 108724 157332 108730 157344
rect 210510 157332 210516 157344
rect 108724 157304 210516 157332
rect 108724 157292 108730 157304
rect 210510 157292 210516 157304
rect 210568 157292 210574 157344
rect 217042 157292 217048 157344
rect 217100 157332 217106 157344
rect 290734 157332 290740 157344
rect 217100 157304 290740 157332
rect 217100 157292 217106 157304
rect 290734 157292 290740 157304
rect 290792 157292 290798 157344
rect 327166 157292 327172 157344
rect 327224 157332 327230 157344
rect 372338 157332 372344 157344
rect 327224 157304 372344 157332
rect 327224 157292 327230 157304
rect 372338 157292 372344 157304
rect 372396 157292 372402 157344
rect 379146 157292 379152 157344
rect 379204 157332 379210 157344
rect 408494 157332 408500 157344
rect 379204 157304 408500 157332
rect 379204 157292 379210 157304
rect 408494 157292 408500 157304
rect 408552 157292 408558 157344
rect 103514 157224 103520 157276
rect 103572 157264 103578 157276
rect 103572 157236 205680 157264
rect 103572 157224 103578 157236
rect 106090 157156 106096 157208
rect 106148 157196 106154 157208
rect 205545 157199 205603 157205
rect 205545 157196 205557 157199
rect 106148 157168 205557 157196
rect 106148 157156 106154 157168
rect 205545 157165 205557 157168
rect 205591 157165 205603 157199
rect 205652 157196 205680 157236
rect 205818 157224 205824 157276
rect 205876 157264 205882 157276
rect 282454 157264 282460 157276
rect 205876 157236 282460 157264
rect 205876 157224 205882 157236
rect 282454 157224 282460 157236
rect 282512 157224 282518 157276
rect 283006 157224 283012 157276
rect 283064 157264 283070 157276
rect 331858 157264 331864 157276
rect 283064 157236 331864 157264
rect 283064 157224 283070 157236
rect 331858 157224 331864 157236
rect 331916 157224 331922 157276
rect 335814 157224 335820 157276
rect 335872 157264 335878 157276
rect 337194 157264 337200 157276
rect 335872 157236 337200 157264
rect 335872 157224 335878 157236
rect 337194 157224 337200 157236
rect 337252 157224 337258 157276
rect 348786 157224 348792 157276
rect 348844 157264 348850 157276
rect 388346 157264 388352 157276
rect 348844 157236 388352 157264
rect 348844 157224 348850 157236
rect 388346 157224 388352 157236
rect 388404 157224 388410 157276
rect 388438 157224 388444 157276
rect 388496 157264 388502 157276
rect 406378 157264 406384 157276
rect 388496 157236 406384 157264
rect 388496 157224 388502 157236
rect 406378 157224 406384 157236
rect 406436 157224 406442 157276
rect 206646 157196 206652 157208
rect 205652 157168 206652 157196
rect 205545 157159 205603 157165
rect 206646 157156 206652 157168
rect 206704 157156 206710 157208
rect 209222 157156 209228 157208
rect 209280 157196 209286 157208
rect 284938 157196 284944 157208
rect 209280 157168 284944 157196
rect 209280 157156 209286 157168
rect 284938 157156 284944 157168
rect 284996 157156 285002 157208
rect 316770 157156 316776 157208
rect 316828 157196 316834 157208
rect 364610 157196 364616 157208
rect 316828 157168 364616 157196
rect 316828 157156 316834 157168
rect 364610 157156 364616 157168
rect 364668 157156 364674 157208
rect 367830 157156 367836 157208
rect 367888 157196 367894 157208
rect 402422 157196 402428 157208
rect 367888 157168 402428 157196
rect 367888 157156 367894 157168
rect 402422 157156 402428 157168
rect 402480 157156 402486 157208
rect 28902 157088 28908 157140
rect 28960 157128 28966 157140
rect 134058 157128 134064 157140
rect 28960 157100 134064 157128
rect 28960 157088 28966 157100
rect 134058 157088 134064 157100
rect 134116 157088 134122 157140
rect 137278 157088 137284 157140
rect 137336 157128 137342 157140
rect 231670 157128 231676 157140
rect 137336 157100 231676 157128
rect 137336 157088 137342 157100
rect 231670 157088 231676 157100
rect 231728 157088 231734 157140
rect 231762 157088 231768 157140
rect 231820 157128 231826 157140
rect 295794 157128 295800 157140
rect 231820 157100 295800 157128
rect 231820 157088 231826 157100
rect 295794 157088 295800 157100
rect 295852 157088 295858 157140
rect 306374 157088 306380 157140
rect 306432 157128 306438 157140
rect 356882 157128 356888 157140
rect 306432 157100 356888 157128
rect 306432 157088 306438 157100
rect 356882 157088 356888 157100
rect 356940 157088 356946 157140
rect 360930 157088 360936 157140
rect 360988 157128 360994 157140
rect 397362 157128 397368 157140
rect 360988 157100 397368 157128
rect 360988 157088 360994 157100
rect 397362 157088 397368 157100
rect 397420 157088 397426 157140
rect 81802 157020 81808 157072
rect 81860 157060 81866 157072
rect 190638 157060 190644 157072
rect 81860 157032 190644 157060
rect 81860 157020 81866 157032
rect 190638 157020 190644 157032
rect 190696 157020 190702 157072
rect 202322 157020 202328 157072
rect 202380 157060 202386 157072
rect 279878 157060 279884 157072
rect 202380 157032 279884 157060
rect 202380 157020 202386 157032
rect 279878 157020 279884 157032
rect 279936 157020 279942 157072
rect 299382 157020 299388 157072
rect 299440 157060 299446 157072
rect 351730 157060 351736 157072
rect 299440 157032 351736 157060
rect 299440 157020 299446 157032
rect 351730 157020 351736 157032
rect 351788 157020 351794 157072
rect 357434 157020 357440 157072
rect 357492 157060 357498 157072
rect 394786 157060 394792 157072
rect 357492 157032 394792 157060
rect 357492 157020 357498 157032
rect 394786 157020 394792 157032
rect 394844 157020 394850 157072
rect 74902 156952 74908 157004
rect 74960 156992 74966 157004
rect 185486 156992 185492 157004
rect 74960 156964 185492 156992
rect 74960 156952 74966 156964
rect 185486 156952 185492 156964
rect 185544 156952 185550 157004
rect 192754 156952 192760 157004
rect 192812 156992 192818 157004
rect 272794 156992 272800 157004
rect 192812 156964 272800 156992
rect 192812 156952 192818 156964
rect 272794 156952 272800 156964
rect 272852 156952 272858 157004
rect 295886 156952 295892 157004
rect 295944 156992 295950 157004
rect 349154 156992 349160 157004
rect 295944 156964 349160 156992
rect 295944 156952 295950 156964
rect 349154 156952 349160 156964
rect 349212 156952 349218 157004
rect 355778 156952 355784 157004
rect 355836 156992 355842 157004
rect 393498 156992 393504 157004
rect 355836 156964 393504 156992
rect 355836 156952 355842 156964
rect 393498 156952 393504 156964
rect 393556 156952 393562 157004
rect 410334 156952 410340 157004
rect 410392 156992 410398 157004
rect 429194 156992 429200 157004
rect 410392 156964 429200 156992
rect 410392 156952 410398 156964
rect 429194 156952 429200 156964
rect 429252 156952 429258 157004
rect 78306 156884 78312 156936
rect 78364 156924 78370 156936
rect 188062 156924 188068 156936
rect 78364 156896 188068 156924
rect 78364 156884 78370 156896
rect 188062 156884 188068 156896
rect 188120 156884 188126 156936
rect 191926 156884 191932 156936
rect 191984 156924 191990 156936
rect 272150 156924 272156 156936
rect 191984 156896 272156 156924
rect 191984 156884 191990 156896
rect 272150 156884 272156 156896
rect 272208 156884 272214 156936
rect 285582 156924 285588 156936
rect 277366 156896 285588 156924
rect 61010 156816 61016 156868
rect 61068 156856 61074 156868
rect 175182 156856 175188 156868
rect 61068 156828 175188 156856
rect 61068 156816 61074 156828
rect 175182 156816 175188 156828
rect 175240 156816 175246 156868
rect 183554 156816 183560 156868
rect 183612 156856 183618 156868
rect 184842 156856 184848 156868
rect 183612 156828 184848 156856
rect 183612 156816 183618 156828
rect 184842 156816 184848 156828
rect 184900 156816 184906 156868
rect 188430 156816 188436 156868
rect 188488 156856 188494 156868
rect 269574 156856 269580 156868
rect 188488 156828 269580 156856
rect 188488 156816 188494 156828
rect 269574 156816 269580 156828
rect 269632 156816 269638 156868
rect 276106 156816 276112 156868
rect 276164 156856 276170 156868
rect 277366 156856 277394 156896
rect 285582 156884 285588 156896
rect 285640 156884 285646 156936
rect 288986 156884 288992 156936
rect 289044 156924 289050 156936
rect 340785 156927 340843 156933
rect 340785 156924 340797 156927
rect 289044 156896 340797 156924
rect 289044 156884 289050 156896
rect 340785 156893 340797 156896
rect 340831 156893 340843 156927
rect 341518 156924 341524 156936
rect 340785 156887 340843 156893
rect 340892 156896 341524 156924
rect 276164 156828 277394 156856
rect 276164 156816 276170 156828
rect 285490 156816 285496 156868
rect 285548 156856 285554 156868
rect 340892 156856 340920 156896
rect 341518 156884 341524 156896
rect 341576 156884 341582 156936
rect 347038 156884 347044 156936
rect 347096 156924 347102 156936
rect 387058 156924 387064 156936
rect 347096 156896 387064 156924
rect 347096 156884 347102 156896
rect 387058 156884 387064 156896
rect 387116 156884 387122 156936
rect 402514 156884 402520 156936
rect 402572 156924 402578 156936
rect 428182 156924 428188 156936
rect 402572 156896 428188 156924
rect 402572 156884 402578 156896
rect 428182 156884 428188 156896
rect 428240 156884 428246 156936
rect 285548 156828 340920 156856
rect 285548 156816 285554 156828
rect 340966 156816 340972 156868
rect 341024 156856 341030 156868
rect 382550 156856 382556 156868
rect 341024 156828 382556 156856
rect 341024 156816 341030 156828
rect 382550 156816 382556 156828
rect 382608 156816 382614 156868
rect 392118 156816 392124 156868
rect 392176 156856 392182 156868
rect 420454 156856 420460 156868
rect 392176 156828 420460 156856
rect 392176 156816 392182 156828
rect 420454 156816 420460 156828
rect 420512 156816 420518 156868
rect 438946 156816 438952 156868
rect 439004 156856 439010 156868
rect 455138 156856 455144 156868
rect 439004 156828 455144 156856
rect 439004 156816 439010 156828
rect 455138 156816 455144 156828
rect 455196 156816 455202 156868
rect 22830 156748 22836 156800
rect 22888 156788 22894 156800
rect 146938 156788 146944 156800
rect 22888 156760 146944 156788
rect 22888 156748 22894 156760
rect 146938 156748 146944 156760
rect 146996 156748 147002 156800
rect 154666 156748 154672 156800
rect 154724 156788 154730 156800
rect 244550 156788 244556 156800
rect 154724 156760 244556 156788
rect 154724 156748 154730 156760
rect 244550 156748 244556 156760
rect 244608 156748 244614 156800
rect 248506 156748 248512 156800
rect 248564 156788 248570 156800
rect 249702 156788 249708 156800
rect 248564 156760 249708 156788
rect 248564 156748 248570 156760
rect 249702 156748 249708 156760
rect 249760 156748 249766 156800
rect 258074 156748 258080 156800
rect 258132 156788 258138 156800
rect 259270 156788 259276 156800
rect 258132 156760 259276 156788
rect 258132 156748 258138 156760
rect 259270 156748 259276 156760
rect 259328 156748 259334 156800
rect 278590 156748 278596 156800
rect 278648 156788 278654 156800
rect 336366 156788 336372 156800
rect 278648 156760 336372 156788
rect 278648 156748 278654 156760
rect 336366 156748 336372 156760
rect 336424 156748 336430 156800
rect 337562 156748 337568 156800
rect 337620 156788 337626 156800
rect 379974 156788 379980 156800
rect 337620 156760 379980 156788
rect 337620 156748 337626 156760
rect 379974 156748 379980 156760
rect 380032 156748 380038 156800
rect 386414 156748 386420 156800
rect 386472 156788 386478 156800
rect 415946 156788 415952 156800
rect 386472 156760 415952 156788
rect 386472 156748 386478 156760
rect 415946 156748 415952 156760
rect 416004 156748 416010 156800
rect 420730 156748 420736 156800
rect 420788 156788 420794 156800
rect 440234 156788 440240 156800
rect 420788 156760 440240 156788
rect 420788 156748 420794 156760
rect 440234 156748 440240 156760
rect 440292 156748 440298 156800
rect 6362 156680 6368 156732
rect 6420 156720 6426 156732
rect 134702 156720 134708 156732
rect 6420 156692 134708 156720
rect 6420 156680 6426 156692
rect 134702 156680 134708 156692
rect 134760 156680 134766 156732
rect 143350 156680 143356 156732
rect 143408 156720 143414 156732
rect 233421 156723 233479 156729
rect 233421 156720 233433 156723
rect 143408 156692 233433 156720
rect 143408 156680 143414 156692
rect 233421 156689 233433 156692
rect 233467 156689 233479 156723
rect 233421 156683 233479 156689
rect 233510 156680 233516 156732
rect 233568 156680 233574 156732
rect 240410 156680 240416 156732
rect 240468 156720 240474 156732
rect 308122 156720 308128 156732
rect 240468 156692 308128 156720
rect 240468 156680 240474 156692
rect 308122 156680 308128 156692
rect 308180 156680 308186 156732
rect 309778 156680 309784 156732
rect 309836 156680 309842 156732
rect 313274 156680 313280 156732
rect 313332 156720 313338 156732
rect 362034 156720 362040 156732
rect 313332 156692 362040 156720
rect 313332 156680 313338 156692
rect 362034 156680 362040 156692
rect 362092 156680 362098 156732
rect 372246 156680 372252 156732
rect 372304 156720 372310 156732
rect 405734 156720 405740 156732
rect 372304 156692 405740 156720
rect 372304 156680 372310 156692
rect 405734 156680 405740 156692
rect 405792 156680 405798 156732
rect 417326 156680 417332 156732
rect 417384 156720 417390 156732
rect 439038 156720 439044 156732
rect 417384 156692 439044 156720
rect 417384 156680 417390 156692
rect 439038 156680 439044 156692
rect 439096 156680 439102 156732
rect 441522 156680 441528 156732
rect 441580 156720 441586 156732
rect 457070 156720 457076 156732
rect 441580 156692 457076 156720
rect 441580 156680 441586 156692
rect 457070 156680 457076 156692
rect 457128 156680 457134 156732
rect 2038 156612 2044 156664
rect 2096 156652 2102 156664
rect 131482 156652 131488 156664
rect 2096 156624 131488 156652
rect 2096 156612 2102 156624
rect 131482 156612 131488 156624
rect 131540 156612 131546 156664
rect 136450 156612 136456 156664
rect 136508 156652 136514 156664
rect 231026 156652 231032 156664
rect 136508 156624 231032 156652
rect 136508 156612 136514 156624
rect 231026 156612 231032 156624
rect 231084 156612 231090 156664
rect 233528 156652 233556 156680
rect 302970 156652 302976 156664
rect 233528 156624 302976 156652
rect 302970 156612 302976 156624
rect 303028 156612 303034 156664
rect 309796 156652 309824 156680
rect 359458 156652 359464 156664
rect 309796 156624 359464 156652
rect 359458 156612 359464 156624
rect 359516 156612 359522 156664
rect 361850 156612 361856 156664
rect 361908 156652 361914 156664
rect 398006 156652 398012 156664
rect 361908 156624 398012 156652
rect 361908 156612 361914 156624
rect 398006 156612 398012 156624
rect 398064 156612 398070 156664
rect 399110 156612 399116 156664
rect 399168 156652 399174 156664
rect 425606 156652 425612 156664
rect 399168 156624 425612 156652
rect 399168 156612 399174 156624
rect 425606 156612 425612 156624
rect 425664 156612 425670 156664
rect 434622 156612 434628 156664
rect 434680 156652 434686 156664
rect 449894 156652 449900 156664
rect 434680 156624 449900 156652
rect 434680 156612 434686 156624
rect 449894 156612 449900 156624
rect 449952 156612 449958 156664
rect 99374 156544 99380 156596
rect 99432 156584 99438 156596
rect 194597 156587 194655 156593
rect 194597 156584 194609 156587
rect 99432 156556 194609 156584
rect 99432 156544 99438 156556
rect 194597 156553 194609 156556
rect 194643 156553 194655 156587
rect 194597 156547 194655 156553
rect 194686 156544 194692 156596
rect 194744 156584 194750 156596
rect 195698 156584 195704 156596
rect 194744 156556 195704 156584
rect 194744 156544 194750 156556
rect 195698 156544 195704 156556
rect 195756 156544 195762 156596
rect 198826 156544 198832 156596
rect 198884 156584 198890 156596
rect 277302 156584 277308 156596
rect 198884 156556 277308 156584
rect 198884 156544 198890 156556
rect 277302 156544 277308 156556
rect 277360 156544 277366 156596
rect 282178 156544 282184 156596
rect 282236 156584 282242 156596
rect 321554 156584 321560 156596
rect 282236 156556 321560 156584
rect 282236 156544 282242 156556
rect 321554 156544 321560 156556
rect 321612 156544 321618 156596
rect 330570 156544 330576 156596
rect 330628 156584 330634 156596
rect 374914 156584 374920 156596
rect 330628 156556 374920 156584
rect 330628 156544 330634 156556
rect 374914 156544 374920 156556
rect 374972 156544 374978 156596
rect 123386 156476 123392 156528
rect 123444 156516 123450 156528
rect 221458 156516 221464 156528
rect 123444 156488 221464 156516
rect 123444 156476 123450 156488
rect 221458 156476 221464 156488
rect 221516 156476 221522 156528
rect 223390 156476 223396 156528
rect 223448 156516 223454 156528
rect 295242 156516 295248 156528
rect 223448 156488 295248 156516
rect 223448 156476 223454 156488
rect 295242 156476 295248 156488
rect 295300 156476 295306 156528
rect 308306 156476 308312 156528
rect 308364 156516 308370 156528
rect 344738 156516 344744 156528
rect 308364 156488 344744 156516
rect 308364 156476 308370 156488
rect 344738 156476 344744 156488
rect 344796 156476 344802 156528
rect 165614 156408 165620 156460
rect 165672 156448 165678 156460
rect 166810 156448 166816 156460
rect 165672 156420 166816 156448
rect 165672 156408 165678 156420
rect 166810 156408 166816 156420
rect 166868 156408 166874 156460
rect 183462 156408 183468 156460
rect 183520 156448 183526 156460
rect 191282 156448 191288 156460
rect 183520 156420 191288 156448
rect 183520 156408 183526 156420
rect 191282 156408 191288 156420
rect 191340 156408 191346 156460
rect 194597 156451 194655 156457
rect 194597 156417 194609 156451
rect 194643 156448 194655 156451
rect 197630 156448 197636 156460
rect 194643 156420 197636 156448
rect 194643 156417 194655 156420
rect 194597 156411 194655 156417
rect 197630 156408 197636 156420
rect 197688 156408 197694 156460
rect 205545 156451 205603 156457
rect 205545 156417 205557 156451
rect 205591 156448 205603 156451
rect 208578 156448 208584 156460
rect 205591 156420 208584 156448
rect 205591 156417 205603 156420
rect 205545 156411 205603 156417
rect 208578 156408 208584 156420
rect 208636 156408 208642 156460
rect 233421 156451 233479 156457
rect 233421 156417 233433 156451
rect 233467 156448 233479 156451
rect 236178 156448 236184 156460
rect 233467 156420 236184 156448
rect 233467 156417 233479 156420
rect 233421 156411 233479 156417
rect 236178 156408 236184 156420
rect 236236 156408 236242 156460
rect 253198 156408 253204 156460
rect 253256 156448 253262 156460
rect 303614 156448 303620 156460
rect 253256 156420 303620 156448
rect 253256 156408 253262 156420
rect 303614 156408 303620 156420
rect 303672 156408 303678 156460
rect 340785 156451 340843 156457
rect 340785 156417 340797 156451
rect 340831 156448 340843 156451
rect 344094 156448 344100 156460
rect 340831 156420 344100 156448
rect 340831 156417 340843 156420
rect 340785 156411 340843 156417
rect 344094 156408 344100 156420
rect 344152 156408 344158 156460
rect 365254 156448 365260 156460
rect 344986 156420 365260 156448
rect 272058 156340 272064 156392
rect 272116 156380 272122 156392
rect 316402 156380 316408 156392
rect 272116 156352 316408 156380
rect 272116 156340 272122 156352
rect 316402 156340 316408 156352
rect 316460 156340 316466 156392
rect 342254 156340 342260 156392
rect 342312 156380 342318 156392
rect 344986 156380 345014 156420
rect 365254 156408 365260 156420
rect 365312 156408 365318 156460
rect 342312 156352 345014 156380
rect 342312 156340 342318 156352
rect 272426 156272 272432 156324
rect 272484 156312 272490 156324
rect 311342 156312 311348 156324
rect 272484 156284 311348 156312
rect 272484 156272 272490 156284
rect 311342 156272 311348 156284
rect 311400 156272 311406 156324
rect 174078 155932 174084 155984
rect 174136 155972 174142 155984
rect 176470 155972 176476 155984
rect 174136 155944 176476 155972
rect 174136 155932 174142 155944
rect 176470 155932 176476 155944
rect 176528 155932 176534 155984
rect 356422 155932 356428 155984
rect 356480 155972 356486 155984
rect 358170 155972 358176 155984
rect 356480 155944 358176 155972
rect 356480 155932 356486 155944
rect 358170 155932 358176 155944
rect 358228 155932 358234 155984
rect 397270 155932 397276 155984
rect 397328 155972 397334 155984
rect 401870 155972 401876 155984
rect 397328 155944 401876 155972
rect 397328 155932 397334 155944
rect 401870 155932 401876 155944
rect 401928 155932 401934 155984
rect 120810 155864 120816 155916
rect 120868 155904 120874 155916
rect 219526 155904 219532 155916
rect 120868 155876 219532 155904
rect 120868 155864 120874 155876
rect 219526 155864 219532 155876
rect 219584 155864 219590 155916
rect 226610 155864 226616 155916
rect 226668 155904 226674 155916
rect 297818 155904 297824 155916
rect 226668 155876 297824 155904
rect 226668 155864 226674 155876
rect 297818 155864 297824 155876
rect 297876 155864 297882 155916
rect 326246 155864 326252 155916
rect 326304 155904 326310 155916
rect 371694 155904 371700 155916
rect 326304 155876 371700 155904
rect 326304 155864 326310 155876
rect 371694 155864 371700 155876
rect 371752 155864 371758 155916
rect 378042 155864 378048 155916
rect 378100 155904 378106 155916
rect 401226 155904 401232 155916
rect 378100 155876 401232 155904
rect 378100 155864 378106 155876
rect 401226 155864 401232 155876
rect 401284 155864 401290 155916
rect 430574 155864 430580 155916
rect 430632 155904 430638 155916
rect 446766 155904 446772 155916
rect 430632 155876 446772 155904
rect 430632 155864 430638 155876
rect 446766 155864 446772 155876
rect 446824 155864 446830 155916
rect 446858 155864 446864 155916
rect 446916 155904 446922 155916
rect 448054 155904 448060 155916
rect 446916 155876 448060 155904
rect 446916 155864 446922 155876
rect 448054 155864 448060 155876
rect 448112 155864 448118 155916
rect 122558 155796 122564 155848
rect 122616 155836 122622 155848
rect 220814 155836 220820 155848
rect 122616 155808 220820 155836
rect 122616 155796 122622 155808
rect 220814 155796 220820 155808
rect 220872 155796 220878 155848
rect 220906 155796 220912 155848
rect 220964 155836 220970 155848
rect 293310 155836 293316 155848
rect 220964 155808 293316 155836
rect 220964 155796 220970 155808
rect 293310 155796 293316 155808
rect 293368 155796 293374 155848
rect 297634 155796 297640 155848
rect 297692 155836 297698 155848
rect 298094 155836 298100 155848
rect 297692 155808 298100 155836
rect 297692 155796 297698 155808
rect 298094 155796 298100 155808
rect 298152 155796 298158 155848
rect 302878 155796 302884 155848
rect 302936 155836 302942 155848
rect 354306 155836 354312 155848
rect 302936 155808 354312 155836
rect 302936 155796 302942 155808
rect 354306 155796 354312 155808
rect 354364 155796 354370 155848
rect 362678 155796 362684 155848
rect 362736 155836 362742 155848
rect 398650 155836 398656 155848
rect 362736 155808 398656 155836
rect 362736 155796 362742 155808
rect 398650 155796 398656 155808
rect 398708 155796 398714 155848
rect 437474 155796 437480 155848
rect 437532 155836 437538 155848
rect 449342 155836 449348 155848
rect 437532 155808 449348 155836
rect 437532 155796 437538 155808
rect 449342 155796 449348 155808
rect 449400 155796 449406 155848
rect 41414 155728 41420 155780
rect 41472 155768 41478 155780
rect 144362 155768 144368 155780
rect 41472 155740 144368 155768
rect 41472 155728 41478 155740
rect 144362 155728 144368 155740
rect 144420 155728 144426 155780
rect 150342 155728 150348 155780
rect 150400 155768 150406 155780
rect 241330 155768 241336 155780
rect 150400 155740 241336 155768
rect 150400 155728 150406 155740
rect 241330 155728 241336 155740
rect 241388 155728 241394 155780
rect 245654 155728 245660 155780
rect 245712 155768 245718 155780
rect 250346 155768 250352 155780
rect 245712 155740 250352 155768
rect 245712 155728 245718 155740
rect 250346 155728 250352 155740
rect 250404 155728 250410 155780
rect 275094 155728 275100 155780
rect 275152 155768 275158 155780
rect 333790 155768 333796 155780
rect 275152 155740 333796 155768
rect 275152 155728 275158 155740
rect 333790 155728 333796 155740
rect 333848 155728 333854 155780
rect 334894 155728 334900 155780
rect 334952 155768 334958 155780
rect 351914 155768 351920 155780
rect 334952 155740 351920 155768
rect 334952 155728 334958 155740
rect 351914 155728 351920 155740
rect 351972 155728 351978 155780
rect 354858 155728 354864 155780
rect 354916 155768 354922 155780
rect 392854 155768 392860 155780
rect 354916 155740 392860 155768
rect 354916 155728 354922 155740
rect 392854 155728 392860 155740
rect 392912 155728 392918 155780
rect 413830 155728 413836 155780
rect 413888 155768 413894 155780
rect 415489 155771 415547 155777
rect 415489 155768 415501 155771
rect 413888 155740 415501 155768
rect 413888 155728 413894 155740
rect 415489 155737 415501 155740
rect 415535 155737 415547 155771
rect 415489 155731 415547 155737
rect 429378 155728 429384 155780
rect 429436 155768 429442 155780
rect 446122 155768 446128 155780
rect 429436 155740 446128 155768
rect 429436 155728 429442 155740
rect 446122 155728 446128 155740
rect 446180 155728 446186 155780
rect 446398 155728 446404 155780
rect 446456 155768 446462 155780
rect 455782 155768 455788 155780
rect 446456 155740 455788 155768
rect 446456 155728 446462 155740
rect 455782 155728 455788 155740
rect 455840 155728 455846 155780
rect 92198 155660 92204 155712
rect 92256 155700 92262 155712
rect 198274 155700 198280 155712
rect 92256 155672 198280 155700
rect 92256 155660 92262 155672
rect 198274 155660 198280 155672
rect 198332 155660 198338 155712
rect 198734 155660 198740 155712
rect 198792 155700 198798 155712
rect 209222 155700 209228 155712
rect 198792 155672 209228 155700
rect 198792 155660 198798 155672
rect 209222 155660 209228 155672
rect 209280 155660 209286 155712
rect 216214 155660 216220 155712
rect 216272 155700 216278 155712
rect 290090 155700 290096 155712
rect 216272 155672 290096 155700
rect 216272 155660 216278 155672
rect 290090 155660 290096 155672
rect 290148 155660 290154 155712
rect 298554 155660 298560 155712
rect 298612 155700 298618 155712
rect 351086 155700 351092 155712
rect 298612 155672 351092 155700
rect 298612 155660 298618 155672
rect 351086 155660 351092 155672
rect 351144 155660 351150 155712
rect 351362 155660 351368 155712
rect 351420 155700 351426 155712
rect 390278 155700 390284 155712
rect 351420 155672 390284 155700
rect 351420 155660 351426 155672
rect 390278 155660 390284 155672
rect 390336 155660 390342 155712
rect 405642 155660 405648 155712
rect 405700 155700 405706 155712
rect 428826 155700 428832 155712
rect 405700 155672 428832 155700
rect 405700 155660 405706 155672
rect 428826 155660 428832 155672
rect 428884 155660 428890 155712
rect 430298 155660 430304 155712
rect 430356 155700 430362 155712
rect 448698 155700 448704 155712
rect 430356 155672 448704 155700
rect 430356 155660 430362 155672
rect 448698 155660 448704 155672
rect 448756 155660 448762 155712
rect 85298 155592 85304 155644
rect 85356 155632 85362 155644
rect 193122 155632 193128 155644
rect 85356 155604 193128 155632
rect 85356 155592 85362 155604
rect 193122 155592 193128 155604
rect 193180 155592 193186 155644
rect 197354 155592 197360 155644
rect 197412 155632 197418 155644
rect 204070 155632 204076 155644
rect 197412 155604 204076 155632
rect 197412 155592 197418 155604
rect 204070 155592 204076 155604
rect 204128 155592 204134 155644
rect 204898 155592 204904 155644
rect 204956 155632 204962 155644
rect 281810 155632 281816 155644
rect 204956 155604 281816 155632
rect 204956 155592 204962 155604
rect 281810 155592 281816 155604
rect 281868 155592 281874 155644
rect 282086 155592 282092 155644
rect 282144 155632 282150 155644
rect 338942 155632 338948 155644
rect 282144 155604 338948 155632
rect 282144 155592 282150 155604
rect 338942 155592 338948 155604
rect 339000 155592 339006 155644
rect 343634 155592 343640 155644
rect 343692 155632 343698 155644
rect 384482 155632 384488 155644
rect 343692 155604 384488 155632
rect 343692 155592 343698 155604
rect 384482 155592 384488 155604
rect 384540 155592 384546 155644
rect 393314 155592 393320 155644
rect 393372 155632 393378 155644
rect 421098 155632 421104 155644
rect 393372 155604 421104 155632
rect 393372 155592 393378 155604
rect 421098 155592 421104 155604
rect 421156 155592 421162 155644
rect 424226 155592 424232 155644
rect 424284 155632 424290 155644
rect 444190 155632 444196 155644
rect 424284 155604 444196 155632
rect 424284 155592 424290 155604
rect 444190 155592 444196 155604
rect 444248 155592 444254 155644
rect 447226 155592 447232 155644
rect 447284 155632 447290 155644
rect 459002 155632 459008 155644
rect 447284 155604 459008 155632
rect 447284 155592 447290 155604
rect 459002 155592 459008 155604
rect 459060 155592 459066 155644
rect 67910 155524 67916 155576
rect 67968 155564 67974 155576
rect 180334 155564 180340 155576
rect 67968 155536 180340 155564
rect 67968 155524 67974 155536
rect 180334 155524 180340 155536
rect 180392 155524 180398 155576
rect 195330 155524 195336 155576
rect 195388 155564 195394 155576
rect 274726 155564 274732 155576
rect 195388 155536 274732 155564
rect 195388 155524 195394 155536
rect 274726 155524 274732 155536
rect 274784 155524 274790 155576
rect 277762 155524 277768 155576
rect 277820 155564 277826 155576
rect 335722 155564 335728 155576
rect 277820 155536 335728 155564
rect 277820 155524 277826 155536
rect 335722 155524 335728 155536
rect 335780 155524 335786 155576
rect 340138 155524 340144 155576
rect 340196 155564 340202 155576
rect 381906 155564 381912 155576
rect 340196 155536 381912 155564
rect 340196 155524 340202 155536
rect 381906 155524 381912 155536
rect 381964 155524 381970 155576
rect 388714 155524 388720 155576
rect 388772 155564 388778 155576
rect 417878 155564 417884 155576
rect 388772 155536 417884 155564
rect 388772 155524 388778 155536
rect 417878 155524 417884 155536
rect 417936 155524 417942 155576
rect 419902 155524 419908 155576
rect 419960 155564 419966 155576
rect 440970 155564 440976 155576
rect 419960 155536 440976 155564
rect 419960 155524 419966 155536
rect 440970 155524 440976 155536
rect 441028 155524 441034 155576
rect 447134 155524 447140 155576
rect 447192 155564 447198 155576
rect 459646 155564 459652 155576
rect 447192 155536 459652 155564
rect 447192 155524 447198 155536
rect 459646 155524 459652 155536
rect 459704 155524 459710 155576
rect 57514 155456 57520 155508
rect 57572 155496 57578 155508
rect 172606 155496 172612 155508
rect 57572 155468 172612 155496
rect 57572 155456 57578 155468
rect 172606 155456 172612 155468
rect 172664 155456 172670 155508
rect 181530 155456 181536 155508
rect 181588 155496 181594 155508
rect 264422 155496 264428 155508
rect 181588 155468 264428 155496
rect 181588 155456 181594 155468
rect 264422 155456 264428 155468
rect 264480 155456 264486 155508
rect 270770 155456 270776 155508
rect 270828 155496 270834 155508
rect 330570 155496 330576 155508
rect 270828 155468 330576 155496
rect 270828 155456 270834 155468
rect 330570 155456 330576 155468
rect 330628 155456 330634 155508
rect 336642 155456 336648 155508
rect 336700 155496 336706 155508
rect 379330 155496 379336 155508
rect 336700 155468 379336 155496
rect 336700 155456 336706 155468
rect 379330 155456 379336 155468
rect 379388 155456 379394 155508
rect 384206 155456 384212 155508
rect 384264 155496 384270 155508
rect 413370 155496 413376 155508
rect 384264 155468 413376 155496
rect 384264 155456 384270 155468
rect 413370 155456 413376 155468
rect 413428 155456 413434 155508
rect 435910 155496 435916 155508
rect 415412 155468 435916 155496
rect 44542 155388 44548 155440
rect 44600 155428 44606 155440
rect 162946 155428 162952 155440
rect 44600 155400 162952 155428
rect 44600 155388 44606 155400
rect 162946 155388 162952 155400
rect 163004 155388 163010 155440
rect 171410 155388 171416 155440
rect 171468 155428 171474 155440
rect 256694 155428 256700 155440
rect 171468 155400 256700 155428
rect 171468 155388 171474 155400
rect 256694 155388 256700 155400
rect 256752 155388 256758 155440
rect 267366 155388 267372 155440
rect 267424 155428 267430 155440
rect 327994 155428 328000 155440
rect 267424 155400 328000 155428
rect 267424 155388 267430 155400
rect 327994 155388 328000 155400
rect 328052 155388 328058 155440
rect 333238 155388 333244 155440
rect 333296 155428 333302 155440
rect 376754 155428 376760 155440
rect 333296 155400 376760 155428
rect 333296 155388 333302 155400
rect 376754 155388 376760 155400
rect 376812 155388 376818 155440
rect 385218 155388 385224 155440
rect 385276 155428 385282 155440
rect 415302 155428 415308 155440
rect 385276 155400 415308 155428
rect 385276 155388 385282 155400
rect 415302 155388 415308 155400
rect 415360 155388 415366 155440
rect 29822 155320 29828 155372
rect 29880 155360 29886 155372
rect 152090 155360 152096 155372
rect 29880 155332 152096 155360
rect 29880 155320 29886 155332
rect 152090 155320 152096 155332
rect 152148 155320 152154 155372
rect 165062 155320 165068 155372
rect 165120 155360 165126 155372
rect 252278 155360 252284 155372
rect 165120 155332 252284 155360
rect 165120 155320 165126 155332
rect 252278 155320 252284 155332
rect 252336 155320 252342 155372
rect 260374 155320 260380 155372
rect 260432 155360 260438 155372
rect 322842 155360 322848 155372
rect 260432 155332 322848 155360
rect 260432 155320 260438 155332
rect 322842 155320 322848 155332
rect 322900 155320 322906 155372
rect 329742 155320 329748 155372
rect 329800 155360 329806 155372
rect 374270 155360 374276 155372
rect 329800 155332 374276 155360
rect 329800 155320 329806 155332
rect 374270 155320 374276 155332
rect 374328 155320 374334 155372
rect 381722 155320 381728 155372
rect 381780 155360 381786 155372
rect 412726 155360 412732 155372
rect 381780 155332 412732 155360
rect 381780 155320 381786 155332
rect 412726 155320 412732 155332
rect 412784 155320 412790 155372
rect 412910 155320 412916 155372
rect 412968 155360 412974 155372
rect 415412 155360 415440 155468
rect 435910 155456 435916 155468
rect 435968 155456 435974 155508
rect 445662 155456 445668 155508
rect 445720 155496 445726 155508
rect 457714 155496 457720 155508
rect 445720 155468 457720 155496
rect 445720 155456 445726 155468
rect 457714 155456 457720 155468
rect 457772 155456 457778 155508
rect 416406 155388 416412 155440
rect 416464 155428 416470 155440
rect 438394 155428 438400 155440
rect 416464 155400 438400 155428
rect 416464 155388 416470 155400
rect 438394 155388 438400 155400
rect 438452 155388 438458 155440
rect 440694 155388 440700 155440
rect 440752 155428 440758 155440
rect 456426 155428 456432 155440
rect 440752 155400 456432 155428
rect 440752 155388 440758 155400
rect 456426 155388 456432 155400
rect 456484 155388 456490 155440
rect 412968 155332 415440 155360
rect 415489 155363 415547 155369
rect 412968 155320 412974 155332
rect 415489 155329 415501 155363
rect 415535 155360 415547 155363
rect 436554 155360 436560 155372
rect 415535 155332 436560 155360
rect 415535 155329 415547 155332
rect 415489 155323 415547 155329
rect 436554 155320 436560 155332
rect 436612 155320 436618 155372
rect 438118 155320 438124 155372
rect 438176 155360 438182 155372
rect 454494 155360 454500 155372
rect 438176 155332 454500 155360
rect 438176 155320 438182 155332
rect 454494 155320 454500 155332
rect 454552 155320 454558 155372
rect 25498 155252 25504 155304
rect 25556 155292 25562 155304
rect 148870 155292 148876 155304
rect 25556 155264 148876 155292
rect 25556 155252 25562 155264
rect 148870 155252 148876 155264
rect 148928 155252 148934 155304
rect 151170 155252 151176 155304
rect 151228 155292 151234 155304
rect 241974 155292 241980 155304
rect 151228 155264 241980 155292
rect 151228 155252 151234 155264
rect 241974 155252 241980 155264
rect 242032 155252 242038 155304
rect 261938 155252 261944 155304
rect 261996 155292 262002 155304
rect 323486 155292 323492 155304
rect 261996 155264 323492 155292
rect 261996 155252 262002 155264
rect 323486 155252 323492 155264
rect 323544 155252 323550 155304
rect 323670 155252 323676 155304
rect 323728 155292 323734 155304
rect 369762 155292 369768 155304
rect 323728 155264 369768 155292
rect 323728 155252 323734 155264
rect 369762 155252 369768 155264
rect 369820 155252 369826 155304
rect 371326 155252 371332 155304
rect 371384 155292 371390 155304
rect 405090 155292 405096 155304
rect 371384 155264 405096 155292
rect 371384 155252 371390 155264
rect 405090 155252 405096 155264
rect 405148 155252 405154 155304
rect 407114 155252 407120 155304
rect 407172 155292 407178 155304
rect 431402 155292 431408 155304
rect 407172 155264 431408 155292
rect 407172 155252 407178 155264
rect 431402 155252 431408 155264
rect 431460 155252 431466 155304
rect 437198 155252 437204 155304
rect 437256 155292 437262 155304
rect 453850 155292 453856 155304
rect 437256 155264 453856 155292
rect 437256 155252 437262 155264
rect 453850 155252 453856 155264
rect 453908 155252 453914 155304
rect 13814 155184 13820 155236
rect 13872 155224 13878 155236
rect 139210 155224 139216 155236
rect 13872 155196 139216 155224
rect 13872 155184 13878 155196
rect 139210 155184 139216 155196
rect 139268 155184 139274 155236
rect 145098 155184 145104 155236
rect 145156 155224 145162 155236
rect 237466 155224 237472 155236
rect 145156 155196 237472 155224
rect 145156 155184 145162 155196
rect 237466 155184 237472 155196
rect 237524 155184 237530 155236
rect 247954 155184 247960 155236
rect 248012 155224 248018 155236
rect 313274 155224 313280 155236
rect 248012 155196 313280 155224
rect 248012 155184 248018 155196
rect 313274 155184 313280 155196
rect 313332 155184 313338 155236
rect 319346 155184 319352 155236
rect 319404 155224 319410 155236
rect 366542 155224 366548 155236
rect 319404 155196 366548 155224
rect 319404 155184 319410 155196
rect 366542 155184 366548 155196
rect 366600 155184 366606 155236
rect 369578 155184 369584 155236
rect 369636 155224 369642 155236
rect 372614 155224 372620 155236
rect 369636 155196 372620 155224
rect 369636 155184 369642 155196
rect 372614 155184 372620 155196
rect 372672 155184 372678 155236
rect 374822 155184 374828 155236
rect 374880 155224 374886 155236
rect 407574 155224 407580 155236
rect 374880 155196 407580 155224
rect 374880 155184 374886 155196
rect 407574 155184 407580 155196
rect 407632 155184 407638 155236
rect 409506 155184 409512 155236
rect 409564 155224 409570 155236
rect 433334 155224 433340 155236
rect 409564 155196 433340 155224
rect 409564 155184 409570 155196
rect 433334 155184 433340 155196
rect 433392 155184 433398 155236
rect 433794 155184 433800 155236
rect 433852 155224 433858 155236
rect 451274 155224 451280 155236
rect 433852 155196 451280 155224
rect 433852 155184 433858 155196
rect 451274 155184 451280 155196
rect 451332 155184 451338 155236
rect 129458 155116 129464 155168
rect 129516 155156 129522 155168
rect 225874 155156 225880 155168
rect 129516 155128 225880 155156
rect 129516 155116 129522 155128
rect 225874 155116 225880 155128
rect 225932 155116 225938 155168
rect 237006 155116 237012 155168
rect 237064 155156 237070 155168
rect 305546 155156 305552 155168
rect 237064 155128 305552 155156
rect 237064 155116 237070 155128
rect 305546 155116 305552 155128
rect 305604 155116 305610 155168
rect 311066 155116 311072 155168
rect 311124 155156 311130 155168
rect 339586 155156 339592 155168
rect 311124 155128 339592 155156
rect 311124 155116 311130 155128
rect 339586 155116 339592 155128
rect 339644 155116 339650 155168
rect 352282 155116 352288 155168
rect 352340 155156 352346 155168
rect 387794 155156 387800 155168
rect 352340 155128 387800 155156
rect 352340 155116 352346 155128
rect 387794 155116 387800 155128
rect 387852 155116 387858 155168
rect 175826 155048 175832 155100
rect 175884 155088 175890 155100
rect 186130 155088 186136 155100
rect 175884 155060 186136 155088
rect 175884 155048 175890 155060
rect 186130 155048 186136 155060
rect 186188 155048 186194 155100
rect 186222 155048 186228 155100
rect 186280 155088 186286 155100
rect 196342 155088 196348 155100
rect 186280 155060 196348 155088
rect 186280 155048 186286 155060
rect 196342 155048 196348 155060
rect 196400 155048 196406 155100
rect 213638 155048 213644 155100
rect 213696 155088 213702 155100
rect 287514 155088 287520 155100
rect 213696 155060 287520 155088
rect 213696 155048 213702 155060
rect 287514 155048 287520 155060
rect 287572 155048 287578 155100
rect 288250 155048 288256 155100
rect 288308 155088 288314 155100
rect 343450 155088 343456 155100
rect 288308 155060 343456 155088
rect 288308 155048 288314 155060
rect 343450 155048 343456 155060
rect 343508 155048 343514 155100
rect 346302 155048 346308 155100
rect 346360 155088 346366 155100
rect 360102 155088 360108 155100
rect 346360 155060 360108 155088
rect 346360 155048 346366 155060
rect 360102 155048 360108 155060
rect 360160 155048 360166 155100
rect 372706 155048 372712 155100
rect 372764 155088 372770 155100
rect 375558 155088 375564 155100
rect 372764 155060 375564 155088
rect 372764 155048 372770 155060
rect 375558 155048 375564 155060
rect 375616 155048 375622 155100
rect 116486 154980 116492 155032
rect 116544 155020 116550 155032
rect 216306 155020 216312 155032
rect 116544 154992 216312 155020
rect 116544 154980 116550 154992
rect 216306 154980 216312 154992
rect 216364 154980 216370 155032
rect 293954 154980 293960 155032
rect 294012 155020 294018 155032
rect 334434 155020 334440 155032
rect 294012 154992 334440 155020
rect 294012 154980 294018 154992
rect 334434 154980 334440 154992
rect 334492 154980 334498 155032
rect 332594 154912 332600 154964
rect 332652 154952 332658 154964
rect 349798 154952 349804 154964
rect 332652 154924 349804 154952
rect 332652 154912 332658 154924
rect 349798 154912 349804 154924
rect 349856 154912 349862 154964
rect 225046 154776 225052 154828
rect 225104 154816 225110 154828
rect 227162 154816 227168 154828
rect 225104 154788 227168 154816
rect 225104 154776 225110 154788
rect 227162 154776 227168 154788
rect 227220 154776 227226 154828
rect 264974 154776 264980 154828
rect 265032 154816 265038 154828
rect 267642 154816 267648 154828
rect 265032 154788 267648 154816
rect 265032 154776 265038 154788
rect 267642 154776 267648 154788
rect 267700 154776 267706 154828
rect 238754 154572 238760 154624
rect 238812 154612 238818 154624
rect 240042 154612 240048 154624
rect 238812 154584 240048 154612
rect 238812 154572 238818 154584
rect 240042 154572 240048 154584
rect 240100 154572 240106 154624
rect 231578 154504 231584 154556
rect 231636 154544 231642 154556
rect 301682 154544 301688 154556
rect 231636 154516 301688 154544
rect 231636 154504 231642 154516
rect 301682 154504 301688 154516
rect 301740 154504 301746 154556
rect 301774 154504 301780 154556
rect 301832 154544 301838 154556
rect 311986 154544 311992 154556
rect 301832 154516 311992 154544
rect 301832 154504 301838 154516
rect 311986 154504 311992 154516
rect 312044 154504 312050 154556
rect 313734 154504 313740 154556
rect 313792 154544 313798 154556
rect 360746 154544 360752 154556
rect 313792 154516 360752 154544
rect 313792 154504 313798 154516
rect 360746 154504 360752 154516
rect 360804 154504 360810 154556
rect 376662 154504 376668 154556
rect 376720 154544 376726 154556
rect 380618 154544 380624 154556
rect 376720 154516 380624 154544
rect 376720 154504 376726 154516
rect 380618 154504 380624 154516
rect 380676 154504 380682 154556
rect 385954 154504 385960 154556
rect 386012 154544 386018 154556
rect 391566 154544 391572 154556
rect 386012 154516 391572 154544
rect 386012 154504 386018 154516
rect 391566 154504 391572 154516
rect 391624 154504 391630 154556
rect 391934 154504 391940 154556
rect 391992 154544 391998 154556
rect 408862 154544 408868 154556
rect 391992 154516 408868 154544
rect 391992 154504 391998 154516
rect 408862 154504 408868 154516
rect 408920 154504 408926 154556
rect 456886 154504 456892 154556
rect 456944 154544 456950 154556
rect 460290 154544 460296 154556
rect 456944 154516 460296 154544
rect 456944 154504 456950 154516
rect 460290 154504 460296 154516
rect 460348 154504 460354 154556
rect 462222 154504 462228 154556
rect 462280 154544 462286 154556
rect 463510 154544 463516 154556
rect 462280 154516 463516 154544
rect 462280 154504 462286 154516
rect 463510 154504 463516 154516
rect 463568 154504 463574 154556
rect 473262 154504 473268 154556
rect 473320 154544 473326 154556
rect 475654 154544 475660 154556
rect 473320 154516 475660 154544
rect 473320 154504 473326 154516
rect 475654 154504 475660 154516
rect 475712 154504 475718 154556
rect 475746 154504 475752 154556
rect 475804 154544 475810 154556
rect 478230 154544 478236 154556
rect 475804 154516 478236 154544
rect 475804 154504 475810 154516
rect 478230 154504 478236 154516
rect 478288 154504 478294 154556
rect 487798 154504 487804 154556
rect 487856 154544 487862 154556
rect 489822 154544 489828 154556
rect 487856 154516 489828 154544
rect 487856 154504 487862 154516
rect 489822 154504 489828 154516
rect 489880 154504 489886 154556
rect 491570 154504 491576 154556
rect 491628 154544 491634 154556
rect 493042 154544 493048 154556
rect 491628 154516 493048 154544
rect 491628 154504 491634 154516
rect 493042 154504 493048 154516
rect 493100 154504 493106 154556
rect 495434 154504 495440 154556
rect 495492 154544 495498 154556
rect 496906 154544 496912 154556
rect 495492 154516 496912 154544
rect 495492 154504 495498 154516
rect 496906 154504 496912 154516
rect 496964 154504 496970 154556
rect 498746 154504 498752 154556
rect 498804 154544 498810 154556
rect 499482 154544 499488 154556
rect 498804 154516 499488 154544
rect 498804 154504 498810 154516
rect 499482 154504 499488 154516
rect 499540 154504 499546 154556
rect 512270 154504 512276 154556
rect 512328 154544 512334 154556
rect 516134 154544 516140 154556
rect 512328 154516 516140 154544
rect 512328 154504 512334 154516
rect 516134 154504 516140 154516
rect 516192 154504 516198 154556
rect 519998 154504 520004 154556
rect 520056 154544 520062 154556
rect 525794 154544 525800 154556
rect 520056 154516 525800 154544
rect 520056 154504 520062 154516
rect 525794 154504 525800 154516
rect 525852 154504 525858 154556
rect 527726 154504 527732 154556
rect 527784 154544 527790 154556
rect 532786 154544 532792 154556
rect 527784 154516 532792 154544
rect 527784 154504 527790 154516
rect 532786 154504 532792 154516
rect 532844 154504 532850 154556
rect 224862 154436 224868 154488
rect 224920 154476 224926 154488
rect 296530 154476 296536 154488
rect 224920 154448 296536 154476
rect 224920 154436 224926 154448
rect 296530 154436 296536 154448
rect 296588 154436 296594 154488
rect 296622 154436 296628 154488
rect 296680 154476 296686 154488
rect 301501 154479 301559 154485
rect 301501 154476 301513 154479
rect 296680 154448 301513 154476
rect 296680 154436 296686 154448
rect 301501 154445 301513 154448
rect 301547 154445 301559 154479
rect 301501 154439 301559 154445
rect 308858 154436 308864 154488
rect 308916 154476 308922 154488
rect 357526 154476 357532 154488
rect 308916 154448 357532 154476
rect 308916 154436 308922 154448
rect 357526 154436 357532 154448
rect 357584 154436 357590 154488
rect 360194 154436 360200 154488
rect 360252 154476 360258 154488
rect 388990 154476 388996 154488
rect 360252 154448 388996 154476
rect 360252 154436 360258 154448
rect 388990 154436 388996 154448
rect 389048 154436 389054 154488
rect 390554 154436 390560 154488
rect 390612 154476 390618 154488
rect 414658 154476 414664 154488
rect 390612 154448 414664 154476
rect 390612 154436 390618 154448
rect 414658 154436 414664 154448
rect 414716 154436 414722 154488
rect 486970 154436 486976 154488
rect 487028 154476 487034 154488
rect 489178 154476 489184 154488
rect 487028 154448 489184 154476
rect 487028 154436 487034 154448
rect 489178 154436 489184 154448
rect 489236 154436 489242 154488
rect 510338 154436 510344 154488
rect 510396 154476 510402 154488
rect 513466 154476 513472 154488
rect 510396 154448 513472 154476
rect 510396 154436 510402 154448
rect 513466 154436 513472 154448
rect 513524 154436 513530 154488
rect 513558 154436 513564 154488
rect 513616 154476 513622 154488
rect 517606 154476 517612 154488
rect 513616 154448 517612 154476
rect 513616 154436 513622 154448
rect 517606 154436 517612 154448
rect 517664 154436 517670 154488
rect 521286 154436 521292 154488
rect 521344 154476 521350 154488
rect 528278 154476 528284 154488
rect 521344 154448 528284 154476
rect 521344 154436 521350 154448
rect 528278 154436 528284 154448
rect 528336 154436 528342 154488
rect 528370 154436 528376 154488
rect 528428 154476 528434 154488
rect 533154 154476 533160 154488
rect 528428 154448 533160 154476
rect 528428 154436 528434 154448
rect 533154 154436 533160 154448
rect 533212 154436 533218 154488
rect 217870 154368 217876 154420
rect 217928 154408 217934 154420
rect 291378 154408 291384 154420
rect 217928 154380 291384 154408
rect 217928 154368 217934 154380
rect 291378 154368 291384 154380
rect 291436 154368 291442 154420
rect 291838 154368 291844 154420
rect 291896 154408 291902 154420
rect 304258 154408 304264 154420
rect 291896 154380 304264 154408
rect 291896 154368 291902 154380
rect 304258 154368 304264 154380
rect 304316 154368 304322 154420
rect 304902 154368 304908 154420
rect 304960 154408 304966 154420
rect 355594 154408 355600 154420
rect 304960 154380 355600 154408
rect 304960 154368 304966 154380
rect 355594 154368 355600 154380
rect 355652 154368 355658 154420
rect 366910 154368 366916 154420
rect 366968 154408 366974 154420
rect 368474 154408 368480 154420
rect 366968 154380 368480 154408
rect 366968 154368 366974 154380
rect 368474 154368 368480 154380
rect 368532 154368 368538 154420
rect 372614 154368 372620 154420
rect 372672 154408 372678 154420
rect 403802 154408 403808 154420
rect 372672 154380 403808 154408
rect 372672 154368 372678 154380
rect 403802 154368 403808 154380
rect 403860 154368 403866 154420
rect 415578 154368 415584 154420
rect 415636 154408 415642 154420
rect 437842 154408 437848 154420
rect 415636 154380 437848 154408
rect 415636 154368 415642 154380
rect 437842 154368 437848 154380
rect 437900 154368 437906 154420
rect 471882 154368 471888 154420
rect 471940 154408 471946 154420
rect 475010 154408 475016 154420
rect 471940 154380 475016 154408
rect 471940 154368 471946 154380
rect 475010 154368 475016 154380
rect 475068 154368 475074 154420
rect 476114 154368 476120 154420
rect 476172 154408 476178 154420
rect 479518 154408 479524 154420
rect 476172 154380 479524 154408
rect 476172 154368 476178 154380
rect 479518 154368 479524 154380
rect 479576 154368 479582 154420
rect 512914 154368 512920 154420
rect 512972 154408 512978 154420
rect 516962 154408 516968 154420
rect 512972 154380 516968 154408
rect 512972 154368 512978 154380
rect 516962 154368 516968 154380
rect 517020 154368 517026 154420
rect 518710 154408 518716 154420
rect 517072 154380 518716 154408
rect 34422 154300 34428 154352
rect 34480 154340 34486 154352
rect 155310 154340 155316 154352
rect 34480 154312 155316 154340
rect 34480 154300 34486 154312
rect 155310 154300 155316 154312
rect 155368 154300 155374 154352
rect 215110 154300 215116 154352
rect 215168 154340 215174 154352
rect 288802 154340 288808 154352
rect 215168 154312 288808 154340
rect 215168 154300 215174 154312
rect 288802 154300 288808 154312
rect 288860 154300 288866 154352
rect 298094 154300 298100 154352
rect 298152 154340 298158 154352
rect 350442 154340 350448 154352
rect 298152 154312 350448 154340
rect 298152 154300 298158 154312
rect 350442 154300 350448 154312
rect 350500 154300 350506 154352
rect 366266 154300 366272 154352
rect 366324 154340 366330 154352
rect 399294 154340 399300 154352
rect 366324 154312 399300 154340
rect 366324 154300 366330 154312
rect 399294 154300 399300 154312
rect 399352 154300 399358 154352
rect 399386 154300 399392 154352
rect 399444 154340 399450 154352
rect 424962 154340 424968 154352
rect 399444 154312 424968 154340
rect 399444 154300 399450 154312
rect 424962 154300 424968 154312
rect 425020 154300 425026 154352
rect 428550 154300 428556 154352
rect 428608 154340 428614 154352
rect 447410 154340 447416 154352
rect 428608 154312 447416 154340
rect 428608 154300 428614 154312
rect 447410 154300 447416 154312
rect 447468 154300 447474 154352
rect 514202 154300 514208 154352
rect 514260 154340 514266 154352
rect 517072 154340 517100 154380
rect 518710 154368 518716 154380
rect 518768 154368 518774 154420
rect 519354 154368 519360 154420
rect 519412 154408 519418 154420
rect 523126 154408 523132 154420
rect 519412 154380 523132 154408
rect 519412 154368 519418 154380
rect 523126 154368 523132 154380
rect 523184 154368 523190 154420
rect 524506 154368 524512 154420
rect 524564 154408 524570 154420
rect 531774 154408 531780 154420
rect 524564 154380 531780 154408
rect 524564 154368 524570 154380
rect 531774 154368 531780 154380
rect 531832 154368 531838 154420
rect 514260 154312 517100 154340
rect 514260 154300 514266 154312
rect 518066 154300 518072 154352
rect 518124 154340 518130 154352
rect 521654 154340 521660 154352
rect 518124 154312 521660 154340
rect 518124 154300 518130 154312
rect 521654 154300 521660 154312
rect 521712 154300 521718 154352
rect 525794 154300 525800 154352
rect 525852 154340 525858 154352
rect 533982 154340 533988 154352
rect 525852 154312 533988 154340
rect 525852 154300 525858 154312
rect 533982 154300 533988 154312
rect 534040 154300 534046 154352
rect 30650 154232 30656 154284
rect 30708 154272 30714 154284
rect 152734 154272 152740 154284
rect 30708 154244 152740 154272
rect 30708 154232 30714 154244
rect 152734 154232 152740 154244
rect 152792 154232 152798 154284
rect 210970 154232 210976 154284
rect 211028 154272 211034 154284
rect 286226 154272 286232 154284
rect 211028 154244 286232 154272
rect 211028 154232 211034 154244
rect 286226 154232 286232 154244
rect 286284 154232 286290 154284
rect 289722 154232 289728 154284
rect 289780 154272 289786 154284
rect 299106 154272 299112 154284
rect 289780 154244 299112 154272
rect 289780 154232 289786 154244
rect 299106 154232 299112 154244
rect 299164 154232 299170 154284
rect 300302 154232 300308 154284
rect 300360 154272 300366 154284
rect 352374 154272 352380 154284
rect 300360 154244 352380 154272
rect 300360 154232 300366 154244
rect 352374 154232 352380 154244
rect 352432 154232 352438 154284
rect 352466 154232 352472 154284
rect 352524 154272 352530 154284
rect 386414 154272 386420 154284
rect 352524 154244 386420 154272
rect 352524 154232 352530 154244
rect 386414 154232 386420 154244
rect 386472 154232 386478 154284
rect 394602 154232 394608 154284
rect 394660 154272 394666 154284
rect 396074 154272 396080 154284
rect 394660 154244 396080 154272
rect 394660 154232 394666 154244
rect 396074 154232 396080 154244
rect 396132 154232 396138 154284
rect 404262 154232 404268 154284
rect 404320 154272 404326 154284
rect 429470 154272 429476 154284
rect 404320 154244 429476 154272
rect 404320 154232 404326 154244
rect 429470 154232 429476 154244
rect 429528 154232 429534 154284
rect 436002 154232 436008 154284
rect 436060 154272 436066 154284
rect 437385 154275 437443 154281
rect 437385 154272 437397 154275
rect 436060 154244 437397 154272
rect 436060 154232 436066 154244
rect 437385 154241 437397 154244
rect 437431 154241 437443 154275
rect 437385 154235 437443 154241
rect 465626 154232 465632 154284
rect 465684 154272 465690 154284
rect 470502 154272 470508 154284
rect 465684 154244 470508 154272
rect 465684 154232 465690 154244
rect 470502 154232 470508 154244
rect 470560 154232 470566 154284
rect 473722 154232 473728 154284
rect 473780 154272 473786 154284
rect 476942 154272 476948 154284
rect 473780 154244 476948 154272
rect 473780 154232 473786 154244
rect 476942 154232 476948 154244
rect 477000 154232 477006 154284
rect 477494 154232 477500 154284
rect 477552 154272 477558 154284
rect 480162 154272 480168 154284
rect 477552 154244 480168 154272
rect 477552 154232 477558 154244
rect 480162 154232 480168 154244
rect 480220 154232 480226 154284
rect 491294 154232 491300 154284
rect 491352 154272 491358 154284
rect 493686 154272 493692 154284
rect 491352 154244 493692 154272
rect 491352 154232 491358 154244
rect 493686 154232 493692 154244
rect 493744 154232 493750 154284
rect 511626 154232 511632 154284
rect 511684 154272 511690 154284
rect 514754 154272 514760 154284
rect 511684 154244 514760 154272
rect 511684 154232 511690 154244
rect 514754 154232 514760 154244
rect 514812 154232 514818 154284
rect 525150 154232 525156 154284
rect 525208 154272 525214 154284
rect 531406 154272 531412 154284
rect 525208 154244 531412 154272
rect 525208 154232 525214 154244
rect 531406 154232 531412 154244
rect 531464 154232 531470 154284
rect 27522 154164 27528 154216
rect 27580 154204 27586 154216
rect 150158 154204 150164 154216
rect 27580 154176 150164 154204
rect 27580 154164 27586 154176
rect 150158 154164 150164 154176
rect 150216 154164 150222 154216
rect 207474 154164 207480 154216
rect 207532 154204 207538 154216
rect 283742 154204 283748 154216
rect 207532 154176 283748 154204
rect 207532 154164 207538 154176
rect 283742 154164 283748 154176
rect 283800 154164 283806 154216
rect 292758 154164 292764 154216
rect 292816 154204 292822 154216
rect 345382 154204 345388 154216
rect 292816 154176 345388 154204
rect 292816 154164 292822 154176
rect 345382 154164 345388 154176
rect 345440 154164 345446 154216
rect 350166 154164 350172 154216
rect 350224 154204 350230 154216
rect 353018 154204 353024 154216
rect 350224 154176 353024 154204
rect 350224 154164 350230 154176
rect 353018 154164 353024 154176
rect 353076 154164 353082 154216
rect 357618 154164 357624 154216
rect 357676 154204 357682 154216
rect 394142 154204 394148 154216
rect 357676 154176 394148 154204
rect 357676 154164 357682 154176
rect 394142 154164 394148 154176
rect 394200 154164 394206 154216
rect 397454 154164 397460 154216
rect 397512 154204 397518 154216
rect 424318 154204 424324 154216
rect 397512 154176 424324 154204
rect 397512 154164 397518 154176
rect 424318 154164 424324 154176
rect 424376 154164 424382 154216
rect 425054 154164 425060 154216
rect 425112 154204 425118 154216
rect 444834 154204 444840 154216
rect 425112 154176 444840 154204
rect 425112 154164 425118 154176
rect 444834 154164 444840 154176
rect 444892 154164 444898 154216
rect 518710 154164 518716 154216
rect 518768 154204 518774 154216
rect 524782 154204 524788 154216
rect 518768 154176 524788 154204
rect 518768 154164 518774 154176
rect 524782 154164 524788 154176
rect 524840 154164 524846 154216
rect 526438 154164 526444 154216
rect 526496 154204 526502 154216
rect 532694 154204 532700 154216
rect 526496 154176 532700 154204
rect 526496 154164 526502 154176
rect 532694 154164 532700 154176
rect 532752 154164 532758 154216
rect 23750 154096 23756 154148
rect 23808 154136 23814 154148
rect 147582 154136 147588 154148
rect 23808 154108 147588 154136
rect 23808 154096 23814 154108
rect 147582 154096 147588 154108
rect 147640 154096 147646 154148
rect 154482 154096 154488 154148
rect 154540 154136 154546 154148
rect 158530 154136 158536 154148
rect 154540 154108 158536 154136
rect 154540 154096 154546 154108
rect 158530 154096 158536 154108
rect 158588 154096 158594 154148
rect 204162 154096 204168 154148
rect 204220 154136 204226 154148
rect 281166 154136 281172 154148
rect 204220 154108 281172 154136
rect 204220 154096 204226 154108
rect 281166 154096 281172 154108
rect 281224 154096 281230 154148
rect 281442 154096 281448 154148
rect 281500 154136 281506 154148
rect 335078 154136 335084 154148
rect 281500 154108 335084 154136
rect 281500 154096 281506 154108
rect 335078 154096 335084 154108
rect 335136 154096 335142 154148
rect 337194 154096 337200 154148
rect 337252 154136 337258 154148
rect 337252 154108 340368 154136
rect 337252 154096 337258 154108
rect 20622 154028 20628 154080
rect 20680 154068 20686 154080
rect 145006 154068 145012 154080
rect 20680 154040 145012 154068
rect 20680 154028 20686 154040
rect 145006 154028 145012 154040
rect 145064 154028 145070 154080
rect 200574 154028 200580 154080
rect 200632 154068 200638 154080
rect 278590 154068 278596 154080
rect 200632 154040 278596 154068
rect 200632 154028 200638 154040
rect 278590 154028 278596 154040
rect 278648 154028 278654 154080
rect 285674 154028 285680 154080
rect 285732 154068 285738 154080
rect 340230 154068 340236 154080
rect 285732 154040 340236 154068
rect 285732 154028 285738 154040
rect 340230 154028 340236 154040
rect 340288 154028 340294 154080
rect 340340 154068 340368 154108
rect 340782 154096 340788 154148
rect 340840 154136 340846 154148
rect 342162 154136 342168 154148
rect 340840 154108 342168 154136
rect 340840 154096 340846 154108
rect 342162 154096 342168 154108
rect 342220 154096 342226 154148
rect 378686 154136 378692 154148
rect 342272 154108 378692 154136
rect 342272 154068 342300 154108
rect 378686 154096 378692 154108
rect 378744 154096 378750 154148
rect 391290 154096 391296 154148
rect 391348 154136 391354 154148
rect 419810 154136 419816 154148
rect 391348 154108 419816 154136
rect 391348 154096 391354 154108
rect 419810 154096 419816 154108
rect 419868 154096 419874 154148
rect 422478 154096 422484 154148
rect 422536 154136 422542 154148
rect 442902 154136 442908 154148
rect 422536 154108 442908 154136
rect 422536 154096 422542 154108
rect 442902 154096 442908 154108
rect 442960 154096 442966 154148
rect 462130 154096 462136 154148
rect 462188 154136 462194 154148
rect 464154 154136 464160 154148
rect 462188 154108 464160 154136
rect 462188 154096 462194 154108
rect 464154 154096 464160 154108
rect 464212 154096 464218 154148
rect 473170 154096 473176 154148
rect 473228 154136 473234 154148
rect 476298 154136 476304 154148
rect 473228 154108 476304 154136
rect 473228 154096 473234 154108
rect 476298 154096 476304 154108
rect 476356 154096 476362 154148
rect 485498 154096 485504 154148
rect 485556 154136 485562 154148
rect 487890 154136 487896 154148
rect 485556 154108 487896 154136
rect 485556 154096 485562 154108
rect 487890 154096 487896 154108
rect 487948 154096 487954 154148
rect 491202 154096 491208 154148
rect 491260 154136 491266 154148
rect 492398 154136 492404 154148
rect 491260 154108 492404 154136
rect 491260 154096 491266 154108
rect 492398 154096 492404 154108
rect 492456 154096 492462 154148
rect 517422 154096 517428 154148
rect 517480 154136 517486 154148
rect 523034 154136 523040 154148
rect 517480 154108 523040 154136
rect 517480 154096 517486 154108
rect 523034 154096 523040 154108
rect 523092 154096 523098 154148
rect 523862 154096 523868 154148
rect 523920 154136 523926 154148
rect 531314 154136 531320 154148
rect 523920 154108 531320 154136
rect 523920 154096 523926 154108
rect 531314 154096 531320 154108
rect 531372 154096 531378 154148
rect 340340 154040 342300 154068
rect 343542 154028 343548 154080
rect 343600 154068 343606 154080
rect 383194 154068 383200 154080
rect 343600 154040 383200 154068
rect 343600 154028 343606 154040
rect 383194 154028 383200 154040
rect 383252 154028 383258 154080
rect 390370 154028 390376 154080
rect 390428 154068 390434 154080
rect 419166 154068 419172 154080
rect 390428 154040 419172 154068
rect 390428 154028 390434 154040
rect 419166 154028 419172 154040
rect 419224 154028 419230 154080
rect 419258 154028 419264 154080
rect 419316 154068 419322 154080
rect 440326 154068 440332 154080
rect 419316 154040 440332 154068
rect 419316 154028 419322 154040
rect 440326 154028 440332 154040
rect 440384 154028 440390 154080
rect 442810 154028 442816 154080
rect 442868 154068 442874 154080
rect 452562 154068 452568 154080
rect 442868 154040 452568 154068
rect 442868 154028 442874 154040
rect 452562 154028 452568 154040
rect 452620 154028 452626 154080
rect 469306 154028 469312 154080
rect 469364 154068 469370 154080
rect 473722 154068 473728 154080
rect 469364 154040 473728 154068
rect 469364 154028 469370 154040
rect 473722 154028 473728 154040
rect 473780 154028 473786 154080
rect 523218 154028 523224 154080
rect 523276 154068 523282 154080
rect 527174 154068 527180 154080
rect 523276 154040 527180 154068
rect 523276 154028 523282 154040
rect 527174 154028 527180 154040
rect 527232 154028 527238 154080
rect 16850 153960 16856 154012
rect 16908 154000 16914 154012
rect 142430 154000 142436 154012
rect 16908 153972 142436 154000
rect 16908 153960 16914 153972
rect 142430 153960 142436 153972
rect 142488 153960 142494 154012
rect 187602 153960 187608 154012
rect 187660 154000 187666 154012
rect 268286 154000 268292 154012
rect 187660 153972 268292 154000
rect 187660 153960 187666 153972
rect 268286 153960 268292 153972
rect 268344 153960 268350 154012
rect 269942 153960 269948 154012
rect 270000 154000 270006 154012
rect 329926 154000 329932 154012
rect 270000 153972 329932 154000
rect 270000 153960 270006 153972
rect 329926 153960 329932 153972
rect 329984 153960 329990 154012
rect 332318 153960 332324 154012
rect 332376 154000 332382 154012
rect 376202 154000 376208 154012
rect 332376 153972 376208 154000
rect 332376 153960 332382 153972
rect 376202 153960 376208 153972
rect 376260 153960 376266 154012
rect 379422 153960 379428 154012
rect 379480 154000 379486 154012
rect 409506 154000 409512 154012
rect 379480 153972 409512 154000
rect 379480 153960 379486 153972
rect 409506 153960 409512 153972
rect 409564 153960 409570 154012
rect 411254 153960 411260 154012
rect 411312 154000 411318 154012
rect 434622 154000 434628 154012
rect 411312 153972 434628 154000
rect 411312 153960 411318 153972
rect 434622 153960 434628 153972
rect 434680 153960 434686 154012
rect 436370 153960 436376 154012
rect 436428 154000 436434 154012
rect 437385 154003 437443 154009
rect 436428 153972 437336 154000
rect 436428 153960 436434 153972
rect 13722 153892 13728 153944
rect 13780 153932 13786 153944
rect 139854 153932 139860 153944
rect 13780 153904 139860 153932
rect 13780 153892 13786 153904
rect 139854 153892 139860 153904
rect 139912 153892 139918 153944
rect 179782 153892 179788 153944
rect 179840 153932 179846 153944
rect 263134 153932 263140 153944
rect 179840 153904 263140 153932
rect 179840 153892 179846 153904
rect 263134 153892 263140 153904
rect 263192 153892 263198 153944
rect 263226 153892 263232 153944
rect 263284 153932 263290 153944
rect 324774 153932 324780 153944
rect 263284 153904 324780 153932
rect 263284 153892 263290 153904
rect 324774 153892 324780 153904
rect 324832 153892 324838 153944
rect 325418 153892 325424 153944
rect 325476 153932 325482 153944
rect 371050 153932 371056 153944
rect 325476 153904 371056 153932
rect 325476 153892 325482 153904
rect 371050 153892 371056 153904
rect 371108 153892 371114 153944
rect 383470 153892 383476 153944
rect 383528 153932 383534 153944
rect 414014 153932 414020 153944
rect 383528 153904 414020 153932
rect 383528 153892 383534 153904
rect 414014 153892 414020 153904
rect 414072 153892 414078 153944
rect 414750 153892 414756 153944
rect 414808 153932 414814 153944
rect 437198 153932 437204 153944
rect 414808 153904 437204 153932
rect 414808 153892 414814 153904
rect 437198 153892 437204 153904
rect 437256 153892 437262 153944
rect 437308 153932 437336 153972
rect 437385 153969 437397 154003
rect 437431 154000 437443 154003
rect 449986 154000 449992 154012
rect 437431 153972 449992 154000
rect 437431 153969 437443 153972
rect 437385 153963 437443 153969
rect 449986 153960 449992 153972
rect 450044 153960 450050 154012
rect 474734 153960 474740 154012
rect 474792 154000 474798 154012
rect 477586 154000 477592 154012
rect 474792 153972 477592 154000
rect 474792 153960 474798 153972
rect 477586 153960 477592 153972
rect 477644 153960 477650 154012
rect 482002 153960 482008 154012
rect 482060 154000 482066 154012
rect 483382 154000 483388 154012
rect 482060 153972 483388 154000
rect 482060 153960 482066 153972
rect 483382 153960 483388 153972
rect 483440 153960 483446 154012
rect 529658 153960 529664 154012
rect 529716 154000 529722 154012
rect 539505 154003 539563 154009
rect 539505 154000 539517 154003
rect 529716 153972 539517 154000
rect 529716 153960 529722 153972
rect 539505 153969 539517 153972
rect 539551 153969 539563 154003
rect 539505 153963 539563 153969
rect 453206 153932 453212 153944
rect 437308 153904 453212 153932
rect 453206 153892 453212 153904
rect 453264 153892 453270 153944
rect 529014 153892 529020 153944
rect 529072 153932 529078 153944
rect 538677 153935 538735 153941
rect 538677 153932 538689 153935
rect 529072 153904 538689 153932
rect 529072 153892 529078 153904
rect 538677 153901 538689 153904
rect 538723 153901 538735 153935
rect 538677 153895 538735 153901
rect 9858 153824 9864 153876
rect 9916 153864 9922 153876
rect 137278 153864 137284 153876
rect 9916 153836 137284 153864
rect 9916 153824 9922 153836
rect 137278 153824 137284 153836
rect 137336 153824 137342 153876
rect 154390 153824 154396 153876
rect 154448 153864 154454 153876
rect 163590 153864 163596 153876
rect 154448 153836 163596 153864
rect 154448 153824 154454 153836
rect 163590 153824 163596 153836
rect 163648 153824 163654 153876
rect 169478 153824 169484 153876
rect 169536 153864 169542 153876
rect 255406 153864 255412 153876
rect 169536 153836 255412 153864
rect 169536 153824 169542 153836
rect 255406 153824 255412 153836
rect 255464 153824 255470 153876
rect 256050 153824 256056 153876
rect 256108 153864 256114 153876
rect 319622 153864 319628 153876
rect 256108 153836 319628 153864
rect 256108 153824 256114 153836
rect 319622 153824 319628 153836
rect 319680 153824 319686 153876
rect 321738 153824 321744 153876
rect 321796 153864 321802 153876
rect 367830 153864 367836 153876
rect 321796 153836 367836 153864
rect 321796 153824 321802 153836
rect 367830 153824 367836 153836
rect 367888 153824 367894 153876
rect 370498 153824 370504 153876
rect 370556 153864 370562 153876
rect 404446 153864 404452 153876
rect 370556 153836 404452 153864
rect 370556 153824 370562 153836
rect 404446 153824 404452 153836
rect 404504 153824 404510 153876
rect 408494 153824 408500 153876
rect 408552 153864 408558 153876
rect 410794 153864 410800 153876
rect 408552 153836 410800 153864
rect 408552 153824 408558 153836
rect 410794 153824 410800 153836
rect 410852 153824 410858 153876
rect 430114 153864 430120 153876
rect 412606 153836 430120 153864
rect 242158 153756 242164 153808
rect 242216 153796 242222 153808
rect 309410 153796 309416 153808
rect 242216 153768 309416 153796
rect 242216 153756 242222 153768
rect 309410 153756 309416 153768
rect 309468 153756 309474 153808
rect 316218 153756 316224 153808
rect 316276 153796 316282 153808
rect 327350 153796 327356 153808
rect 316276 153768 327356 153796
rect 316276 153756 316282 153768
rect 327350 153756 327356 153768
rect 327408 153756 327414 153808
rect 330754 153756 330760 153808
rect 330812 153796 330818 153808
rect 372982 153796 372988 153808
rect 330812 153768 372988 153796
rect 330812 153756 330818 153768
rect 372982 153756 372988 153768
rect 373040 153756 373046 153808
rect 405182 153756 405188 153808
rect 405240 153796 405246 153808
rect 412606 153796 412634 153836
rect 430114 153824 430120 153836
rect 430172 153824 430178 153876
rect 433242 153824 433248 153876
rect 433300 153864 433306 153876
rect 450630 153864 450636 153876
rect 433300 153836 450636 153864
rect 433300 153824 433306 153836
rect 450630 153824 450636 153836
rect 450688 153824 450694 153876
rect 451734 153824 451740 153876
rect 451792 153864 451798 153876
rect 460934 153864 460940 153876
rect 451792 153836 460940 153864
rect 451792 153824 451798 153836
rect 460934 153824 460940 153836
rect 460992 153824 460998 153876
rect 463694 153824 463700 153876
rect 463752 153864 463758 153876
rect 466086 153864 466092 153876
rect 463752 153836 466092 153864
rect 463752 153824 463758 153836
rect 466086 153824 466092 153836
rect 466144 153824 466150 153876
rect 469214 153824 469220 153876
rect 469272 153864 469278 153876
rect 474366 153864 474372 153876
rect 469272 153836 474372 153864
rect 469272 153824 469278 153836
rect 474366 153824 474372 153836
rect 474424 153824 474430 153876
rect 527082 153824 527088 153876
rect 527140 153864 527146 153876
rect 535546 153864 535552 153876
rect 527140 153836 535552 153864
rect 527140 153824 527146 153836
rect 535546 153824 535552 153836
rect 535604 153824 535610 153876
rect 405240 153768 412634 153796
rect 405240 153756 405246 153768
rect 249150 153688 249156 153740
rect 249208 153728 249214 153740
rect 314562 153728 314568 153740
rect 249208 153700 314568 153728
rect 249208 153688 249214 153700
rect 314562 153688 314568 153700
rect 314620 153688 314626 153740
rect 324314 153688 324320 153740
rect 324372 153728 324378 153740
rect 365898 153728 365904 153740
rect 324372 153700 365904 153728
rect 324372 153688 324378 153700
rect 365898 153688 365904 153700
rect 365956 153688 365962 153740
rect 415210 153688 415216 153740
rect 415268 153728 415274 153740
rect 416590 153728 416596 153740
rect 415268 153700 416596 153728
rect 415268 153688 415274 153700
rect 416590 153688 416596 153700
rect 416648 153688 416654 153740
rect 280982 153620 280988 153672
rect 281040 153660 281046 153672
rect 293954 153660 293960 153672
rect 281040 153632 293960 153660
rect 281040 153620 281046 153632
rect 293954 153620 293960 153632
rect 294012 153620 294018 153672
rect 301501 153663 301559 153669
rect 301501 153629 301513 153663
rect 301547 153660 301559 153663
rect 306834 153660 306840 153672
rect 301547 153632 306840 153660
rect 301547 153629 301559 153632
rect 301501 153623 301559 153629
rect 306834 153620 306840 153632
rect 306892 153620 306898 153672
rect 311894 153620 311900 153672
rect 311952 153660 311958 153672
rect 322198 153660 322204 153672
rect 311952 153632 322204 153660
rect 311952 153620 311958 153632
rect 322198 153620 322204 153632
rect 322256 153620 322262 153672
rect 328362 153620 328368 153672
rect 328420 153660 328426 153672
rect 332502 153660 332508 153672
rect 328420 153632 332508 153660
rect 328420 153620 328426 153632
rect 332502 153620 332508 153632
rect 332560 153620 332566 153672
rect 351914 153620 351920 153672
rect 351972 153660 351978 153672
rect 378042 153660 378048 153672
rect 351972 153632 378048 153660
rect 351972 153620 351978 153632
rect 378042 153620 378048 153632
rect 378100 153620 378106 153672
rect 462866 153552 462872 153604
rect 462924 153592 462930 153604
rect 464798 153592 464804 153604
rect 462924 153564 464804 153592
rect 462924 153552 462930 153564
rect 464798 153552 464804 153564
rect 464856 153552 464862 153604
rect 481082 153552 481088 153604
rect 481140 153592 481146 153604
rect 482094 153592 482100 153604
rect 481140 153564 482100 153592
rect 481140 153552 481146 153564
rect 482094 153552 482100 153564
rect 482152 153552 482158 153604
rect 515490 153552 515496 153604
rect 515548 153592 515554 153604
rect 520182 153592 520188 153604
rect 515548 153564 520188 153592
rect 515548 153552 515554 153564
rect 520182 153552 520188 153564
rect 520240 153552 520246 153604
rect 520642 153552 520648 153604
rect 520700 153592 520706 153604
rect 527358 153592 527364 153604
rect 520700 153564 527364 153592
rect 520700 153552 520706 153564
rect 527358 153552 527364 153564
rect 527416 153552 527422 153604
rect 43806 153484 43812 153536
rect 43864 153524 43870 153536
rect 118050 153524 118056 153536
rect 43864 153496 118056 153524
rect 43864 153484 43870 153496
rect 118050 153484 118056 153496
rect 118108 153484 118114 153536
rect 387794 153484 387800 153536
rect 387852 153524 387858 153536
rect 390922 153524 390928 153536
rect 387852 153496 390928 153524
rect 387852 153484 387858 153496
rect 390922 153484 390928 153496
rect 390980 153484 390986 153536
rect 95142 153416 95148 153468
rect 95200 153456 95206 153468
rect 126698 153456 126704 153468
rect 95200 153428 126704 153456
rect 95200 153416 95206 153428
rect 126698 153416 126704 153428
rect 126756 153416 126762 153468
rect 463786 153416 463792 153468
rect 463844 153456 463850 153468
rect 465442 153456 465448 153468
rect 463844 153428 465448 153456
rect 463844 153416 463850 153428
rect 465442 153416 465448 153428
rect 465500 153416 465506 153468
rect 466822 153416 466828 153468
rect 466880 153456 466886 153468
rect 471790 153456 471796 153468
rect 466880 153428 471796 153456
rect 466880 153416 466886 153428
rect 471790 153416 471796 153428
rect 471848 153416 471854 153468
rect 488258 153416 488264 153468
rect 488316 153456 488322 153468
rect 490466 153456 490472 153468
rect 488316 153428 490472 153456
rect 488316 153416 488322 153428
rect 490466 153416 490472 153428
rect 490524 153416 490530 153468
rect 514846 153416 514852 153468
rect 514904 153456 514910 153468
rect 518894 153456 518900 153468
rect 514904 153428 518900 153456
rect 514904 153416 514910 153428
rect 518894 153416 518900 153428
rect 518952 153416 518958 153468
rect 50614 153348 50620 153400
rect 50672 153388 50678 153400
rect 115290 153388 115296 153400
rect 50672 153360 115296 153388
rect 50672 153348 50678 153360
rect 115290 153348 115296 153360
rect 115348 153348 115354 153400
rect 459554 153348 459560 153400
rect 459612 153388 459618 153400
rect 462866 153388 462872 153400
rect 459612 153360 462872 153388
rect 459612 153348 459618 153360
rect 462866 153348 462872 153360
rect 462924 153348 462930 153400
rect 468110 153348 468116 153400
rect 468168 153388 468174 153400
rect 473078 153388 473084 153400
rect 468168 153360 473084 153388
rect 468168 153348 468174 153360
rect 473078 153348 473084 153360
rect 473136 153348 473142 153400
rect 488534 153348 488540 153400
rect 488592 153388 488598 153400
rect 491754 153388 491760 153400
rect 488592 153360 491760 153388
rect 488592 153348 488598 153360
rect 491754 153348 491760 153360
rect 491812 153348 491818 153400
rect 516134 153348 516140 153400
rect 516192 153388 516198 153400
rect 520734 153388 520740 153400
rect 516192 153360 520740 153388
rect 516192 153348 516198 153360
rect 520734 153348 520740 153360
rect 520792 153348 520798 153400
rect 522574 153348 522580 153400
rect 522632 153388 522638 153400
rect 529934 153388 529940 153400
rect 522632 153360 529940 153388
rect 522632 153348 522638 153360
rect 529934 153348 529940 153360
rect 529992 153348 529998 153400
rect 46750 153280 46756 153332
rect 46808 153320 46814 153332
rect 117222 153320 117228 153332
rect 46808 153292 117228 153320
rect 46808 153280 46814 153292
rect 117222 153280 117228 153292
rect 117280 153280 117286 153332
rect 379514 153280 379520 153332
rect 379572 153320 379578 153332
rect 385770 153320 385776 153332
rect 379572 153292 385776 153320
rect 379572 153280 379578 153292
rect 385770 153280 385776 153292
rect 385828 153280 385834 153332
rect 459830 153280 459836 153332
rect 459888 153320 459894 153332
rect 462222 153320 462228 153332
rect 459888 153292 462228 153320
rect 459888 153280 459894 153292
rect 462222 153280 462228 153292
rect 462280 153280 462286 153332
rect 468202 153280 468208 153332
rect 468260 153320 468266 153332
rect 472434 153320 472440 153332
rect 468260 153292 472440 153320
rect 468260 153280 468266 153292
rect 472434 153280 472440 153292
rect 472492 153280 472498 153332
rect 478874 153280 478880 153332
rect 478932 153320 478938 153332
rect 481450 153320 481456 153332
rect 478932 153292 481456 153320
rect 478932 153280 478938 153292
rect 481450 153280 481456 153292
rect 481508 153280 481514 153332
rect 521930 153280 521936 153332
rect 521988 153320 521994 153332
rect 528554 153320 528560 153332
rect 521988 153292 528560 153320
rect 521988 153280 521994 153292
rect 528554 153280 528560 153292
rect 528612 153280 528618 153332
rect 108942 153212 108948 153264
rect 109000 153252 109006 153264
rect 119890 153252 119896 153264
rect 109000 153224 119896 153252
rect 109000 153212 109006 153224
rect 119890 153212 119896 153224
rect 119948 153212 119954 153264
rect 277228 153224 277394 153252
rect 114646 153144 114652 153196
rect 114704 153184 114710 153196
rect 182910 153184 182916 153196
rect 114704 153156 182916 153184
rect 114704 153144 114710 153156
rect 182910 153144 182916 153156
rect 182968 153144 182974 153196
rect 184106 153144 184112 153196
rect 184164 153184 184170 153196
rect 266354 153184 266360 153196
rect 184164 153156 266360 153184
rect 184164 153144 184170 153156
rect 266354 153144 266360 153156
rect 266412 153144 266418 153196
rect 274542 153144 274548 153196
rect 274600 153184 274606 153196
rect 277228 153184 277256 153224
rect 274600 153156 277256 153184
rect 277366 153184 277394 153224
rect 310238 153212 310244 153264
rect 310296 153252 310302 153264
rect 317046 153252 317052 153264
rect 310296 153224 317052 153252
rect 310296 153212 310302 153224
rect 317046 153212 317052 153224
rect 317104 153212 317110 153264
rect 382274 153212 382280 153264
rect 382332 153252 382338 153264
rect 383838 153252 383844 153264
rect 382332 153224 383844 153252
rect 382332 153212 382338 153224
rect 383838 153212 383844 153224
rect 383896 153212 383902 153264
rect 420914 153212 420920 153264
rect 420972 153252 420978 153264
rect 422386 153252 422392 153264
rect 420972 153224 422392 153252
rect 420972 153212 420978 153224
rect 422386 153212 422392 153224
rect 422444 153212 422450 153264
rect 429194 153212 429200 153264
rect 429252 153252 429258 153264
rect 433978 153252 433984 153264
rect 429252 153224 433984 153252
rect 429252 153212 429258 153224
rect 433978 153212 433984 153224
rect 434036 153212 434042 153264
rect 440234 153212 440240 153264
rect 440292 153252 440298 153264
rect 441614 153252 441620 153264
rect 440292 153224 441620 153252
rect 440292 153212 440298 153224
rect 441614 153212 441620 153224
rect 441672 153212 441678 153264
rect 449894 153212 449900 153264
rect 449952 153252 449958 153264
rect 451918 153252 451924 153264
rect 449952 153224 451924 153252
rect 449952 153212 449958 153224
rect 451918 153212 451924 153224
rect 451976 153212 451982 153264
rect 458174 153212 458180 153264
rect 458232 153252 458238 153264
rect 461578 153252 461584 153264
rect 458232 153224 461584 153252
rect 458232 153212 458238 153224
rect 461578 153212 461584 153224
rect 461636 153212 461642 153264
rect 476390 153212 476396 153264
rect 476448 153252 476454 153264
rect 476448 153224 478920 153252
rect 476448 153212 476454 153224
rect 478892 153196 478920 153224
rect 478966 153212 478972 153264
rect 479024 153252 479030 153264
rect 480806 153252 480812 153264
rect 479024 153224 480812 153252
rect 479024 153212 479030 153224
rect 480806 153212 480812 153224
rect 480864 153212 480870 153264
rect 488626 153212 488632 153264
rect 488684 153252 488690 153264
rect 491110 153252 491116 153264
rect 488684 153224 491116 153252
rect 488684 153212 488690 153224
rect 491110 153212 491116 153224
rect 491168 153212 491174 153264
rect 516778 153212 516784 153264
rect 516836 153252 516842 153264
rect 520550 153252 520556 153264
rect 516836 153224 520556 153252
rect 516836 153212 516842 153224
rect 520550 153212 520556 153224
rect 520608 153212 520614 153264
rect 333146 153184 333152 153196
rect 277366 153156 333152 153184
rect 274600 153144 274606 153156
rect 333146 153144 333152 153156
rect 333204 153144 333210 153196
rect 478874 153144 478880 153196
rect 478932 153144 478938 153196
rect 118694 153076 118700 153128
rect 118752 153116 118758 153128
rect 175826 153116 175832 153128
rect 118752 153088 175832 153116
rect 118752 153076 118758 153088
rect 175826 153076 175832 153088
rect 175884 153076 175890 153128
rect 177206 153076 177212 153128
rect 177264 153116 177270 153128
rect 261202 153116 261208 153128
rect 177264 153088 261208 153116
rect 177264 153076 177270 153088
rect 261202 153076 261208 153088
rect 261260 153076 261266 153128
rect 272245 153119 272303 153125
rect 272245 153085 272257 153119
rect 272291 153116 272303 153119
rect 324130 153116 324136 153128
rect 272291 153088 324136 153116
rect 272291 153085 272303 153088
rect 272245 153079 272303 153085
rect 324130 153076 324136 153088
rect 324188 153076 324194 153128
rect 62114 153008 62120 153060
rect 62172 153048 62178 153060
rect 146294 153048 146300 153060
rect 62172 153020 146300 153048
rect 62172 153008 62178 153020
rect 146294 153008 146300 153020
rect 146352 153008 146358 153060
rect 250717 153051 250775 153057
rect 250717 153017 250729 153051
rect 250763 153048 250775 153051
rect 250763 153020 306374 153048
rect 250763 153017 250775 153020
rect 250717 153011 250775 153017
rect 143258 152940 143264 152992
rect 143316 152980 143322 152992
rect 235534 152980 235540 152992
rect 143316 152952 235540 152980
rect 143316 152940 143322 152952
rect 235534 152940 235540 152952
rect 235592 152940 235598 152992
rect 236086 152940 236092 152992
rect 236144 152980 236150 152992
rect 304902 152980 304908 152992
rect 236144 152952 304908 152980
rect 236144 152940 236150 152952
rect 304902 152940 304908 152952
rect 304960 152940 304966 152992
rect 222286 152872 222292 152924
rect 222344 152912 222350 152924
rect 222344 152884 229094 152912
rect 222344 152872 222350 152884
rect 125502 152804 125508 152856
rect 125560 152844 125566 152856
rect 222654 152844 222660 152856
rect 125560 152816 222660 152844
rect 125560 152804 125566 152816
rect 222654 152804 222660 152816
rect 222712 152804 222718 152856
rect 229066 152844 229094 152884
rect 229186 152872 229192 152924
rect 229244 152912 229250 152924
rect 299750 152912 299756 152924
rect 229244 152884 299756 152912
rect 229244 152872 229250 152884
rect 299750 152872 299756 152884
rect 299808 152872 299814 152924
rect 306346 152912 306374 153020
rect 308766 152912 308772 152924
rect 306346 152884 308772 152912
rect 308766 152872 308772 152884
rect 308824 152872 308830 152924
rect 294598 152844 294604 152856
rect 229066 152816 294604 152844
rect 294598 152804 294604 152816
rect 294656 152804 294662 152856
rect 118602 152736 118608 152788
rect 118660 152776 118666 152788
rect 217594 152776 217600 152788
rect 118660 152748 217600 152776
rect 118660 152736 118666 152748
rect 217594 152736 217600 152748
rect 217652 152736 217658 152788
rect 218790 152736 218796 152788
rect 218848 152776 218854 152788
rect 292022 152776 292028 152788
rect 218848 152748 292028 152776
rect 218848 152736 218854 152748
rect 292022 152736 292028 152748
rect 292080 152736 292086 152788
rect 111702 152668 111708 152720
rect 111760 152708 111766 152720
rect 212442 152708 212448 152720
rect 111760 152680 212448 152708
rect 111760 152668 111766 152680
rect 212442 152668 212448 152680
rect 212500 152668 212506 152720
rect 215294 152668 215300 152720
rect 215352 152708 215358 152720
rect 289446 152708 289452 152720
rect 215352 152680 289452 152708
rect 215352 152668 215358 152680
rect 289446 152668 289452 152680
rect 289504 152668 289510 152720
rect 93946 152600 93952 152652
rect 94004 152640 94010 152652
rect 199562 152640 199568 152652
rect 94004 152612 199568 152640
rect 94004 152600 94010 152612
rect 199562 152600 199568 152612
rect 199620 152600 199626 152652
rect 208394 152600 208400 152652
rect 208452 152640 208458 152652
rect 284294 152640 284300 152652
rect 208452 152612 284300 152640
rect 208452 152600 208458 152612
rect 284294 152600 284300 152612
rect 284352 152600 284358 152652
rect 87046 152532 87052 152584
rect 87104 152572 87110 152584
rect 194410 152572 194416 152584
rect 87104 152544 194416 152572
rect 87104 152532 87110 152544
rect 194410 152532 194416 152544
rect 194468 152532 194474 152584
rect 197998 152532 198004 152584
rect 198056 152572 198062 152584
rect 276658 152572 276664 152584
rect 198056 152544 276664 152572
rect 198056 152532 198062 152544
rect 276658 152532 276664 152544
rect 276716 152532 276722 152584
rect 279418 152532 279424 152584
rect 279476 152572 279482 152584
rect 337010 152572 337016 152584
rect 279476 152544 337016 152572
rect 279476 152532 279482 152544
rect 337010 152532 337016 152544
rect 337068 152532 337074 152584
rect 2958 152464 2964 152516
rect 3016 152504 3022 152516
rect 132126 152504 132132 152516
rect 3016 152476 132132 152504
rect 3016 152464 3022 152476
rect 132126 152464 132132 152476
rect 132184 152464 132190 152516
rect 227714 152464 227720 152516
rect 227772 152504 227778 152516
rect 298462 152504 298468 152516
rect 227772 152476 298468 152504
rect 227772 152464 227778 152476
rect 298462 152464 298468 152476
rect 298520 152464 298526 152516
rect 151998 152396 152004 152448
rect 152056 152436 152062 152448
rect 242618 152436 242624 152448
rect 152056 152408 242624 152436
rect 152056 152396 152062 152408
rect 242618 152396 242624 152408
rect 242676 152396 242682 152448
rect 262214 152396 262220 152448
rect 262272 152436 262278 152448
rect 272245 152439 272303 152445
rect 272245 152436 272257 152439
rect 262272 152408 272257 152436
rect 262272 152396 262278 152408
rect 272245 152405 272257 152408
rect 272291 152405 272303 152439
rect 272245 152399 272303 152405
rect 132954 152328 132960 152380
rect 133012 152368 133018 152380
rect 228450 152368 228456 152380
rect 133012 152340 228456 152368
rect 133012 152328 133018 152340
rect 228450 152328 228456 152340
rect 228508 152328 228514 152380
rect 241514 152328 241520 152380
rect 241572 152368 241578 152380
rect 250717 152371 250775 152377
rect 250717 152368 250729 152371
rect 241572 152340 250729 152368
rect 241572 152328 241578 152340
rect 250717 152337 250729 152340
rect 250763 152337 250775 152371
rect 250717 152331 250775 152337
rect 16206 152260 16212 152312
rect 16264 152300 16270 152312
rect 124858 152300 124864 152312
rect 16264 152272 124864 152300
rect 16264 152260 16270 152272
rect 124858 152260 124864 152272
rect 124916 152260 124922 152312
rect 135530 152260 135536 152312
rect 135588 152300 135594 152312
rect 230382 152300 230388 152312
rect 135588 152272 230388 152300
rect 135588 152260 135594 152272
rect 230382 152260 230388 152272
rect 230440 152260 230446 152312
rect 101904 152192 101910 152244
rect 101962 152232 101968 152244
rect 118602 152232 118608 152244
rect 101962 152204 118608 152232
rect 101962 152192 101968 152204
rect 118602 152192 118608 152204
rect 118660 152192 118666 152244
rect 91600 152124 91606 152176
rect 91658 152164 91664 152176
rect 116578 152164 116584 152176
rect 91658 152136 116584 152164
rect 91658 152124 91664 152136
rect 116578 152124 116584 152136
rect 116636 152124 116642 152176
rect 39988 152056 39994 152108
rect 40046 152096 40052 152108
rect 115198 152096 115204 152108
rect 40046 152068 115204 152096
rect 40046 152056 40052 152068
rect 115198 152056 115204 152068
rect 115256 152056 115262 152108
rect 36906 151988 36912 152040
rect 36964 152028 36970 152040
rect 120810 152028 120816 152040
rect 36964 152000 120816 152028
rect 36964 151988 36970 152000
rect 120810 151988 120816 152000
rect 120868 151988 120874 152040
rect 30006 151920 30012 151972
rect 30064 151960 30070 151972
rect 122190 151960 122196 151972
rect 30064 151932 122196 151960
rect 30064 151920 30070 151932
rect 122190 151920 122196 151932
rect 122248 151920 122254 151972
rect 19702 151852 19708 151904
rect 19760 151892 19766 151904
rect 123478 151892 123484 151904
rect 19760 151864 123484 151892
rect 19760 151852 19766 151864
rect 123478 151852 123484 151864
rect 123536 151852 123542 151904
rect 105630 151784 105636 151836
rect 105688 151824 105694 151836
rect 114554 151824 114560 151836
rect 105688 151796 114560 151824
rect 105688 151784 105694 151796
rect 114554 151784 114560 151796
rect 114612 151784 114618 151836
rect 531590 151512 531596 151564
rect 531648 151552 531654 151564
rect 534718 151552 534724 151564
rect 531648 151524 534724 151552
rect 531648 151512 531654 151524
rect 534718 151512 534724 151524
rect 534776 151512 534782 151564
rect 60826 151416 60832 151428
rect 60787 151388 60832 151416
rect 60826 151376 60832 151388
rect 60884 151376 60890 151428
rect 64414 151416 64420 151428
rect 64375 151388 64420 151416
rect 64414 151376 64420 151388
rect 64472 151376 64478 151428
rect 53926 151308 53932 151360
rect 53984 151308 53990 151360
rect 57514 151308 57520 151360
rect 57572 151348 57578 151360
rect 67634 151348 67640 151360
rect 57572 151320 64874 151348
rect 67595 151320 67640 151348
rect 57572 151308 57578 151320
rect 53944 151212 53972 151308
rect 64846 151280 64874 151320
rect 67634 151308 67640 151320
rect 67692 151308 67698 151360
rect 71314 151348 71320 151360
rect 71275 151320 71320 151348
rect 71314 151308 71320 151320
rect 71372 151308 71378 151360
rect 74534 151308 74540 151360
rect 74592 151348 74598 151360
rect 78122 151348 78128 151360
rect 74592 151320 74637 151348
rect 78083 151320 78128 151348
rect 74592 151308 74598 151320
rect 78122 151308 78128 151320
rect 78180 151308 78186 151360
rect 81434 151348 81440 151360
rect 81395 151320 81440 151348
rect 81434 151308 81440 151320
rect 81492 151308 81498 151360
rect 85022 151348 85028 151360
rect 84983 151320 85028 151348
rect 85022 151308 85028 151320
rect 85080 151308 85086 151360
rect 88334 151348 88340 151360
rect 88295 151320 88340 151348
rect 88334 151308 88340 151320
rect 88392 151308 88398 151360
rect 98822 151348 98828 151360
rect 98783 151320 98828 151348
rect 98822 151308 98828 151320
rect 98880 151308 98886 151360
rect 116854 151280 116860 151292
rect 64846 151252 116860 151280
rect 116854 151240 116860 151252
rect 116912 151240 116918 151292
rect 123570 151212 123576 151224
rect 53944 151184 123576 151212
rect 123570 151172 123576 151184
rect 123628 151172 123634 151224
rect 88337 151147 88395 151153
rect 88337 151113 88349 151147
rect 88383 151144 88395 151147
rect 115382 151144 115388 151156
rect 88383 151116 115388 151144
rect 88383 151113 88395 151116
rect 88337 151107 88395 151113
rect 115382 151104 115388 151116
rect 115440 151104 115446 151156
rect 120718 151104 120724 151156
rect 120776 151144 120782 151156
rect 127618 151144 127624 151156
rect 120776 151116 127624 151144
rect 120776 151104 120782 151116
rect 127618 151104 127624 151116
rect 127676 151104 127682 151156
rect 85025 151079 85083 151085
rect 85025 151045 85037 151079
rect 85071 151076 85083 151079
rect 123662 151076 123668 151088
rect 85071 151048 123668 151076
rect 85071 151045 85083 151048
rect 85025 151039 85083 151045
rect 123662 151036 123668 151048
rect 123720 151036 123726 151088
rect 81437 151011 81495 151017
rect 81437 150977 81449 151011
rect 81483 151008 81495 151011
rect 122282 151008 122288 151020
rect 81483 150980 122288 151008
rect 81483 150977 81495 150980
rect 81437 150971 81495 150977
rect 122282 150968 122288 150980
rect 122340 150968 122346 151020
rect 78125 150943 78183 150949
rect 78125 150909 78137 150943
rect 78171 150940 78183 150943
rect 119522 150940 119528 150952
rect 78171 150912 119528 150940
rect 78171 150909 78183 150912
rect 78125 150903 78183 150909
rect 119522 150900 119528 150912
rect 119580 150900 119586 150952
rect 74537 150875 74595 150881
rect 74537 150841 74549 150875
rect 74583 150872 74595 150875
rect 116762 150872 116768 150884
rect 74583 150844 116768 150872
rect 74583 150841 74595 150844
rect 74537 150835 74595 150841
rect 116762 150832 116768 150844
rect 116820 150832 116826 150884
rect 71317 150807 71375 150813
rect 71317 150773 71329 150807
rect 71363 150804 71375 150807
rect 118142 150804 118148 150816
rect 71363 150776 118148 150804
rect 71363 150773 71375 150776
rect 71317 150767 71375 150773
rect 118142 150764 118148 150776
rect 118200 150764 118206 150816
rect 67637 150739 67695 150745
rect 67637 150705 67649 150739
rect 67683 150736 67695 150739
rect 120902 150736 120908 150748
rect 67683 150708 120908 150736
rect 67683 150705 67695 150708
rect 67637 150699 67695 150705
rect 120902 150696 120908 150708
rect 120960 150696 120966 150748
rect 112530 150628 112536 150680
rect 112588 150668 112594 150680
rect 126974 150668 126980 150680
rect 112588 150640 126980 150668
rect 112588 150628 112594 150640
rect 126974 150628 126980 150640
rect 127032 150628 127038 150680
rect 64417 150603 64475 150609
rect 64417 150569 64429 150603
rect 64463 150600 64475 150603
rect 126330 150600 126336 150612
rect 64463 150572 126336 150600
rect 64463 150569 64475 150572
rect 64417 150563 64475 150569
rect 126330 150560 126336 150572
rect 126388 150560 126394 150612
rect 60829 150535 60887 150541
rect 60829 150501 60841 150535
rect 60875 150532 60887 150535
rect 124950 150532 124956 150544
rect 60875 150504 124956 150532
rect 60875 150501 60887 150504
rect 60829 150495 60887 150501
rect 124950 150492 124956 150504
rect 125008 150492 125014 150544
rect 98825 150467 98883 150473
rect 98825 150433 98837 150467
rect 98871 150464 98883 150467
rect 124582 150464 124588 150476
rect 98871 150436 124588 150464
rect 98871 150433 98883 150436
rect 98825 150427 98883 150433
rect 124582 150424 124588 150436
rect 124640 150424 124646 150476
rect 126698 150424 126704 150476
rect 126756 150464 126762 150476
rect 127894 150464 127900 150476
rect 126756 150436 127900 150464
rect 126756 150424 126762 150436
rect 127894 150424 127900 150436
rect 127952 150424 127958 150476
rect 532602 149880 532608 149932
rect 532660 149920 532666 149932
rect 536098 149920 536104 149932
rect 532660 149892 536104 149920
rect 532660 149880 532666 149892
rect 536098 149880 536104 149892
rect 536156 149880 536162 149932
rect 117222 149676 117228 149728
rect 117280 149716 117286 149728
rect 127710 149716 127716 149728
rect 117280 149688 127716 149716
rect 117280 149676 117286 149688
rect 127710 149676 127716 149688
rect 127768 149676 127774 149728
rect 119890 148996 119896 149048
rect 119948 149036 119954 149048
rect 126974 149036 126980 149048
rect 119948 149008 126980 149036
rect 119948 148996 119954 149008
rect 126974 148996 126980 149008
rect 127032 148996 127038 149048
rect 532326 148996 532332 149048
rect 532384 149036 532390 149048
rect 536190 149036 536196 149048
rect 532384 149008 536196 149036
rect 532384 148996 532390 149008
rect 536190 148996 536196 149008
rect 536248 148996 536254 149048
rect 114554 147568 114560 147620
rect 114612 147608 114618 147620
rect 126974 147608 126980 147620
rect 114612 147580 126980 147608
rect 114612 147568 114618 147580
rect 126974 147568 126980 147580
rect 127032 147568 127038 147620
rect 118602 146208 118608 146260
rect 118660 146248 118666 146260
rect 126974 146248 126980 146260
rect 118660 146220 126980 146248
rect 118660 146208 118666 146220
rect 126974 146208 126980 146220
rect 127032 146208 127038 146260
rect 532142 146072 532148 146124
rect 532200 146112 532206 146124
rect 535362 146112 535368 146124
rect 532200 146084 535368 146112
rect 532200 146072 532206 146084
rect 535362 146072 535368 146084
rect 535420 146072 535426 146124
rect 116670 145188 116676 145240
rect 116728 145228 116734 145240
rect 120718 145228 120724 145240
rect 116728 145200 120724 145228
rect 116728 145188 116734 145200
rect 120718 145188 120724 145200
rect 120776 145188 120782 145240
rect 531774 144848 531780 144900
rect 531832 144888 531838 144900
rect 536282 144888 536288 144900
rect 531832 144860 536288 144888
rect 531832 144848 531838 144860
rect 536282 144848 536288 144860
rect 536340 144848 536346 144900
rect 124582 143488 124588 143540
rect 124640 143528 124646 143540
rect 126974 143528 126980 143540
rect 124640 143500 126980 143528
rect 124640 143488 124646 143500
rect 126974 143488 126980 143500
rect 127032 143488 127038 143540
rect 531682 143216 531688 143268
rect 531740 143256 531746 143268
rect 535270 143256 535276 143268
rect 531740 143228 535276 143256
rect 531740 143216 531746 143228
rect 535270 143216 535276 143228
rect 535328 143216 535334 143268
rect 531958 141856 531964 141908
rect 532016 141896 532022 141908
rect 534902 141896 534908 141908
rect 532016 141868 534908 141896
rect 532016 141856 532022 141868
rect 534902 141856 534908 141868
rect 534960 141856 534966 141908
rect 116578 140700 116584 140752
rect 116636 140740 116642 140752
rect 126974 140740 126980 140752
rect 116636 140712 126980 140740
rect 116636 140700 116642 140712
rect 126974 140700 126980 140712
rect 127032 140700 127038 140752
rect 531958 140700 531964 140752
rect 532016 140740 532022 140752
rect 535178 140740 535184 140752
rect 532016 140712 535184 140740
rect 532016 140700 532022 140712
rect 535178 140700 535184 140712
rect 535236 140700 535242 140752
rect 531590 139340 531596 139392
rect 531648 139380 531654 139392
rect 534718 139380 534724 139392
rect 531648 139352 534724 139380
rect 531648 139340 531654 139352
rect 534718 139340 534724 139352
rect 534776 139340 534782 139392
rect 115382 137912 115388 137964
rect 115440 137952 115446 137964
rect 126974 137952 126980 137964
rect 115440 137924 126980 137952
rect 115440 137912 115446 137924
rect 126974 137912 126980 137924
rect 127032 137912 127038 137964
rect 531406 137912 531412 137964
rect 531464 137952 531470 137964
rect 534810 137952 534816 137964
rect 531464 137924 534816 137952
rect 531464 137912 531470 137924
rect 534810 137912 534816 137924
rect 534868 137912 534874 137964
rect 123662 136552 123668 136604
rect 123720 136592 123726 136604
rect 126974 136592 126980 136604
rect 123720 136564 126980 136592
rect 123720 136552 123726 136564
rect 126974 136552 126980 136564
rect 127032 136552 127038 136604
rect 532142 136348 532148 136400
rect 532200 136388 532206 136400
rect 535086 136388 535092 136400
rect 532200 136360 535092 136388
rect 532200 136348 532206 136360
rect 535086 136348 535092 136360
rect 535144 136348 535150 136400
rect 531774 134852 531780 134904
rect 531832 134892 531838 134904
rect 534994 134892 535000 134904
rect 531832 134864 535000 134892
rect 531832 134852 531838 134864
rect 534994 134852 535000 134864
rect 535052 134852 535058 134904
rect 122282 133832 122288 133884
rect 122340 133872 122346 133884
rect 126974 133872 126980 133884
rect 122340 133844 126980 133872
rect 122340 133832 122346 133844
rect 126974 133832 126980 133844
rect 127032 133832 127038 133884
rect 531774 133492 531780 133544
rect 531832 133532 531838 133544
rect 536190 133532 536196 133544
rect 531832 133504 536196 133532
rect 531832 133492 531838 133504
rect 536190 133492 536196 133504
rect 536248 133492 536254 133544
rect 119522 132404 119528 132456
rect 119580 132444 119586 132456
rect 126974 132444 126980 132456
rect 119580 132416 126980 132444
rect 119580 132404 119586 132416
rect 126974 132404 126980 132416
rect 127032 132404 127038 132456
rect 531406 131996 531412 132048
rect 531464 132036 531470 132048
rect 536006 132036 536012 132048
rect 531464 132008 536012 132036
rect 531464 131996 531470 132008
rect 536006 131996 536012 132008
rect 536064 131996 536070 132048
rect 116670 131044 116676 131096
rect 116728 131084 116734 131096
rect 126974 131084 126980 131096
rect 116728 131056 126980 131084
rect 116728 131044 116734 131056
rect 126974 131044 126980 131056
rect 127032 131044 127038 131096
rect 532602 130636 532608 130688
rect 532660 130676 532666 130688
rect 536742 130676 536748 130688
rect 532660 130648 536748 130676
rect 532660 130636 532666 130648
rect 536742 130636 536748 130648
rect 536800 130636 536806 130688
rect 531590 129412 531596 129464
rect 531648 129452 531654 129464
rect 536650 129452 536656 129464
rect 531648 129424 536656 129452
rect 531648 129412 531654 129424
rect 536650 129412 536656 129424
rect 536708 129412 536714 129464
rect 118142 128256 118148 128308
rect 118200 128296 118206 128308
rect 126974 128296 126980 128308
rect 118200 128268 126980 128296
rect 118200 128256 118206 128268
rect 126974 128256 126980 128268
rect 127032 128256 127038 128308
rect 531958 128052 531964 128104
rect 532016 128092 532022 128104
rect 536558 128092 536564 128104
rect 532016 128064 536564 128092
rect 532016 128052 532022 128064
rect 536558 128052 536564 128064
rect 536616 128052 536622 128104
rect 120902 126896 120908 126948
rect 120960 126936 120966 126948
rect 126974 126936 126980 126948
rect 120960 126908 126980 126936
rect 120960 126896 120966 126908
rect 126974 126896 126980 126908
rect 127032 126896 127038 126948
rect 531866 126556 531872 126608
rect 531924 126596 531930 126608
rect 536466 126596 536472 126608
rect 531924 126568 536472 126596
rect 531924 126556 531930 126568
rect 536466 126556 536472 126568
rect 536524 126556 536530 126608
rect 532602 125196 532608 125248
rect 532660 125236 532666 125248
rect 536374 125236 536380 125248
rect 532660 125208 536380 125236
rect 532660 125196 532666 125208
rect 536374 125196 536380 125208
rect 536432 125196 536438 125248
rect 531774 123836 531780 123888
rect 531832 123876 531838 123888
rect 536098 123876 536104 123888
rect 531832 123848 536104 123876
rect 531832 123836 531838 123848
rect 536098 123836 536104 123848
rect 536156 123836 536162 123888
rect 532602 122476 532608 122528
rect 532660 122516 532666 122528
rect 536282 122516 536288 122528
rect 532660 122488 536288 122516
rect 532660 122476 532666 122488
rect 536282 122476 536288 122488
rect 536340 122476 536346 122528
rect 124950 122408 124956 122460
rect 125008 122448 125014 122460
rect 126974 122448 126980 122460
rect 125008 122420 126980 122448
rect 125008 122408 125014 122420
rect 126974 122408 126980 122420
rect 127032 122408 127038 122460
rect 116762 121388 116768 121440
rect 116820 121428 116826 121440
rect 126974 121428 126980 121440
rect 116820 121400 126980 121428
rect 116820 121388 116826 121400
rect 126974 121388 126980 121400
rect 127032 121388 127038 121440
rect 532142 121116 532148 121168
rect 532200 121156 532206 121168
rect 536190 121156 536196 121168
rect 532200 121128 536196 121156
rect 532200 121116 532206 121128
rect 536190 121116 536196 121128
rect 536248 121116 536254 121168
rect 532510 119892 532516 119944
rect 532568 119932 532574 119944
rect 536650 119932 536656 119944
rect 532568 119904 536656 119932
rect 532568 119892 532574 119904
rect 536650 119892 536656 119904
rect 536708 119892 536714 119944
rect 123570 118600 123576 118652
rect 123628 118640 123634 118652
rect 126974 118640 126980 118652
rect 123628 118612 126980 118640
rect 123628 118600 123634 118612
rect 126974 118600 126980 118612
rect 127032 118600 127038 118652
rect 532602 118396 532608 118448
rect 532660 118436 532666 118448
rect 536742 118436 536748 118448
rect 532660 118408 536748 118436
rect 532660 118396 532666 118408
rect 536742 118396 536748 118408
rect 536800 118396 536806 118448
rect 115290 117240 115296 117292
rect 115348 117280 115354 117292
rect 126974 117280 126980 117292
rect 115348 117252 126980 117280
rect 115348 117240 115354 117252
rect 126974 117240 126980 117252
rect 127032 117240 127038 117292
rect 532326 117036 532332 117088
rect 532384 117076 532390 117088
rect 535454 117076 535460 117088
rect 532384 117048 535460 117076
rect 532384 117036 532390 117048
rect 535454 117036 535460 117048
rect 535512 117036 535518 117088
rect 532602 115676 532608 115728
rect 532660 115716 532666 115728
rect 536374 115716 536380 115728
rect 532660 115688 536380 115716
rect 532660 115676 532666 115688
rect 536374 115676 536380 115688
rect 536432 115676 536438 115728
rect 531682 114316 531688 114368
rect 531740 114356 531746 114368
rect 535638 114356 535644 114368
rect 531740 114328 535644 114356
rect 531740 114316 531746 114328
rect 535638 114316 535644 114328
rect 535696 114316 535702 114368
rect 118050 113092 118056 113144
rect 118108 113132 118114 113144
rect 126974 113132 126980 113144
rect 118108 113104 126980 113132
rect 118108 113092 118114 113104
rect 126974 113092 126980 113104
rect 127032 113092 127038 113144
rect 531774 112888 531780 112940
rect 531832 112928 531838 112940
rect 536282 112928 536288 112940
rect 531832 112900 536288 112928
rect 531832 112888 531838 112900
rect 536282 112888 536288 112900
rect 536340 112888 536346 112940
rect 532510 111800 532516 111852
rect 532568 111840 532574 111852
rect 535454 111840 535460 111852
rect 532568 111812 535460 111840
rect 532568 111800 532574 111812
rect 535454 111800 535460 111812
rect 535512 111800 535518 111852
rect 115198 111732 115204 111784
rect 115256 111772 115262 111784
rect 126974 111772 126980 111784
rect 115256 111744 126980 111772
rect 115256 111732 115262 111744
rect 126974 111732 126980 111744
rect 127032 111732 127038 111784
rect 532602 111460 532608 111512
rect 532660 111500 532666 111512
rect 536466 111500 536472 111512
rect 532660 111472 536472 111500
rect 532660 111460 532666 111472
rect 536466 111460 536472 111472
rect 536524 111460 536530 111512
rect 532602 110440 532608 110492
rect 532660 110480 532666 110492
rect 535454 110480 535460 110492
rect 532660 110452 535460 110480
rect 532660 110440 532666 110452
rect 535454 110440 535460 110452
rect 535512 110440 535518 110492
rect 531958 110100 531964 110152
rect 532016 110140 532022 110152
rect 536190 110140 536196 110152
rect 532016 110112 536196 110140
rect 532016 110100 532022 110112
rect 536190 110100 536196 110112
rect 536248 110100 536254 110152
rect 532418 109012 532424 109064
rect 532476 109052 532482 109064
rect 535454 109052 535460 109064
rect 532476 109024 535460 109052
rect 532476 109012 532482 109024
rect 535454 109012 535460 109024
rect 535512 109012 535518 109064
rect 120810 108944 120816 108996
rect 120868 108984 120874 108996
rect 126974 108984 126980 108996
rect 120868 108956 126980 108984
rect 120868 108944 120874 108956
rect 126974 108944 126980 108956
rect 127032 108944 127038 108996
rect 531774 108876 531780 108928
rect 531832 108916 531838 108928
rect 536650 108916 536656 108928
rect 531832 108888 536656 108916
rect 531832 108876 531838 108888
rect 536650 108876 536656 108888
rect 536708 108876 536714 108928
rect 532234 107652 532240 107704
rect 532292 107692 532298 107704
rect 535454 107692 535460 107704
rect 532292 107664 535460 107692
rect 532292 107652 532298 107664
rect 535454 107652 535460 107664
rect 535512 107652 535518 107704
rect 119430 107584 119436 107636
rect 119488 107624 119494 107636
rect 126974 107624 126980 107636
rect 119488 107596 126980 107624
rect 119488 107584 119494 107596
rect 126974 107584 126980 107596
rect 127032 107584 127038 107636
rect 531774 107380 531780 107432
rect 531832 107420 531838 107432
rect 535546 107420 535552 107432
rect 531832 107392 535552 107420
rect 531832 107380 531838 107392
rect 535546 107380 535552 107392
rect 535604 107380 535610 107432
rect 532142 106292 532148 106344
rect 532200 106332 532206 106344
rect 535454 106332 535460 106344
rect 532200 106304 535460 106332
rect 532200 106292 532206 106304
rect 535454 106292 535460 106304
rect 535512 106292 535518 106344
rect 532510 104864 532516 104916
rect 532568 104904 532574 104916
rect 535454 104904 535460 104916
rect 532568 104876 535460 104904
rect 532568 104864 532574 104876
rect 535454 104864 535460 104876
rect 535512 104864 535518 104916
rect 122190 104796 122196 104848
rect 122248 104836 122254 104848
rect 126974 104836 126980 104848
rect 122248 104808 126980 104836
rect 122248 104796 122254 104808
rect 126974 104796 126980 104808
rect 127032 104796 127038 104848
rect 532602 103708 532608 103760
rect 532660 103748 532666 103760
rect 535454 103748 535460 103760
rect 532660 103720 535460 103748
rect 532660 103708 532666 103720
rect 535454 103708 535460 103720
rect 535512 103708 535518 103760
rect 117958 103436 117964 103488
rect 118016 103476 118022 103488
rect 126974 103476 126980 103488
rect 118016 103448 126980 103476
rect 118016 103436 118022 103448
rect 126974 103436 126980 103448
rect 127032 103436 127038 103488
rect 532050 102144 532056 102196
rect 532108 102184 532114 102196
rect 535454 102184 535460 102196
rect 532108 102156 535460 102184
rect 532108 102144 532114 102156
rect 535454 102144 535460 102156
rect 535512 102144 535518 102196
rect 122098 102076 122104 102128
rect 122156 102116 122162 102128
rect 126974 102116 126980 102128
rect 122156 102088 126980 102116
rect 122156 102076 122162 102088
rect 126974 102076 126980 102088
rect 127032 102076 127038 102128
rect 532602 100716 532608 100768
rect 532660 100756 532666 100768
rect 535454 100756 535460 100768
rect 532660 100728 535460 100756
rect 532660 100716 532666 100728
rect 535454 100716 535460 100728
rect 535512 100716 535518 100768
rect 116946 99424 116952 99476
rect 117004 99464 117010 99476
rect 122098 99464 122104 99476
rect 117004 99436 122104 99464
rect 117004 99424 117010 99436
rect 122098 99424 122104 99436
rect 122156 99424 122162 99476
rect 123478 99288 123484 99340
rect 123536 99328 123542 99340
rect 126974 99328 126980 99340
rect 123536 99300 126980 99328
rect 123536 99288 123542 99300
rect 126974 99288 126980 99300
rect 127032 99288 127038 99340
rect 532234 97996 532240 98048
rect 532292 98036 532298 98048
rect 535454 98036 535460 98048
rect 532292 98008 535460 98036
rect 532292 97996 532298 98008
rect 535454 97996 535460 98008
rect 535512 97996 535518 98048
rect 124858 97928 124864 97980
rect 124916 97968 124922 97980
rect 126974 97968 126980 97980
rect 124916 97940 126980 97968
rect 124916 97928 124922 97940
rect 126974 97928 126980 97940
rect 127032 97928 127038 97980
rect 532142 96636 532148 96688
rect 532200 96676 532206 96688
rect 535454 96676 535460 96688
rect 532200 96648 535460 96676
rect 532200 96636 532206 96648
rect 535454 96636 535460 96648
rect 535512 96636 535518 96688
rect 119338 96568 119344 96620
rect 119396 96608 119402 96620
rect 126974 96608 126980 96620
rect 119396 96580 126980 96608
rect 119396 96568 119402 96580
rect 126974 96568 126980 96580
rect 127032 96568 127038 96620
rect 532050 95208 532056 95260
rect 532108 95248 532114 95260
rect 535454 95248 535460 95260
rect 532108 95220 535460 95248
rect 532108 95208 532114 95220
rect 535454 95208 535460 95220
rect 535512 95208 535518 95260
rect 532510 94188 532516 94240
rect 532568 94228 532574 94240
rect 535454 94228 535460 94240
rect 532568 94200 535460 94228
rect 532568 94188 532574 94200
rect 535454 94188 535460 94200
rect 535512 94188 535518 94240
rect 532418 92488 532424 92540
rect 532476 92528 532482 92540
rect 535454 92528 535460 92540
rect 532476 92500 535460 92528
rect 532476 92488 532482 92500
rect 535454 92488 535460 92500
rect 535512 92488 535518 92540
rect 531958 91060 531964 91112
rect 532016 91100 532022 91112
rect 535454 91100 535460 91112
rect 532016 91072 535460 91100
rect 532016 91060 532022 91072
rect 535454 91060 535460 91072
rect 535512 91060 535518 91112
rect 532602 89700 532608 89752
rect 532660 89740 532666 89752
rect 535454 89740 535460 89752
rect 532660 89712 535460 89740
rect 532660 89700 532666 89712
rect 535454 89700 535460 89712
rect 535512 89700 535518 89752
rect 120718 89632 120724 89684
rect 120776 89672 120782 89684
rect 126974 89672 126980 89684
rect 120776 89644 126980 89672
rect 120776 89632 120782 89644
rect 126974 89632 126980 89644
rect 127032 89632 127038 89684
rect 115934 88544 115940 88596
rect 115992 88584 115998 88596
rect 117958 88584 117964 88596
rect 115992 88556 117964 88584
rect 115992 88544 115998 88556
rect 117958 88544 117964 88556
rect 118016 88544 118022 88596
rect 532050 88340 532056 88392
rect 532108 88380 532114 88392
rect 535454 88380 535460 88392
rect 532108 88352 535460 88380
rect 532108 88340 532114 88352
rect 535454 88340 535460 88352
rect 535512 88340 535518 88392
rect 116578 88272 116584 88324
rect 116636 88312 116642 88324
rect 126974 88312 126980 88324
rect 116636 88284 126980 88312
rect 116636 88272 116642 88284
rect 126974 88272 126980 88284
rect 127032 88272 127038 88324
rect 532326 86980 532332 87032
rect 532384 87020 532390 87032
rect 535454 87020 535460 87032
rect 532384 86992 535460 87020
rect 532384 86980 532390 86992
rect 535454 86980 535460 86992
rect 535512 86980 535518 87032
rect 116670 86912 116676 86964
rect 116728 86952 116734 86964
rect 126974 86952 126980 86964
rect 116728 86924 126980 86952
rect 116728 86912 116734 86924
rect 126974 86912 126980 86924
rect 127032 86912 127038 86964
rect 532510 85552 532516 85604
rect 532568 85592 532574 85604
rect 535454 85592 535460 85604
rect 532568 85564 535460 85592
rect 532568 85552 532574 85564
rect 535454 85552 535460 85564
rect 535512 85552 535518 85604
rect 532602 84192 532608 84244
rect 532660 84232 532666 84244
rect 535454 84232 535460 84244
rect 532660 84204 535460 84232
rect 532660 84192 532666 84204
rect 535454 84192 535460 84204
rect 535512 84192 535518 84244
rect 116762 84124 116768 84176
rect 116820 84164 116826 84176
rect 126974 84164 126980 84176
rect 116820 84136 126980 84164
rect 116820 84124 116826 84136
rect 126974 84124 126980 84136
rect 127032 84124 127038 84176
rect 122098 82764 122104 82816
rect 122156 82804 122162 82816
rect 126974 82804 126980 82816
rect 122156 82776 126980 82804
rect 122156 82764 122162 82776
rect 126974 82764 126980 82776
rect 127032 82764 127038 82816
rect 117958 79976 117964 80028
rect 118016 80016 118022 80028
rect 126974 80016 126980 80028
rect 118016 79988 126980 80016
rect 118016 79976 118022 79988
rect 126974 79976 126980 79988
rect 127032 79976 127038 80028
rect 532142 78684 532148 78736
rect 532200 78724 532206 78736
rect 535638 78724 535644 78736
rect 532200 78696 535644 78724
rect 532200 78684 532206 78696
rect 535638 78684 535644 78696
rect 535696 78684 535702 78736
rect 116118 77936 116124 77988
rect 116176 77976 116182 77988
rect 126974 77976 126980 77988
rect 116176 77948 126980 77976
rect 116176 77936 116182 77948
rect 126974 77936 126980 77948
rect 127032 77936 127038 77988
rect 532602 77188 532608 77240
rect 532660 77228 532666 77240
rect 535546 77228 535552 77240
rect 532660 77200 535552 77228
rect 532660 77188 532666 77200
rect 535546 77188 535552 77200
rect 535604 77188 535610 77240
rect 116578 75896 116584 75948
rect 116636 75936 116642 75948
rect 126974 75936 126980 75948
rect 116636 75908 126980 75936
rect 116636 75896 116642 75908
rect 126974 75896 126980 75908
rect 127032 75896 127038 75948
rect 532602 75828 532608 75880
rect 532660 75868 532666 75880
rect 535454 75868 535460 75880
rect 532660 75840 535460 75868
rect 532660 75828 532666 75840
rect 535454 75828 535460 75840
rect 535512 75828 535518 75880
rect 532602 74468 532608 74520
rect 532660 74508 532666 74520
rect 536282 74508 536288 74520
rect 532660 74480 536288 74508
rect 532660 74468 532666 74480
rect 536282 74468 536288 74480
rect 536340 74468 536346 74520
rect 116762 73176 116768 73228
rect 116820 73216 116826 73228
rect 126974 73216 126980 73228
rect 116820 73188 126980 73216
rect 116820 73176 116826 73188
rect 126974 73176 126980 73188
rect 127032 73176 127038 73228
rect 532418 73108 532424 73160
rect 532476 73148 532482 73160
rect 535546 73148 535552 73160
rect 532476 73120 535552 73148
rect 532476 73108 532482 73120
rect 535546 73108 535552 73120
rect 535604 73108 535610 73160
rect 116670 71748 116676 71800
rect 116728 71788 116734 71800
rect 126974 71788 126980 71800
rect 116728 71760 126980 71788
rect 116728 71748 116734 71760
rect 126974 71748 126980 71760
rect 127032 71748 127038 71800
rect 532418 71680 532424 71732
rect 532476 71720 532482 71732
rect 535638 71720 535644 71732
rect 532476 71692 535644 71720
rect 532476 71680 532482 71692
rect 535638 71680 535644 71692
rect 535696 71680 535702 71732
rect 531774 70524 531780 70576
rect 531832 70564 531838 70576
rect 535730 70564 535736 70576
rect 531832 70536 535736 70564
rect 531832 70524 531838 70536
rect 535730 70524 535736 70536
rect 535788 70524 535794 70576
rect 531958 69776 531964 69828
rect 532016 69816 532022 69828
rect 535546 69816 535552 69828
rect 532016 69788 535552 69816
rect 532016 69776 532022 69788
rect 535546 69776 535552 69788
rect 535604 69776 535610 69828
rect 120810 69028 120816 69080
rect 120868 69068 120874 69080
rect 126974 69068 126980 69080
rect 120868 69040 126980 69068
rect 120868 69028 120874 69040
rect 126974 69028 126980 69040
rect 127032 69028 127038 69080
rect 531958 68144 531964 68196
rect 532016 68184 532022 68196
rect 535454 68184 535460 68196
rect 532016 68156 535460 68184
rect 532016 68144 532022 68156
rect 535454 68144 535460 68156
rect 535512 68144 535518 68196
rect 118050 67600 118056 67652
rect 118108 67640 118114 67652
rect 126974 67640 126980 67652
rect 118108 67612 126980 67640
rect 118108 67600 118114 67612
rect 126974 67600 126980 67612
rect 127032 67600 127038 67652
rect 531958 67532 531964 67584
rect 532016 67572 532022 67584
rect 535546 67572 535552 67584
rect 532016 67544 535552 67572
rect 532016 67532 532022 67544
rect 535546 67532 535552 67544
rect 535604 67532 535610 67584
rect 124858 66240 124864 66292
rect 124916 66280 124922 66292
rect 127434 66280 127440 66292
rect 124916 66252 127440 66280
rect 124916 66240 124922 66252
rect 127434 66240 127440 66252
rect 127492 66240 127498 66292
rect 535454 66280 535460 66292
rect 532712 66252 535460 66280
rect 532142 66172 532148 66224
rect 532200 66212 532206 66224
rect 532712 66212 532740 66252
rect 535454 66240 535460 66252
rect 535512 66240 535518 66292
rect 532200 66184 532740 66212
rect 532200 66172 532206 66184
rect 535454 64920 535460 64932
rect 532712 64892 535460 64920
rect 531314 64812 531320 64864
rect 531372 64852 531378 64864
rect 532712 64852 532740 64892
rect 535454 64880 535460 64892
rect 535512 64880 535518 64932
rect 531372 64824 532740 64852
rect 531372 64812 531378 64824
rect 119338 63520 119344 63572
rect 119396 63560 119402 63572
rect 126974 63560 126980 63572
rect 119396 63532 126980 63560
rect 119396 63520 119402 63532
rect 126974 63520 126980 63532
rect 127032 63520 127038 63572
rect 535454 63560 535460 63572
rect 532712 63532 535460 63560
rect 532142 63452 532148 63504
rect 532200 63492 532206 63504
rect 532712 63492 532740 63532
rect 535454 63520 535460 63532
rect 535512 63520 535518 63572
rect 532200 63464 532740 63492
rect 532200 63452 532206 63464
rect 115198 62092 115204 62144
rect 115256 62132 115262 62144
rect 126974 62132 126980 62144
rect 115256 62104 126980 62132
rect 115256 62092 115262 62104
rect 126974 62092 126980 62104
rect 127032 62092 127038 62144
rect 535454 62132 535460 62144
rect 532712 62104 535460 62132
rect 532326 62024 532332 62076
rect 532384 62064 532390 62076
rect 532712 62064 532740 62104
rect 535454 62092 535460 62104
rect 535512 62092 535518 62144
rect 532384 62036 532740 62064
rect 532384 62024 532390 62036
rect 535454 60772 535460 60784
rect 533724 60744 535460 60772
rect 532510 60664 532516 60716
rect 532568 60704 532574 60716
rect 533724 60704 533752 60744
rect 535454 60732 535460 60744
rect 535512 60732 535518 60784
rect 532568 60676 533752 60704
rect 532568 60664 532574 60676
rect 535454 59412 535460 59424
rect 532712 59384 535460 59412
rect 532602 59304 532608 59356
rect 532660 59344 532666 59356
rect 532712 59344 532740 59384
rect 535454 59372 535460 59384
rect 535512 59372 535518 59424
rect 532660 59316 532740 59344
rect 532660 59304 532666 59316
rect 535454 57984 535460 57996
rect 532712 57956 535460 57984
rect 532418 57876 532424 57928
rect 532476 57916 532482 57928
rect 532712 57916 532740 57956
rect 535454 57944 535460 57956
rect 535512 57944 535518 57996
rect 532476 57888 532740 57916
rect 532476 57876 532482 57888
rect 115290 57196 115296 57248
rect 115348 57236 115354 57248
rect 126974 57236 126980 57248
rect 115348 57208 126980 57236
rect 115348 57196 115354 57208
rect 126974 57196 126980 57208
rect 127032 57196 127038 57248
rect 535454 56624 535460 56636
rect 532712 56596 535460 56624
rect 532602 56516 532608 56568
rect 532660 56556 532666 56568
rect 532712 56556 532740 56596
rect 535454 56584 535460 56596
rect 535512 56584 535518 56636
rect 532660 56528 532740 56556
rect 532660 56516 532666 56528
rect 535454 55264 535460 55276
rect 532712 55236 535460 55264
rect 531314 55156 531320 55208
rect 531372 55196 531378 55208
rect 532712 55196 532740 55236
rect 535454 55224 535460 55236
rect 535512 55224 535518 55276
rect 531372 55168 532740 55196
rect 531372 55156 531378 55168
rect 116578 53796 116584 53848
rect 116636 53836 116642 53848
rect 126974 53836 126980 53848
rect 116636 53808 126980 53836
rect 116636 53796 116642 53808
rect 126974 53796 126980 53808
rect 127032 53796 127038 53848
rect 117958 53048 117964 53100
rect 118016 53088 118022 53100
rect 127802 53088 127808 53100
rect 118016 53060 127808 53088
rect 118016 53048 118022 53060
rect 127802 53048 127808 53060
rect 127860 53048 127866 53100
rect 532142 52980 532148 53032
rect 532200 53020 532206 53032
rect 535454 53020 535460 53032
rect 532200 52992 535460 53020
rect 532200 52980 532206 52992
rect 535454 52980 535460 52992
rect 535512 52980 535518 53032
rect 532602 51280 532608 51332
rect 532660 51320 532666 51332
rect 535454 51320 535460 51332
rect 532660 51292 535460 51320
rect 532660 51280 532666 51292
rect 535454 51280 535460 51292
rect 535512 51280 535518 51332
rect 120718 51076 120724 51128
rect 120776 51116 120782 51128
rect 126974 51116 126980 51128
rect 120776 51088 126980 51116
rect 120776 51076 120782 51088
rect 126974 51076 126980 51088
rect 127032 51076 127038 51128
rect 532510 49988 532516 50040
rect 532568 50028 532574 50040
rect 535454 50028 535460 50040
rect 532568 50000 535460 50028
rect 532568 49988 532574 50000
rect 535454 49988 535460 50000
rect 535512 49988 535518 50040
rect 531958 48628 531964 48680
rect 532016 48668 532022 48680
rect 535454 48668 535460 48680
rect 532016 48640 535460 48668
rect 532016 48628 532022 48640
rect 535454 48628 535460 48640
rect 535512 48628 535518 48680
rect 532602 47404 532608 47456
rect 532660 47444 532666 47456
rect 535454 47444 535460 47456
rect 532660 47416 535460 47444
rect 532660 47404 532666 47416
rect 535454 47404 535460 47416
rect 535512 47404 535518 47456
rect 123478 46928 123484 46980
rect 123536 46968 123542 46980
rect 126974 46968 126980 46980
rect 123536 46940 126980 46968
rect 123536 46928 123542 46940
rect 126974 46928 126980 46940
rect 127032 46928 127038 46980
rect 532602 45772 532608 45824
rect 532660 45812 532666 45824
rect 535454 45812 535460 45824
rect 532660 45784 535460 45812
rect 532660 45772 532666 45784
rect 535454 45772 535460 45784
rect 535512 45772 535518 45824
rect 532510 44548 532516 44600
rect 532568 44588 532574 44600
rect 535454 44588 535460 44600
rect 532568 44560 535460 44588
rect 532568 44548 532574 44560
rect 535454 44548 535460 44560
rect 535512 44548 535518 44600
rect 122098 44140 122104 44192
rect 122156 44180 122162 44192
rect 126974 44180 126980 44192
rect 122156 44152 126980 44180
rect 122156 44140 122162 44152
rect 126974 44140 126980 44152
rect 127032 44140 127038 44192
rect 532602 43052 532608 43104
rect 532660 43092 532666 43104
rect 535454 43092 535460 43104
rect 532660 43064 535460 43092
rect 532660 43052 532666 43064
rect 535454 43052 535460 43064
rect 535512 43052 535518 43104
rect 119430 42780 119436 42832
rect 119488 42820 119494 42832
rect 126974 42820 126980 42832
rect 119488 42792 126980 42820
rect 119488 42780 119494 42792
rect 126974 42780 126980 42792
rect 127032 42780 127038 42832
rect 532602 41692 532608 41744
rect 532660 41732 532666 41744
rect 535454 41732 535460 41744
rect 532660 41704 535460 41732
rect 532660 41692 532666 41704
rect 535454 41692 535460 41704
rect 535512 41692 535518 41744
rect 124950 41420 124956 41472
rect 125008 41460 125014 41472
rect 126974 41460 126980 41472
rect 125008 41432 126980 41460
rect 125008 41420 125014 41432
rect 126974 41420 126980 41432
rect 127032 41420 127038 41472
rect 532602 40128 532608 40180
rect 532660 40168 532666 40180
rect 535454 40168 535460 40180
rect 532660 40140 535460 40168
rect 532660 40128 532666 40140
rect 535454 40128 535460 40140
rect 535512 40128 535518 40180
rect 532602 38768 532608 38820
rect 532660 38808 532666 38820
rect 535454 38808 535460 38820
rect 532660 38780 535460 38808
rect 532660 38768 532666 38780
rect 535454 38768 535460 38780
rect 535512 38768 535518 38820
rect 118142 38632 118148 38684
rect 118200 38672 118206 38684
rect 126974 38672 126980 38684
rect 118200 38644 126980 38672
rect 118200 38632 118206 38644
rect 126974 38632 126980 38644
rect 127032 38632 127038 38684
rect 532602 37408 532608 37460
rect 532660 37448 532666 37460
rect 535362 37448 535368 37460
rect 532660 37420 535368 37448
rect 532660 37408 532666 37420
rect 535362 37408 535368 37420
rect 535420 37408 535426 37460
rect 116670 37272 116676 37324
rect 116728 37312 116734 37324
rect 126974 37312 126980 37324
rect 116728 37284 126980 37312
rect 116728 37272 116734 37284
rect 126974 37272 126980 37284
rect 127032 37272 127038 37324
rect 532326 36048 532332 36100
rect 532384 36088 532390 36100
rect 535362 36088 535368 36100
rect 532384 36060 535368 36088
rect 532384 36048 532390 36060
rect 535362 36048 535368 36060
rect 535420 36048 535426 36100
rect 532602 34688 532608 34740
rect 532660 34728 532666 34740
rect 535362 34728 535368 34740
rect 532660 34700 535368 34728
rect 532660 34688 532666 34700
rect 535362 34688 535368 34700
rect 535420 34688 535426 34740
rect 116854 33328 116860 33380
rect 116912 33368 116918 33380
rect 120810 33368 120816 33380
rect 116912 33340 120816 33368
rect 116912 33328 116918 33340
rect 120810 33328 120816 33340
rect 120868 33328 120874 33380
rect 531958 33328 531964 33380
rect 532016 33368 532022 33380
rect 535362 33368 535368 33380
rect 532016 33340 535368 33368
rect 532016 33328 532022 33340
rect 535362 33328 535368 33340
rect 535420 33328 535426 33380
rect 123570 33124 123576 33176
rect 123628 33164 123634 33176
rect 126974 33164 126980 33176
rect 123628 33136 126980 33164
rect 123628 33124 123634 33136
rect 126974 33124 126980 33136
rect 127032 33124 127038 33176
rect 532602 31968 532608 32020
rect 532660 32008 532666 32020
rect 535362 32008 535368 32020
rect 532660 31980 535368 32008
rect 532660 31968 532666 31980
rect 535362 31968 535368 31980
rect 535420 31968 535426 32020
rect 122190 31764 122196 31816
rect 122248 31804 122254 31816
rect 126974 31804 126980 31816
rect 122248 31776 126980 31804
rect 122248 31764 122254 31776
rect 126974 31764 126980 31776
rect 127032 31764 127038 31816
rect 532602 30608 532608 30660
rect 532660 30648 532666 30660
rect 535362 30648 535368 30660
rect 532660 30620 535368 30648
rect 532660 30608 532666 30620
rect 535362 30608 535368 30620
rect 535420 30608 535426 30660
rect 532602 29248 532608 29300
rect 532660 29288 532666 29300
rect 535362 29288 535368 29300
rect 532660 29260 535368 29288
rect 532660 29248 532666 29260
rect 535362 29248 535368 29260
rect 535420 29248 535426 29300
rect 120810 28976 120816 29028
rect 120868 29016 120874 29028
rect 126974 29016 126980 29028
rect 120868 28988 126980 29016
rect 120868 28976 120874 28988
rect 126974 28976 126980 28988
rect 127032 28976 127038 29028
rect 119522 27616 119528 27668
rect 119580 27656 119586 27668
rect 126974 27656 126980 27668
rect 119580 27628 126980 27656
rect 119580 27616 119586 27628
rect 126974 27616 126980 27628
rect 127032 27616 127038 27668
rect 532602 27616 532608 27668
rect 532660 27656 532666 27668
rect 532660 27628 534120 27656
rect 532660 27616 532666 27628
rect 534092 27588 534120 27628
rect 535454 27588 535460 27600
rect 534092 27560 535460 27588
rect 535454 27548 535460 27560
rect 535512 27548 535518 27600
rect 532326 26528 532332 26580
rect 532384 26568 532390 26580
rect 535362 26568 535368 26580
rect 532384 26540 535368 26568
rect 532384 26528 532390 26540
rect 535362 26528 535368 26540
rect 535420 26528 535426 26580
rect 116762 24828 116768 24880
rect 116820 24868 116826 24880
rect 126974 24868 126980 24880
rect 116820 24840 126980 24868
rect 116820 24828 116826 24840
rect 126974 24828 126980 24840
rect 127032 24828 127038 24880
rect 532602 24828 532608 24880
rect 532660 24868 532666 24880
rect 535362 24868 535368 24880
rect 532660 24840 535368 24868
rect 532660 24828 532666 24840
rect 535362 24828 535368 24840
rect 535420 24828 535426 24880
rect 532050 23672 532056 23724
rect 532108 23712 532114 23724
rect 535270 23712 535276 23724
rect 532108 23684 535276 23712
rect 532108 23672 532114 23684
rect 535270 23672 535276 23684
rect 535328 23672 535334 23724
rect 531958 22312 531964 22364
rect 532016 22352 532022 22364
rect 535362 22352 535368 22364
rect 532016 22324 535368 22352
rect 532016 22312 532022 22324
rect 535362 22312 535368 22324
rect 535420 22312 535426 22364
rect 123662 22108 123668 22160
rect 123720 22148 123726 22160
rect 126974 22148 126980 22160
rect 123720 22120 126980 22148
rect 123720 22108 123726 22120
rect 126974 22108 126980 22120
rect 127032 22108 127038 22160
rect 115934 21088 115940 21140
rect 115992 21128 115998 21140
rect 118050 21128 118056 21140
rect 115992 21100 118056 21128
rect 115992 21088 115998 21100
rect 118050 21088 118056 21100
rect 118108 21088 118114 21140
rect 531958 20952 531964 21004
rect 532016 20992 532022 21004
rect 535270 20992 535276 21004
rect 532016 20964 535276 20992
rect 532016 20952 532022 20964
rect 535270 20952 535276 20964
rect 535328 20952 535334 21004
rect 531958 19592 531964 19644
rect 532016 19632 532022 19644
rect 535178 19632 535184 19644
rect 532016 19604 535184 19632
rect 532016 19592 532022 19604
rect 535178 19592 535184 19604
rect 535236 19592 535242 19644
rect 122282 19320 122288 19372
rect 122340 19360 122346 19372
rect 126974 19360 126980 19372
rect 122340 19332 126980 19360
rect 122340 19320 122346 19332
rect 126974 19320 126980 19332
rect 127032 19320 127038 19372
rect 120902 17960 120908 18012
rect 120960 18000 120966 18012
rect 126974 18000 126980 18012
rect 120960 17972 126980 18000
rect 120960 17960 120966 17972
rect 126974 17960 126980 17972
rect 127032 17960 127038 18012
rect 532326 17960 532332 18012
rect 532384 18000 532390 18012
rect 535362 18000 535368 18012
rect 532384 17972 535368 18000
rect 532384 17960 532390 17972
rect 535362 17960 535368 17972
rect 535420 17960 535426 18012
rect 532234 16872 532240 16924
rect 532292 16912 532298 16924
rect 535270 16912 535276 16924
rect 532292 16884 535276 16912
rect 532292 16872 532298 16884
rect 535270 16872 535276 16884
rect 535328 16872 535334 16924
rect 532602 15512 532608 15564
rect 532660 15552 532666 15564
rect 535362 15552 535368 15564
rect 532660 15524 535368 15552
rect 532660 15512 532666 15524
rect 535362 15512 535368 15524
rect 535420 15512 535426 15564
rect 532142 14152 532148 14204
rect 532200 14192 532206 14204
rect 535270 14192 535276 14204
rect 532200 14164 535276 14192
rect 532200 14152 532206 14164
rect 535270 14152 535276 14164
rect 535328 14152 535334 14204
rect 118050 13812 118056 13864
rect 118108 13852 118114 13864
rect 126974 13852 126980 13864
rect 118108 13824 126980 13852
rect 118108 13812 118114 13824
rect 126974 13812 126980 13824
rect 127032 13812 127038 13864
rect 531590 12656 531596 12708
rect 531648 12696 531654 12708
rect 535362 12696 535368 12708
rect 531648 12668 535368 12696
rect 531648 12656 531654 12668
rect 535362 12656 535368 12668
rect 535420 12656 535426 12708
rect 115382 12452 115388 12504
rect 115440 12492 115446 12504
rect 126974 12492 126980 12504
rect 115440 12464 126980 12492
rect 115440 12452 115446 12464
rect 126974 12452 126980 12464
rect 127032 12452 127038 12504
rect 531958 11296 531964 11348
rect 532016 11336 532022 11348
rect 535178 11336 535184 11348
rect 532016 11308 535184 11336
rect 532016 11296 532022 11308
rect 535178 11296 535184 11308
rect 535236 11296 535242 11348
rect 125042 10888 125048 10940
rect 125100 10928 125106 10940
rect 127710 10928 127716 10940
rect 125100 10900 127716 10928
rect 125100 10888 125106 10900
rect 127710 10888 127716 10900
rect 127768 10888 127774 10940
rect 531774 9664 531780 9716
rect 531832 9704 531838 9716
rect 534994 9704 535000 9716
rect 531832 9676 535000 9704
rect 531832 9664 531838 9676
rect 534994 9664 535000 9676
rect 535052 9664 535058 9716
rect 117222 9052 117228 9104
rect 117280 9092 117286 9104
rect 124858 9092 124864 9104
rect 117280 9064 124864 9092
rect 117280 9052 117286 9064
rect 124858 9052 124864 9064
rect 124916 9052 124922 9104
rect 124306 8984 124312 9036
rect 124364 9024 124370 9036
rect 127250 9024 127256 9036
rect 124364 8996 127256 9024
rect 124364 8984 124370 8996
rect 127250 8984 127256 8996
rect 127308 8984 127314 9036
rect 532234 8304 532240 8356
rect 532292 8344 532298 8356
rect 535270 8344 535276 8356
rect 532292 8316 535276 8344
rect 532292 8304 532298 8316
rect 535270 8304 535276 8316
rect 535328 8304 535334 8356
rect 531958 7080 531964 7132
rect 532016 7120 532022 7132
rect 535178 7120 535184 7132
rect 532016 7092 535184 7120
rect 532016 7080 532022 7092
rect 535178 7080 535184 7092
rect 535236 7080 535242 7132
rect 531590 5856 531596 5908
rect 531648 5896 531654 5908
rect 535362 5896 535368 5908
rect 531648 5868 535368 5896
rect 531648 5856 531654 5868
rect 535362 5856 535368 5868
rect 535420 5856 535426 5908
rect 124858 5516 124864 5568
rect 124916 5556 124922 5568
rect 126974 5556 126980 5568
rect 124916 5528 126980 5556
rect 124916 5516 124922 5528
rect 126974 5516 126980 5528
rect 127032 5516 127038 5568
rect 95973 5355 96031 5361
rect 95973 5321 95985 5355
rect 96019 5352 96031 5355
rect 116578 5352 116584 5364
rect 96019 5324 116584 5352
rect 96019 5321 96031 5324
rect 95973 5315 96031 5321
rect 116578 5312 116584 5324
rect 116636 5312 116642 5364
rect 82633 5287 82691 5293
rect 82633 5253 82645 5287
rect 82679 5284 82691 5287
rect 123478 5284 123484 5296
rect 82679 5256 123484 5284
rect 82679 5253 82691 5256
rect 82633 5247 82691 5253
rect 123478 5244 123484 5256
rect 123536 5244 123542 5296
rect 79321 5219 79379 5225
rect 79321 5185 79333 5219
rect 79367 5216 79379 5219
rect 122098 5216 122104 5228
rect 79367 5188 122104 5216
rect 79367 5185 79379 5188
rect 79321 5179 79379 5185
rect 122098 5176 122104 5188
rect 122156 5176 122162 5228
rect 75825 5151 75883 5157
rect 75825 5117 75837 5151
rect 75871 5148 75883 5151
rect 119430 5148 119436 5160
rect 75871 5120 119436 5148
rect 75871 5117 75883 5120
rect 75825 5111 75883 5117
rect 119430 5108 119436 5120
rect 119488 5108 119494 5160
rect 65981 5083 66039 5089
rect 65981 5049 65993 5083
rect 66027 5080 66039 5083
rect 116670 5080 116676 5092
rect 66027 5052 116676 5080
rect 66027 5049 66039 5052
rect 65981 5043 66039 5049
rect 116670 5040 116676 5052
rect 116728 5040 116734 5092
rect 62669 5015 62727 5021
rect 62669 4981 62681 5015
rect 62715 5012 62727 5015
rect 126330 5012 126336 5024
rect 62715 4984 126336 5012
rect 62715 4981 62727 4984
rect 62669 4975 62727 4981
rect 126330 4972 126336 4984
rect 126388 4972 126394 5024
rect 55953 4947 56011 4953
rect 55953 4913 55965 4947
rect 55999 4944 56011 4947
rect 123570 4944 123576 4956
rect 55999 4916 123576 4944
rect 55999 4913 56011 4916
rect 55953 4907 56011 4913
rect 123570 4904 123576 4916
rect 123628 4904 123634 4956
rect 52641 4879 52699 4885
rect 52641 4845 52653 4879
rect 52687 4876 52699 4879
rect 120810 4876 120816 4888
rect 52687 4848 120816 4876
rect 52687 4845 52699 4848
rect 52641 4839 52699 4845
rect 120810 4836 120816 4848
rect 120868 4836 120874 4888
rect 124858 4808 124864 4820
rect 16546 4780 48314 4808
rect 9306 4632 9312 4684
rect 9364 4672 9370 4684
rect 16546 4672 16574 4780
rect 48286 4740 48314 4780
rect 57946 4780 124864 4808
rect 57946 4740 57974 4780
rect 124858 4768 124864 4780
rect 124916 4768 124922 4820
rect 48286 4712 57974 4740
rect 9364 4644 16574 4672
rect 9364 4632 9370 4644
rect 49326 4632 49332 4684
rect 49384 4672 49390 4684
rect 52641 4675 52699 4681
rect 52641 4672 52653 4675
rect 49384 4644 52653 4672
rect 49384 4632 49390 4644
rect 52641 4641 52653 4644
rect 52687 4641 52699 4675
rect 55950 4672 55956 4684
rect 55911 4644 55956 4672
rect 52641 4635 52699 4641
rect 55950 4632 55956 4644
rect 56008 4632 56014 4684
rect 62666 4672 62672 4684
rect 62627 4644 62672 4672
rect 62666 4632 62672 4644
rect 62724 4632 62730 4684
rect 65978 4672 65984 4684
rect 65939 4644 65984 4672
rect 65978 4632 65984 4644
rect 66036 4632 66042 4684
rect 75822 4672 75828 4684
rect 75783 4644 75828 4672
rect 75822 4632 75828 4644
rect 75880 4632 75886 4684
rect 79318 4672 79324 4684
rect 79279 4644 79324 4672
rect 79318 4632 79324 4644
rect 79376 4632 79382 4684
rect 82630 4672 82636 4684
rect 82591 4644 82636 4672
rect 82630 4632 82636 4644
rect 82688 4632 82694 4684
rect 95970 4672 95976 4684
rect 95931 4644 95976 4672
rect 95970 4632 95976 4644
rect 96028 4632 96034 4684
rect 532602 4496 532608 4548
rect 532660 4536 532666 4548
rect 535454 4536 535460 4548
rect 532660 4508 535460 4536
rect 532660 4496 532666 4508
rect 535454 4496 535460 4508
rect 535512 4496 535518 4548
rect 117222 4156 117228 4208
rect 117280 4196 117286 4208
rect 126974 4196 126980 4208
rect 117280 4168 126980 4196
rect 117280 4156 117286 4168
rect 126974 4156 126980 4168
rect 127032 4156 127038 4208
rect 5994 3544 6000 3596
rect 6052 3584 6058 3596
rect 117222 3584 117228 3596
rect 6052 3556 117228 3584
rect 6052 3544 6058 3556
rect 117222 3544 117228 3556
rect 117280 3544 117286 3596
rect 105630 3476 105636 3528
rect 105688 3516 105694 3528
rect 127618 3516 127624 3528
rect 105688 3488 127624 3516
rect 105688 3476 105694 3488
rect 127618 3476 127624 3488
rect 127676 3476 127682 3528
rect 91094 3408 91100 3460
rect 91152 3448 91158 3460
rect 127802 3448 127808 3460
rect 91152 3420 127808 3448
rect 91152 3408 91158 3420
rect 127802 3408 127808 3420
rect 127860 3408 127866 3460
rect 33686 3340 33692 3392
rect 33744 3380 33750 3392
rect 128354 3380 128360 3392
rect 33744 3352 128360 3380
rect 33744 3340 33750 3352
rect 128354 3340 128360 3352
rect 128412 3340 128418 3392
rect 89346 3272 89352 3324
rect 89404 3312 89410 3324
rect 120718 3312 120724 3324
rect 89404 3284 120724 3312
rect 89404 3272 89410 3284
rect 120718 3272 120724 3284
rect 120776 3272 120782 3324
rect 68922 3204 68928 3256
rect 68980 3244 68986 3256
rect 118142 3244 118148 3256
rect 68980 3216 118148 3244
rect 68980 3204 68986 3216
rect 118142 3204 118148 3216
rect 118200 3204 118206 3256
rect 52362 3136 52368 3188
rect 52420 3176 52426 3188
rect 122190 3176 122196 3188
rect 52420 3148 122196 3176
rect 52420 3136 52426 3148
rect 122190 3136 122196 3148
rect 122248 3136 122254 3188
rect 45922 3068 45928 3120
rect 45980 3108 45986 3120
rect 119522 3108 119528 3120
rect 45980 3080 119528 3108
rect 45980 3068 45986 3080
rect 119522 3068 119528 3080
rect 119580 3068 119586 3120
rect 42610 3000 42616 3052
rect 42668 3040 42674 3052
rect 116762 3040 116768 3052
rect 42668 3012 116768 3040
rect 42668 3000 42674 3012
rect 116762 3000 116768 3012
rect 116820 3000 116826 3052
rect 39298 2932 39304 2984
rect 39356 2972 39362 2984
rect 126422 2972 126428 2984
rect 39356 2944 126428 2972
rect 39356 2932 39362 2944
rect 126422 2932 126428 2944
rect 126480 2932 126486 2984
rect 101122 2864 101128 2916
rect 101180 2904 101186 2916
rect 101180 2876 129780 2904
rect 101180 2864 101186 2876
rect 15930 2796 15936 2848
rect 15988 2836 15994 2848
rect 127710 2836 127716 2848
rect 15988 2808 127716 2836
rect 15988 2796 15994 2808
rect 127710 2796 127716 2808
rect 127768 2796 127774 2848
rect 12342 2728 12348 2780
rect 12400 2768 12406 2780
rect 91094 2768 91100 2780
rect 12400 2740 91100 2768
rect 12400 2728 12406 2740
rect 91094 2728 91100 2740
rect 91152 2728 91158 2780
rect 99282 2728 99288 2780
rect 99340 2768 99346 2780
rect 105630 2768 105636 2780
rect 99340 2740 105636 2768
rect 99340 2728 99346 2740
rect 105630 2728 105636 2740
rect 105688 2728 105694 2780
rect 117958 2768 117964 2780
rect 108316 2740 117964 2768
rect 102686 2660 102692 2712
rect 102744 2700 102750 2712
rect 108316 2700 108344 2740
rect 117958 2728 117964 2740
rect 118016 2728 118022 2780
rect 129752 2768 129780 2876
rect 313274 2864 313280 2916
rect 313332 2904 313338 2916
rect 371142 2904 371148 2916
rect 313332 2876 371148 2904
rect 313332 2864 313338 2876
rect 371142 2864 371148 2876
rect 371200 2864 371206 2916
rect 236178 2796 236184 2848
rect 236236 2836 236242 2848
rect 236236 2808 244320 2836
rect 236236 2796 236242 2808
rect 179966 2768 179972 2780
rect 129752 2740 179972 2768
rect 179966 2728 179972 2740
rect 180024 2728 180030 2780
rect 244292 2768 244320 2808
rect 279970 2796 279976 2848
rect 280028 2836 280034 2848
rect 303706 2836 303712 2848
rect 280028 2808 303712 2836
rect 280028 2796 280034 2808
rect 303706 2796 303712 2808
rect 303764 2796 303770 2848
rect 346670 2796 346676 2848
rect 346728 2836 346734 2848
rect 438670 2836 438676 2848
rect 346728 2808 438676 2836
rect 346728 2796 346734 2808
rect 438670 2796 438676 2808
rect 438728 2796 438734 2848
rect 246666 2768 246672 2780
rect 244292 2740 246672 2768
rect 246666 2728 246672 2740
rect 246724 2728 246730 2780
rect 102744 2672 108344 2700
rect 102744 2660 102750 2672
rect 108942 2660 108948 2712
rect 109000 2700 109006 2712
rect 115198 2700 115204 2712
rect 109000 2672 115204 2700
rect 109000 2660 109006 2672
rect 115198 2660 115204 2672
rect 115256 2660 115262 2712
rect 128354 2660 128360 2712
rect 128412 2700 128418 2712
rect 146662 2700 146668 2712
rect 128412 2672 146668 2700
rect 128412 2660 128418 2672
rect 146662 2660 146668 2672
rect 146720 2660 146726 2712
rect 112622 2592 112628 2644
rect 112680 2632 112686 2644
rect 119338 2632 119344 2644
rect 112680 2604 119344 2632
rect 112680 2592 112686 2604
rect 119338 2592 119344 2604
rect 119396 2592 119402 2644
rect 28902 2524 28908 2576
rect 28960 2564 28966 2576
rect 120902 2564 120908 2576
rect 28960 2536 120908 2564
rect 28960 2524 28966 2536
rect 120902 2524 120908 2536
rect 120960 2524 120966 2576
rect 32582 2456 32588 2508
rect 32640 2496 32646 2508
rect 122282 2496 122288 2508
rect 32640 2468 122288 2496
rect 32640 2456 32646 2468
rect 122282 2456 122288 2468
rect 122340 2456 122346 2508
rect 35802 2388 35808 2440
rect 35860 2428 35866 2440
rect 123662 2428 123668 2440
rect 35860 2400 123668 2428
rect 35860 2388 35866 2400
rect 123662 2388 123668 2400
rect 123720 2388 123726 2440
rect 92382 2320 92388 2372
rect 92440 2360 92446 2372
rect 125042 2360 125048 2372
rect 92440 2332 125048 2360
rect 92440 2320 92446 2332
rect 125042 2320 125048 2332
rect 125100 2320 125106 2372
rect 72602 2252 72608 2304
rect 72660 2292 72666 2304
rect 124950 2292 124956 2304
rect 72660 2264 124956 2292
rect 72660 2252 72666 2264
rect 124950 2252 124956 2264
rect 125008 2252 125014 2304
rect 85942 2184 85948 2236
rect 86000 2224 86006 2236
rect 126238 2224 126244 2236
rect 86000 2196 126244 2224
rect 86000 2184 86006 2196
rect 126238 2184 126244 2196
rect 126296 2184 126302 2236
rect 19242 2116 19248 2168
rect 19300 2156 19306 2168
rect 115382 2156 115388 2168
rect 19300 2128 115388 2156
rect 19300 2116 19306 2128
rect 115382 2116 115388 2128
rect 115440 2116 115446 2168
rect 168650 2116 168656 2168
rect 168708 2156 168714 2168
rect 213270 2156 213276 2168
rect 168708 2128 213276 2156
rect 168708 2116 168714 2128
rect 213270 2116 213276 2128
rect 213328 2116 213334 2168
rect 25958 2048 25964 2100
rect 26016 2088 26022 2100
rect 124306 2088 124312 2100
rect 26016 2060 124312 2088
rect 26016 2048 26022 2060
rect 124306 2048 124312 2060
rect 124364 2048 124370 2100
rect 183462 2048 183468 2100
rect 183520 2088 183526 2100
rect 379974 2088 379980 2100
rect 183520 2060 379980 2088
rect 183520 2048 183526 2060
rect 379974 2048 379980 2060
rect 380032 2088 380038 2100
rect 506198 2088 506204 2100
rect 380032 2060 506204 2088
rect 380032 2048 380038 2060
rect 506198 2048 506204 2060
rect 506256 2048 506262 2100
rect 22646 1980 22652 2032
rect 22704 2020 22710 2032
rect 118050 2020 118056 2032
rect 22704 1992 118056 2020
rect 22704 1980 22710 1992
rect 118050 1980 118056 1992
rect 118108 1980 118114 2032
rect 105998 1912 106004 1964
rect 106056 1952 106062 1964
rect 115290 1952 115296 1964
rect 106056 1924 115296 1952
rect 106056 1912 106062 1924
rect 115290 1912 115296 1924
rect 115348 1912 115354 1964
rect 59262 1300 59268 1352
rect 59320 1340 59326 1352
rect 183462 1340 183468 1352
rect 59320 1312 183468 1340
rect 59320 1300 59326 1312
rect 183462 1300 183468 1312
rect 183520 1300 183526 1352
<< via1 >>
rect 60464 163888 60516 163940
rect 63868 163888 63920 163940
rect 174452 163888 174504 163940
rect 177120 163888 177172 163940
rect 56784 163820 56836 163872
rect 171876 163820 171928 163872
rect 53288 163752 53340 163804
rect 169300 163752 169352 163804
rect 49884 163684 49936 163736
rect 165620 163684 165672 163736
rect 42892 163616 42944 163668
rect 161664 163616 161716 163668
rect 46388 163548 46440 163600
rect 164240 163548 164292 163600
rect 35992 163480 36044 163532
rect 156236 163480 156288 163532
rect 39396 163412 39448 163464
rect 159180 163412 159232 163464
rect 167736 163412 167788 163464
rect 254124 163412 254176 163464
rect 114836 163344 114888 163396
rect 214380 163344 214432 163396
rect 112260 163276 112312 163328
rect 212632 163276 212684 163328
rect 110512 163208 110564 163260
rect 211804 163208 211856 163260
rect 98368 163140 98420 163192
rect 202236 163140 202288 163192
rect 87880 163072 87932 163124
rect 195060 163072 195112 163124
rect 84384 163004 84436 163056
rect 192484 163004 192536 163056
rect 88800 162936 88852 162988
rect 194692 162936 194744 162988
rect 80980 162868 81032 162920
rect 189264 162868 189316 162920
rect 77484 162800 77536 162852
rect 186596 162800 186648 162852
rect 79232 162732 79284 162784
rect 188344 162732 188396 162784
rect 73988 162664 74040 162716
rect 183560 162664 183612 162716
rect 70584 162596 70636 162648
rect 182272 162596 182324 162648
rect 184940 162596 184992 162648
rect 267004 162596 267056 162648
rect 165896 162528 165948 162580
rect 252928 162528 252980 162580
rect 67088 162460 67140 162512
rect 179696 162460 179748 162512
rect 58440 162392 58492 162444
rect 172796 162392 172848 162444
rect 174544 162392 174596 162444
rect 258080 162392 258132 162444
rect 160744 162324 160796 162376
rect 249064 162324 249116 162376
rect 164148 162256 164200 162308
rect 251640 162256 251692 162308
rect 149428 162188 149480 162240
rect 240324 162188 240376 162240
rect 153752 162120 153804 162172
rect 243820 162120 243872 162172
rect 141608 162052 141660 162104
rect 234896 162052 234948 162104
rect 139860 161984 139912 162036
rect 233424 161984 233476 162036
rect 124312 161916 124364 161968
rect 221280 161916 221332 161968
rect 126060 161848 126112 161900
rect 223028 161848 223080 161900
rect 31576 161780 31628 161832
rect 153384 161780 153436 161832
rect 182364 161780 182416 161832
rect 265072 161780 265124 161832
rect 28080 161712 28132 161764
rect 150808 161712 150860 161764
rect 178040 161712 178092 161764
rect 261208 161712 261260 161764
rect 24584 161644 24636 161696
rect 148232 161644 148284 161696
rect 161572 161644 161624 161696
rect 248512 161644 248564 161696
rect 21180 161576 21232 161628
rect 145656 161576 145708 161628
rect 158996 161576 159048 161628
rect 247316 161576 247368 161628
rect 17684 161508 17736 161560
rect 142436 161508 142488 161560
rect 157248 161508 157300 161560
rect 246396 161508 246448 161560
rect 14188 161440 14240 161492
rect 140504 161440 140556 161492
rect 146852 161440 146904 161492
rect 238852 161440 238904 161492
rect 243084 161440 243136 161492
rect 309692 161440 309744 161492
rect 163320 161372 163372 161424
rect 250996 161372 251048 161424
rect 253480 161372 253532 161424
rect 317696 161372 317748 161424
rect 121736 161304 121788 161356
rect 220176 161304 220228 161356
rect 225696 161304 225748 161356
rect 297180 161304 297232 161356
rect 105268 161236 105320 161288
rect 207940 161236 207992 161288
rect 211896 161236 211948 161288
rect 286876 161236 286928 161288
rect 90456 161168 90508 161220
rect 196992 161168 197044 161220
rect 199752 161168 199804 161220
rect 277952 161168 278004 161220
rect 80060 161100 80112 161152
rect 189172 161100 189224 161152
rect 191012 161100 191064 161152
rect 271512 161100 271564 161152
rect 66260 161032 66312 161084
rect 179052 161032 179104 161084
rect 180616 161032 180668 161084
rect 263784 161032 263836 161084
rect 265624 161032 265676 161084
rect 326712 161032 326764 161084
rect 37648 160964 37700 161016
rect 157892 160964 157944 161016
rect 166816 160964 166868 161016
rect 253480 160964 253532 161016
rect 255228 160964 255280 161016
rect 318984 160964 319036 161016
rect 26332 160896 26384 160948
rect 149520 160896 149572 160948
rect 159824 160896 159876 160948
rect 248420 160896 248472 160948
rect 249984 160896 250036 160948
rect 315120 160896 315172 160948
rect 18512 160828 18564 160880
rect 143724 160828 143776 160880
rect 152924 160828 152976 160880
rect 243268 160828 243320 160880
rect 246488 160828 246540 160880
rect 312636 160828 312688 160880
rect 11612 160760 11664 160812
rect 138572 160760 138624 160812
rect 145932 160760 145984 160812
rect 4712 160692 4764 160744
rect 133420 160692 133472 160744
rect 139032 160692 139084 160744
rect 232964 160760 233016 160812
rect 239588 160760 239640 160812
rect 307484 160760 307536 160812
rect 232688 160692 232740 160744
rect 302332 160692 302384 160744
rect 170220 160624 170272 160676
rect 255964 160624 256016 160676
rect 256884 160624 256936 160676
rect 320272 160624 320324 160676
rect 173716 160556 173768 160608
rect 258540 160556 258592 160608
rect 263876 160556 263928 160608
rect 325332 160556 325384 160608
rect 238116 160488 238168 160540
rect 100944 160216 100996 160268
rect 165528 160216 165580 160268
rect 50620 160148 50672 160200
rect 167460 160148 167512 160200
rect 28908 160080 28960 160132
rect 151452 160080 151504 160132
rect 138204 160012 138256 160064
rect 232320 160012 232372 160064
rect 259552 160012 259604 160064
rect 311900 160012 311952 160064
rect 338396 160012 338448 160064
rect 376668 160012 376720 160064
rect 418160 160012 418212 160064
rect 439688 160012 439740 160064
rect 452844 160012 452896 160064
rect 463792 160012 463844 160064
rect 484032 160012 484084 160064
rect 486608 160012 486660 160064
rect 488264 160012 488316 160064
rect 61844 159944 61896 159996
rect 118700 159944 118752 159996
rect 131212 159944 131264 159996
rect 225052 159944 225104 159996
rect 245660 159944 245712 159996
rect 301780 159944 301832 159996
rect 331496 159944 331548 159996
rect 372712 159944 372764 159996
rect 408592 159944 408644 159996
rect 432696 159944 432748 159996
rect 445852 159944 445904 159996
rect 456892 159944 456944 159996
rect 458916 159944 458968 159996
rect 469864 159944 469916 159996
rect 475384 159944 475436 159996
rect 481088 159944 481140 159996
rect 488724 159944 488776 159996
rect 41052 159876 41104 159928
rect 56508 159876 56560 159928
rect 89628 159876 89680 159928
rect 186228 159876 186280 159928
rect 196256 159876 196308 159928
rect 260564 159876 260616 159928
rect 266452 159876 266504 159928
rect 316224 159876 316276 159928
rect 339316 159876 339368 159928
rect 381268 159876 381320 159928
rect 394792 159876 394844 159928
rect 420920 159876 420972 159928
rect 451096 159876 451148 159928
rect 462136 159876 462188 159928
rect 468392 159876 468444 159928
rect 33324 159808 33376 159860
rect 49608 159808 49660 159860
rect 71412 159808 71464 159860
rect 114652 159808 114704 159860
rect 119068 159808 119120 159860
rect 218244 159808 218296 159860
rect 235264 159808 235316 159860
rect 291844 159808 291896 159860
rect 321928 159808 321980 159860
rect 366916 159808 366968 159860
rect 376576 159808 376628 159860
rect 391940 159808 391992 159860
rect 393872 159808 393924 159860
rect 421748 159808 421800 159860
rect 432052 159808 432104 159860
rect 436008 159808 436060 159860
rect 450268 159808 450320 159860
rect 462228 159808 462280 159860
rect 470140 159808 470192 159860
rect 471888 159876 471940 159928
rect 476120 159876 476172 159928
rect 477960 159876 478012 159928
rect 484032 159876 484084 159928
rect 473728 159808 473780 159860
rect 19432 159740 19484 159792
rect 41420 159740 41472 159792
rect 47124 159740 47176 159792
rect 100760 159740 100812 159792
rect 113916 159740 113968 159792
rect 214288 159740 214340 159792
rect 238760 159740 238812 159792
rect 296628 159740 296680 159792
rect 324504 159740 324556 159792
rect 370412 159740 370464 159792
rect 380900 159740 380952 159792
rect 411996 159740 412048 159792
rect 425980 159740 426032 159792
rect 445484 159740 445536 159792
rect 451924 159740 451976 159792
rect 462872 159740 462924 159792
rect 465816 159740 465868 159792
rect 471888 159740 471940 159792
rect 478880 159740 478932 159792
rect 484676 159740 484728 159792
rect 32404 159672 32456 159724
rect 69664 159672 69716 159724
rect 82728 159672 82780 159724
rect 183468 159672 183520 159724
rect 185860 159672 185912 159724
rect 264980 159672 265032 159724
rect 273352 159672 273404 159724
rect 328368 159672 328420 159724
rect 328828 159672 328880 159724
rect 373632 159672 373684 159724
rect 379980 159672 380032 159724
rect 411168 159672 411220 159724
rect 412088 159672 412140 159724
rect 435272 159672 435324 159724
rect 448520 159672 448572 159724
rect 459836 159672 459888 159724
rect 475752 159672 475804 159724
rect 22008 159604 22060 159656
rect 62120 159604 62172 159656
rect 101772 159604 101824 159656
rect 205364 159604 205416 159656
rect 221372 159604 221424 159656
rect 280988 159604 281040 159656
rect 308036 159604 308088 159656
rect 356428 159604 356480 159656
rect 367008 159604 367060 159656
rect 397276 159604 397328 159656
rect 401692 159604 401744 159656
rect 427544 159604 427596 159656
rect 431132 159604 431184 159656
rect 437480 159604 437532 159656
rect 442448 159604 442500 159656
rect 445668 159604 445720 159656
rect 447600 159604 447652 159656
rect 458180 159604 458232 159656
rect 460664 159604 460716 159656
rect 471152 159604 471204 159656
rect 5540 159536 5592 159588
rect 28908 159536 28960 159588
rect 34980 159536 35032 159588
rect 80060 159536 80112 159588
rect 100852 159536 100904 159588
rect 204720 159536 204772 159588
rect 213552 159536 213604 159588
rect 224960 159536 225012 159588
rect 228364 159536 228416 159588
rect 289728 159536 289780 159588
rect 301136 159536 301188 159588
rect 350172 159536 350224 159588
rect 353116 159536 353168 159588
rect 385960 159536 386012 159588
rect 386972 159536 387024 159588
rect 415216 159536 415268 159588
rect 421656 159536 421708 159588
rect 442264 159536 442316 159588
rect 449348 159536 449400 159588
rect 1216 159468 1268 159520
rect 89720 159468 89772 159520
rect 91376 159468 91428 159520
rect 99380 159468 99432 159520
rect 104348 159468 104400 159520
rect 207296 159468 207348 159520
rect 210148 159468 210200 159520
rect 276112 159468 276164 159520
rect 294236 159468 294288 159520
rect 347688 159468 347740 159520
rect 360108 159468 360160 159520
rect 396724 159468 396776 159520
rect 400864 159468 400916 159520
rect 426900 159468 426952 159520
rect 429384 159468 429436 159520
rect 446864 159468 446916 159520
rect 457996 159536 458048 159588
rect 469128 159536 469180 159588
rect 469312 159536 469364 159588
rect 474740 159536 474792 159588
rect 459560 159468 459612 159520
rect 462412 159468 462464 159520
rect 468208 159468 468260 159520
rect 479708 159468 479760 159520
rect 485320 159468 485372 159520
rect 388 159400 440 159452
rect 39948 159400 40000 159452
rect 45376 159400 45428 159452
rect 154396 159400 154448 159452
rect 162400 159400 162452 159452
rect 245660 159400 245712 159452
rect 258632 159400 258684 159452
rect 282184 159400 282236 159452
rect 342720 159400 342772 159452
rect 382280 159400 382332 159452
rect 387800 159400 387852 159452
rect 417240 159400 417292 159452
rect 439872 159400 439924 159452
rect 446404 159400 446456 159452
rect 454592 159400 454644 159452
rect 466368 159400 466420 159452
rect 3792 159332 3844 159384
rect 34520 159332 34572 159384
rect 38476 159332 38528 159384
rect 154488 159332 154540 159384
rect 155500 159332 155552 159384
rect 245200 159332 245252 159384
rect 252560 159332 252612 159384
rect 310244 159332 310296 159384
rect 315028 159332 315080 159384
rect 363328 159332 363380 159384
rect 373908 159332 373960 159384
rect 406752 159332 406804 159384
rect 407764 159332 407816 159384
rect 432052 159332 432104 159384
rect 453672 159332 453724 159384
rect 463700 159332 463752 159384
rect 473636 159332 473688 159384
rect 478972 159332 479024 159384
rect 48044 159264 48096 159316
rect 100944 159264 100996 159316
rect 106924 159264 106976 159316
rect 198740 159264 198792 159316
rect 244832 159264 244884 159316
rect 272432 159264 272484 159316
rect 276020 159264 276072 159316
rect 293960 159264 294012 159316
rect 296812 159264 296864 159316
rect 332600 159264 332652 159316
rect 345388 159264 345440 159316
rect 379520 159264 379572 159316
rect 456340 159264 456392 159316
rect 467748 159264 467800 159316
rect 99196 159196 99248 159248
rect 138020 159196 138072 159248
rect 148600 159196 148652 159248
rect 238668 159196 238720 159248
rect 269028 159196 269080 159248
rect 291108 159196 291160 159248
rect 303712 159196 303764 159248
rect 339408 159196 339460 159248
rect 349712 159196 349764 159248
rect 360200 159196 360252 159248
rect 373080 159196 373132 159248
rect 388444 159196 388496 159248
rect 455420 159196 455472 159248
rect 467380 159196 467432 159248
rect 12440 159128 12492 159180
rect 13820 159128 13872 159180
rect 251732 159128 251784 159180
rect 272064 159128 272116 159180
rect 289820 159128 289872 159180
rect 308312 159128 308364 159180
rect 310704 159128 310756 159180
rect 346308 159128 346360 159180
rect 366180 159128 366232 159180
rect 378048 159128 378100 159180
rect 457168 159128 457220 159180
rect 468668 159128 468720 159180
rect 234344 159060 234396 159112
rect 253204 159060 253256 159112
rect 272524 159060 272576 159112
rect 283012 159060 283064 159112
rect 293316 159060 293368 159112
rect 322940 159060 322992 159112
rect 444196 159060 444248 159112
rect 447232 159060 447284 159112
rect 464068 159060 464120 159112
rect 469312 159060 469364 159112
rect 474464 159060 474516 159112
rect 478880 159060 478932 159112
rect 223948 158992 224000 159044
rect 231768 158992 231820 159044
rect 248236 158992 248288 159044
rect 251088 158992 251140 159044
rect 282920 158992 282972 159044
rect 311072 158992 311124 159044
rect 317604 158992 317656 159044
rect 342260 158992 342312 159044
rect 384396 158992 384448 159044
rect 390560 158992 390612 159044
rect 459744 158992 459796 159044
rect 465632 158992 465684 159044
rect 471060 158992 471112 159044
rect 476396 158992 476448 159044
rect 480536 158992 480588 159044
rect 485964 158992 486016 159044
rect 287244 158924 287296 158976
rect 342812 158924 342864 158976
rect 435456 158924 435508 158976
rect 442816 158924 442868 158976
rect 466736 158924 466788 158976
rect 473268 158924 473320 158976
rect 481456 158924 481508 158976
rect 486608 158924 486660 158976
rect 487528 158924 487580 158976
rect 488632 158924 488684 158976
rect 507124 158924 507176 158976
rect 509148 158924 509200 158976
rect 509700 158924 509752 158976
rect 512644 158924 512696 158976
rect 533160 158924 533212 158976
rect 537760 158924 537812 158976
rect 237840 158856 237892 158908
rect 240048 158856 240100 158908
rect 463240 158856 463292 158908
rect 468116 158856 468168 158908
rect 472808 158856 472860 158908
rect 477500 158856 477552 158908
rect 482284 158856 482336 158908
rect 487252 158856 487304 158908
rect 489276 158856 489328 158908
rect 491208 158856 491260 158908
rect 492680 158856 492732 158908
rect 494980 158856 495032 158908
rect 506480 158856 506532 158908
rect 508320 158856 508372 158908
rect 508412 158856 508464 158908
rect 510896 158856 510948 158908
rect 532700 158856 532752 158908
rect 535184 158856 535236 158908
rect 94872 158788 94924 158840
rect 97816 158788 97868 158840
rect 318432 158788 318484 158840
rect 324320 158788 324372 158840
rect 377404 158788 377456 158840
rect 379428 158788 379480 158840
rect 398196 158788 398248 158840
rect 399392 158788 399444 158840
rect 403440 158788 403492 158840
rect 405648 158788 405700 158840
rect 426808 158788 426860 158840
rect 429384 158788 429436 158840
rect 446772 158788 446824 158840
rect 451740 158788 451792 158840
rect 461492 158788 461544 158840
rect 466828 158788 466880 158840
rect 467564 158788 467616 158840
rect 473176 158788 473228 158840
rect 477132 158788 477184 158840
rect 482008 158788 482060 158840
rect 484860 158788 484912 158840
rect 486976 158788 487028 158840
rect 491852 158788 491904 158840
rect 493968 158788 494020 158840
rect 494428 158788 494480 158840
rect 496268 158788 496320 158840
rect 497004 158788 497056 158840
rect 498200 158788 498252 158840
rect 504548 158788 504600 158840
rect 505744 158788 505796 158840
rect 505836 158788 505888 158840
rect 507400 158788 507452 158840
rect 507768 158788 507820 158840
rect 510068 158788 510120 158840
rect 510988 158788 511040 158840
rect 514392 158788 514444 158840
rect 520556 158788 520608 158840
rect 522212 158788 522264 158840
rect 523132 158788 523184 158840
rect 525616 158788 525668 158840
rect 532792 158788 532844 158840
rect 536932 158788 536984 158840
rect 41972 158720 42024 158772
rect 46388 158720 46440 158772
rect 142528 158720 142580 158772
rect 143264 158720 143316 158772
rect 172888 158720 172940 158772
rect 173348 158720 173400 158772
rect 186688 158720 186740 158772
rect 187608 158720 187660 158772
rect 212724 158720 212776 158772
rect 213644 158720 213696 158772
rect 214472 158720 214524 158772
rect 215116 158720 215168 158772
rect 230940 158720 230992 158772
rect 127808 158652 127860 158704
rect 224592 158652 224644 158704
rect 247408 158720 247460 158772
rect 247960 158720 248012 158772
rect 261300 158720 261352 158772
rect 261944 158720 261996 158772
rect 290740 158720 290792 158772
rect 292764 158720 292816 158772
rect 307208 158720 307260 158772
rect 308864 158720 308916 158772
rect 311532 158720 311584 158772
rect 313740 158720 313792 158772
rect 314108 158720 314160 158772
rect 318708 158720 318760 158772
rect 321100 158720 321152 158772
rect 321744 158720 321796 158772
rect 328000 158720 328052 158772
rect 330760 158720 330812 158772
rect 346216 158720 346268 158772
rect 352472 158720 352524 158772
rect 363512 158720 363564 158772
rect 366272 158720 366324 158772
rect 382648 158720 382700 158772
rect 384212 158720 384264 158772
rect 396448 158720 396500 158772
rect 301044 158652 301096 158704
rect 312360 158652 312412 158704
rect 361396 158652 361448 158704
rect 427728 158720 427780 158772
rect 430580 158720 430632 158772
rect 445024 158720 445076 158772
rect 447140 158720 447192 158772
rect 464988 158720 465040 158772
rect 469220 158720 469272 158772
rect 476212 158720 476264 158772
rect 482744 158720 482796 158772
rect 483204 158720 483256 158772
rect 485504 158720 485556 158772
rect 485780 158720 485832 158772
rect 487804 158720 487856 158772
rect 490104 158720 490156 158772
rect 491576 158720 491628 158772
rect 493600 158720 493652 158772
rect 495256 158720 495308 158772
rect 496176 158720 496228 158772
rect 497556 158720 497608 158772
rect 497924 158720 497976 158772
rect 498844 158720 498896 158772
rect 503260 158720 503312 158772
rect 503720 158720 503772 158772
rect 503904 158720 503956 158772
rect 504824 158720 504876 158772
rect 505192 158720 505244 158772
rect 506572 158720 506624 158772
rect 509056 158720 509108 158772
rect 511816 158720 511868 158772
rect 521660 158720 521712 158772
rect 523868 158720 523920 158772
rect 527180 158720 527232 158772
rect 530860 158720 530912 158772
rect 531412 158720 531464 158772
rect 533436 158720 533488 158772
rect 538680 158763 538732 158772
rect 538680 158729 538689 158763
rect 538689 158729 538723 158763
rect 538723 158729 538732 158763
rect 538680 158720 538732 158729
rect 539508 158763 539560 158772
rect 539508 158729 539517 158763
rect 539517 158729 539551 158763
rect 539551 158729 539560 158763
rect 539508 158720 539560 158729
rect 34520 158584 34572 158636
rect 132776 158584 132828 158636
rect 133880 158584 133932 158636
rect 229100 158584 229152 158636
rect 230020 158584 230072 158636
rect 300400 158584 300452 158636
rect 305460 158584 305512 158636
rect 356244 158584 356296 158636
rect 364432 158584 364484 158636
rect 399944 158584 399996 158636
rect 119988 158516 120040 158568
rect 218888 158516 218940 158568
rect 219624 158516 219676 158568
rect 292672 158516 292724 158568
rect 301964 158516 302016 158568
rect 353668 158516 353720 158568
rect 358360 158516 358412 158568
rect 395436 158516 395488 158568
rect 102600 158448 102652 158500
rect 206008 158448 206060 158500
rect 206652 158448 206704 158500
rect 283104 158448 283156 158500
rect 295064 158448 295116 158500
rect 348516 158448 348568 158500
rect 354036 158448 354088 158500
rect 392216 158448 392268 158500
rect 76656 158380 76708 158432
rect 186504 158380 186556 158432
rect 189356 158380 189408 158432
rect 270224 158380 270276 158432
rect 276848 158380 276900 158432
rect 281448 158380 281500 158432
rect 286416 158380 286468 158432
rect 340788 158380 340840 158432
rect 350540 158380 350592 158432
rect 389640 158380 389692 158432
rect 423680 158380 423732 158432
rect 59360 158312 59412 158364
rect 173900 158312 173952 158364
rect 178868 158312 178920 158364
rect 262496 158312 262548 158364
rect 270408 158312 270460 158364
rect 279240 158312 279292 158364
rect 281172 158312 281224 158364
rect 338304 158312 338356 158364
rect 344468 158312 344520 158364
rect 384948 158312 385000 158364
rect 389548 158312 389600 158364
rect 418528 158312 418580 158364
rect 51448 158244 51500 158296
rect 168104 158244 168156 158296
rect 52460 158176 52512 158228
rect 168748 158244 168800 158296
rect 175464 158244 175516 158296
rect 259920 158244 259972 158296
rect 268200 158244 268252 158296
rect 328644 158244 328696 158296
rect 334072 158244 334124 158296
rect 377404 158244 377456 158296
rect 378324 158244 378376 158296
rect 410156 158244 410208 158296
rect 168472 158176 168524 158228
rect 254032 158176 254084 158228
rect 254308 158176 254360 158228
rect 318340 158176 318392 158228
rect 322848 158176 322900 158228
rect 369124 158176 369176 158228
rect 375656 158176 375708 158228
rect 408224 158176 408276 158228
rect 15108 158108 15160 158160
rect 141148 158108 141200 158160
rect 147680 158108 147732 158160
rect 239404 158108 239456 158160
rect 250904 158108 250956 158160
rect 315764 158108 315816 158160
rect 320180 158108 320232 158160
rect 367192 158108 367244 158160
rect 368756 158108 368808 158160
rect 403164 158108 403216 158160
rect 406016 158108 406068 158160
rect 430764 158108 430816 158160
rect 10784 158040 10836 158092
rect 137928 158040 137980 158092
rect 144276 158040 144328 158092
rect 236828 158040 236880 158092
rect 240048 158040 240100 158092
rect 306196 158040 306248 158092
rect 308956 158040 309008 158092
rect 358820 158040 358872 158092
rect 359188 158040 359240 158092
rect 394608 158040 394660 158092
rect 395620 158040 395672 158092
rect 423036 158040 423088 158092
rect 423404 158040 423456 158092
rect 443552 158040 443604 158092
rect 7288 157972 7340 158024
rect 135352 157972 135404 158024
rect 140780 157972 140832 158024
rect 234252 157972 234304 158024
rect 243912 157972 243964 158024
rect 310704 157972 310756 158024
rect 315856 157972 315908 158024
rect 363972 157972 364024 158024
rect 365260 157972 365312 158024
rect 39948 157904 40000 157956
rect 130292 157904 130344 157956
rect 130384 157904 130436 157956
rect 226524 157904 226576 157956
rect 257804 157904 257856 157956
rect 320916 157904 320968 157956
rect 347964 157904 348016 157956
rect 387708 157904 387760 157956
rect 400220 157972 400272 158024
rect 426256 157972 426308 158024
rect 443276 157972 443328 158024
rect 458364 157972 458416 158024
rect 400588 157904 400640 157956
rect 80060 157836 80112 157888
rect 155960 157836 156012 157888
rect 158076 157836 158128 157888
rect 247132 157836 247184 157888
rect 260564 157836 260616 157888
rect 275376 157836 275428 157888
rect 291568 157836 291620 157888
rect 345940 157836 345992 157888
rect 356612 157836 356664 157888
rect 357624 157836 357676 157888
rect 224960 157768 225012 157820
rect 288164 157768 288216 157820
rect 318708 157768 318760 157820
rect 362592 157768 362644 157820
rect 283840 157700 283892 157752
rect 285680 157700 285732 157752
rect 339408 157700 339460 157752
rect 354956 157700 355008 157752
rect 341892 157632 341944 157684
rect 343548 157632 343600 157684
rect 254032 157360 254084 157412
rect 254768 157360 254820 157412
rect 531964 157360 532016 157412
rect 535460 157360 535512 157412
rect 108672 157292 108724 157344
rect 210516 157292 210568 157344
rect 217048 157292 217100 157344
rect 290740 157292 290792 157344
rect 327172 157292 327224 157344
rect 372344 157292 372396 157344
rect 379152 157292 379204 157344
rect 408500 157292 408552 157344
rect 103520 157224 103572 157276
rect 106096 157156 106148 157208
rect 205824 157224 205876 157276
rect 282460 157224 282512 157276
rect 283012 157224 283064 157276
rect 331864 157224 331916 157276
rect 335820 157224 335872 157276
rect 337200 157224 337252 157276
rect 348792 157224 348844 157276
rect 388352 157224 388404 157276
rect 388444 157224 388496 157276
rect 406384 157224 406436 157276
rect 206652 157156 206704 157208
rect 209228 157156 209280 157208
rect 284944 157156 284996 157208
rect 316776 157156 316828 157208
rect 364616 157156 364668 157208
rect 367836 157156 367888 157208
rect 402428 157156 402480 157208
rect 28908 157088 28960 157140
rect 134064 157088 134116 157140
rect 137284 157088 137336 157140
rect 231676 157088 231728 157140
rect 231768 157088 231820 157140
rect 295800 157088 295852 157140
rect 306380 157088 306432 157140
rect 356888 157088 356940 157140
rect 360936 157088 360988 157140
rect 397368 157088 397420 157140
rect 81808 157020 81860 157072
rect 190644 157020 190696 157072
rect 202328 157020 202380 157072
rect 279884 157020 279936 157072
rect 299388 157020 299440 157072
rect 351736 157020 351788 157072
rect 357440 157020 357492 157072
rect 394792 157020 394844 157072
rect 74908 156952 74960 157004
rect 185492 156952 185544 157004
rect 192760 156952 192812 157004
rect 272800 156952 272852 157004
rect 295892 156952 295944 157004
rect 349160 156952 349212 157004
rect 355784 156952 355836 157004
rect 393504 156952 393556 157004
rect 410340 156952 410392 157004
rect 429200 156952 429252 157004
rect 78312 156884 78364 156936
rect 188068 156884 188120 156936
rect 191932 156884 191984 156936
rect 272156 156884 272208 156936
rect 61016 156816 61068 156868
rect 175188 156816 175240 156868
rect 183560 156816 183612 156868
rect 184848 156816 184900 156868
rect 188436 156816 188488 156868
rect 269580 156816 269632 156868
rect 276112 156816 276164 156868
rect 285588 156884 285640 156936
rect 288992 156884 289044 156936
rect 285496 156816 285548 156868
rect 341524 156884 341576 156936
rect 347044 156884 347096 156936
rect 387064 156884 387116 156936
rect 402520 156884 402572 156936
rect 428188 156884 428240 156936
rect 340972 156816 341024 156868
rect 382556 156816 382608 156868
rect 392124 156816 392176 156868
rect 420460 156816 420512 156868
rect 438952 156816 439004 156868
rect 455144 156816 455196 156868
rect 22836 156748 22888 156800
rect 146944 156748 146996 156800
rect 154672 156748 154724 156800
rect 244556 156748 244608 156800
rect 248512 156748 248564 156800
rect 249708 156748 249760 156800
rect 258080 156748 258132 156800
rect 259276 156748 259328 156800
rect 278596 156748 278648 156800
rect 336372 156748 336424 156800
rect 337568 156748 337620 156800
rect 379980 156748 380032 156800
rect 386420 156748 386472 156800
rect 415952 156748 416004 156800
rect 420736 156748 420788 156800
rect 440240 156748 440292 156800
rect 6368 156680 6420 156732
rect 134708 156680 134760 156732
rect 143356 156680 143408 156732
rect 233516 156680 233568 156732
rect 240416 156680 240468 156732
rect 308128 156680 308180 156732
rect 309784 156680 309836 156732
rect 313280 156680 313332 156732
rect 362040 156680 362092 156732
rect 372252 156680 372304 156732
rect 405740 156680 405792 156732
rect 417332 156680 417384 156732
rect 439044 156680 439096 156732
rect 441528 156680 441580 156732
rect 457076 156680 457128 156732
rect 2044 156612 2096 156664
rect 131488 156612 131540 156664
rect 136456 156612 136508 156664
rect 231032 156612 231084 156664
rect 302976 156612 303028 156664
rect 359464 156612 359516 156664
rect 361856 156612 361908 156664
rect 398012 156612 398064 156664
rect 399116 156612 399168 156664
rect 425612 156612 425664 156664
rect 434628 156612 434680 156664
rect 449900 156612 449952 156664
rect 99380 156544 99432 156596
rect 194692 156544 194744 156596
rect 195704 156544 195756 156596
rect 198832 156544 198884 156596
rect 277308 156544 277360 156596
rect 282184 156544 282236 156596
rect 321560 156544 321612 156596
rect 330576 156544 330628 156596
rect 374920 156544 374972 156596
rect 123392 156476 123444 156528
rect 221464 156476 221516 156528
rect 223396 156476 223448 156528
rect 295248 156476 295300 156528
rect 308312 156476 308364 156528
rect 344744 156476 344796 156528
rect 165620 156408 165672 156460
rect 166816 156408 166868 156460
rect 183468 156408 183520 156460
rect 191288 156408 191340 156460
rect 197636 156408 197688 156460
rect 208584 156408 208636 156460
rect 236184 156408 236236 156460
rect 253204 156408 253256 156460
rect 303620 156408 303672 156460
rect 344100 156408 344152 156460
rect 272064 156340 272116 156392
rect 316408 156340 316460 156392
rect 342260 156340 342312 156392
rect 365260 156408 365312 156460
rect 272432 156272 272484 156324
rect 311348 156272 311400 156324
rect 174084 155932 174136 155984
rect 176476 155932 176528 155984
rect 356428 155932 356480 155984
rect 358176 155932 358228 155984
rect 397276 155932 397328 155984
rect 401876 155932 401928 155984
rect 120816 155864 120868 155916
rect 219532 155864 219584 155916
rect 226616 155864 226668 155916
rect 297824 155864 297876 155916
rect 326252 155864 326304 155916
rect 371700 155864 371752 155916
rect 378048 155864 378100 155916
rect 401232 155864 401284 155916
rect 430580 155864 430632 155916
rect 446772 155864 446824 155916
rect 446864 155864 446916 155916
rect 448060 155864 448112 155916
rect 122564 155796 122616 155848
rect 220820 155796 220872 155848
rect 220912 155796 220964 155848
rect 293316 155796 293368 155848
rect 297640 155796 297692 155848
rect 298100 155796 298152 155848
rect 302884 155796 302936 155848
rect 354312 155796 354364 155848
rect 362684 155796 362736 155848
rect 398656 155796 398708 155848
rect 437480 155796 437532 155848
rect 449348 155796 449400 155848
rect 41420 155728 41472 155780
rect 144368 155728 144420 155780
rect 150348 155728 150400 155780
rect 241336 155728 241388 155780
rect 245660 155728 245712 155780
rect 250352 155728 250404 155780
rect 275100 155728 275152 155780
rect 333796 155728 333848 155780
rect 334900 155728 334952 155780
rect 351920 155728 351972 155780
rect 354864 155728 354916 155780
rect 392860 155728 392912 155780
rect 413836 155728 413888 155780
rect 429384 155728 429436 155780
rect 446128 155728 446180 155780
rect 446404 155728 446456 155780
rect 455788 155728 455840 155780
rect 92204 155660 92256 155712
rect 198280 155660 198332 155712
rect 198740 155660 198792 155712
rect 209228 155660 209280 155712
rect 216220 155660 216272 155712
rect 290096 155660 290148 155712
rect 298560 155660 298612 155712
rect 351092 155660 351144 155712
rect 351368 155660 351420 155712
rect 390284 155660 390336 155712
rect 405648 155660 405700 155712
rect 428832 155660 428884 155712
rect 430304 155660 430356 155712
rect 448704 155660 448756 155712
rect 85304 155592 85356 155644
rect 193128 155592 193180 155644
rect 197360 155592 197412 155644
rect 204076 155592 204128 155644
rect 204904 155592 204956 155644
rect 281816 155592 281868 155644
rect 282092 155592 282144 155644
rect 338948 155592 339000 155644
rect 343640 155592 343692 155644
rect 384488 155592 384540 155644
rect 393320 155592 393372 155644
rect 421104 155592 421156 155644
rect 424232 155592 424284 155644
rect 444196 155592 444248 155644
rect 447232 155592 447284 155644
rect 459008 155592 459060 155644
rect 67916 155524 67968 155576
rect 180340 155524 180392 155576
rect 195336 155524 195388 155576
rect 274732 155524 274784 155576
rect 277768 155524 277820 155576
rect 335728 155524 335780 155576
rect 340144 155524 340196 155576
rect 381912 155524 381964 155576
rect 388720 155524 388772 155576
rect 417884 155524 417936 155576
rect 419908 155524 419960 155576
rect 440976 155524 441028 155576
rect 447140 155524 447192 155576
rect 459652 155524 459704 155576
rect 57520 155456 57572 155508
rect 172612 155456 172664 155508
rect 181536 155456 181588 155508
rect 264428 155456 264480 155508
rect 270776 155456 270828 155508
rect 330576 155456 330628 155508
rect 336648 155456 336700 155508
rect 379336 155456 379388 155508
rect 384212 155456 384264 155508
rect 413376 155456 413428 155508
rect 44548 155388 44600 155440
rect 162952 155388 163004 155440
rect 171416 155388 171468 155440
rect 256700 155388 256752 155440
rect 267372 155388 267424 155440
rect 328000 155388 328052 155440
rect 333244 155388 333296 155440
rect 376760 155388 376812 155440
rect 385224 155388 385276 155440
rect 415308 155388 415360 155440
rect 29828 155320 29880 155372
rect 152096 155320 152148 155372
rect 165068 155320 165120 155372
rect 252284 155320 252336 155372
rect 260380 155320 260432 155372
rect 322848 155320 322900 155372
rect 329748 155320 329800 155372
rect 374276 155320 374328 155372
rect 381728 155320 381780 155372
rect 412732 155320 412784 155372
rect 412916 155320 412968 155372
rect 435916 155456 435968 155508
rect 445668 155456 445720 155508
rect 457720 155456 457772 155508
rect 416412 155388 416464 155440
rect 438400 155388 438452 155440
rect 440700 155388 440752 155440
rect 456432 155388 456484 155440
rect 436560 155320 436612 155372
rect 438124 155320 438176 155372
rect 454500 155320 454552 155372
rect 25504 155252 25556 155304
rect 148876 155252 148928 155304
rect 151176 155252 151228 155304
rect 241980 155252 242032 155304
rect 261944 155252 261996 155304
rect 323492 155252 323544 155304
rect 323676 155252 323728 155304
rect 369768 155252 369820 155304
rect 371332 155252 371384 155304
rect 405096 155252 405148 155304
rect 407120 155252 407172 155304
rect 431408 155252 431460 155304
rect 437204 155252 437256 155304
rect 453856 155252 453908 155304
rect 13820 155184 13872 155236
rect 139216 155184 139268 155236
rect 145104 155184 145156 155236
rect 237472 155184 237524 155236
rect 247960 155184 248012 155236
rect 313280 155184 313332 155236
rect 319352 155184 319404 155236
rect 366548 155184 366600 155236
rect 369584 155184 369636 155236
rect 372620 155184 372672 155236
rect 374828 155184 374880 155236
rect 407580 155184 407632 155236
rect 409512 155184 409564 155236
rect 433340 155184 433392 155236
rect 433800 155184 433852 155236
rect 451280 155184 451332 155236
rect 129464 155116 129516 155168
rect 225880 155116 225932 155168
rect 237012 155116 237064 155168
rect 305552 155116 305604 155168
rect 311072 155116 311124 155168
rect 339592 155116 339644 155168
rect 352288 155116 352340 155168
rect 387800 155116 387852 155168
rect 175832 155048 175884 155100
rect 186136 155048 186188 155100
rect 186228 155048 186280 155100
rect 196348 155048 196400 155100
rect 213644 155048 213696 155100
rect 287520 155048 287572 155100
rect 288256 155048 288308 155100
rect 343456 155048 343508 155100
rect 346308 155048 346360 155100
rect 360108 155048 360160 155100
rect 372712 155048 372764 155100
rect 375564 155048 375616 155100
rect 116492 154980 116544 155032
rect 216312 154980 216364 155032
rect 293960 154980 294012 155032
rect 334440 154980 334492 155032
rect 332600 154912 332652 154964
rect 349804 154912 349856 154964
rect 225052 154776 225104 154828
rect 227168 154776 227220 154828
rect 264980 154776 265032 154828
rect 267648 154776 267700 154828
rect 238760 154572 238812 154624
rect 240048 154572 240100 154624
rect 231584 154504 231636 154556
rect 301688 154504 301740 154556
rect 301780 154504 301832 154556
rect 311992 154504 312044 154556
rect 313740 154504 313792 154556
rect 360752 154504 360804 154556
rect 376668 154504 376720 154556
rect 380624 154504 380676 154556
rect 385960 154504 386012 154556
rect 391572 154504 391624 154556
rect 391940 154504 391992 154556
rect 408868 154504 408920 154556
rect 456892 154504 456944 154556
rect 460296 154504 460348 154556
rect 462228 154504 462280 154556
rect 463516 154504 463568 154556
rect 473268 154504 473320 154556
rect 475660 154504 475712 154556
rect 475752 154504 475804 154556
rect 478236 154504 478288 154556
rect 487804 154504 487856 154556
rect 489828 154504 489880 154556
rect 491576 154504 491628 154556
rect 493048 154504 493100 154556
rect 495440 154504 495492 154556
rect 496912 154504 496964 154556
rect 498752 154504 498804 154556
rect 499488 154504 499540 154556
rect 512276 154504 512328 154556
rect 516140 154504 516192 154556
rect 520004 154504 520056 154556
rect 525800 154504 525852 154556
rect 527732 154504 527784 154556
rect 532792 154504 532844 154556
rect 224868 154436 224920 154488
rect 296536 154436 296588 154488
rect 296628 154436 296680 154488
rect 308864 154436 308916 154488
rect 357532 154436 357584 154488
rect 360200 154436 360252 154488
rect 388996 154436 389048 154488
rect 390560 154436 390612 154488
rect 414664 154436 414716 154488
rect 486976 154436 487028 154488
rect 489184 154436 489236 154488
rect 510344 154436 510396 154488
rect 513472 154436 513524 154488
rect 513564 154436 513616 154488
rect 517612 154436 517664 154488
rect 521292 154436 521344 154488
rect 528284 154436 528336 154488
rect 528376 154436 528428 154488
rect 533160 154436 533212 154488
rect 217876 154368 217928 154420
rect 291384 154368 291436 154420
rect 291844 154368 291896 154420
rect 304264 154368 304316 154420
rect 304908 154368 304960 154420
rect 355600 154368 355652 154420
rect 366916 154368 366968 154420
rect 368480 154368 368532 154420
rect 372620 154368 372672 154420
rect 403808 154368 403860 154420
rect 415584 154368 415636 154420
rect 437848 154368 437900 154420
rect 471888 154368 471940 154420
rect 475016 154368 475068 154420
rect 476120 154368 476172 154420
rect 479524 154368 479576 154420
rect 512920 154368 512972 154420
rect 516968 154368 517020 154420
rect 34428 154300 34480 154352
rect 155316 154300 155368 154352
rect 215116 154300 215168 154352
rect 288808 154300 288860 154352
rect 298100 154300 298152 154352
rect 350448 154300 350500 154352
rect 366272 154300 366324 154352
rect 399300 154300 399352 154352
rect 399392 154300 399444 154352
rect 424968 154300 425020 154352
rect 428556 154300 428608 154352
rect 447416 154300 447468 154352
rect 514208 154300 514260 154352
rect 518716 154368 518768 154420
rect 519360 154368 519412 154420
rect 523132 154368 523184 154420
rect 524512 154368 524564 154420
rect 531780 154368 531832 154420
rect 518072 154300 518124 154352
rect 521660 154300 521712 154352
rect 525800 154300 525852 154352
rect 533988 154300 534040 154352
rect 30656 154232 30708 154284
rect 152740 154232 152792 154284
rect 210976 154232 211028 154284
rect 286232 154232 286284 154284
rect 289728 154232 289780 154284
rect 299112 154232 299164 154284
rect 300308 154232 300360 154284
rect 352380 154232 352432 154284
rect 352472 154232 352524 154284
rect 386420 154232 386472 154284
rect 394608 154232 394660 154284
rect 396080 154232 396132 154284
rect 404268 154232 404320 154284
rect 429476 154232 429528 154284
rect 436008 154232 436060 154284
rect 465632 154232 465684 154284
rect 470508 154232 470560 154284
rect 473728 154232 473780 154284
rect 476948 154232 477000 154284
rect 477500 154232 477552 154284
rect 480168 154232 480220 154284
rect 491300 154232 491352 154284
rect 493692 154232 493744 154284
rect 511632 154232 511684 154284
rect 514760 154232 514812 154284
rect 525156 154232 525208 154284
rect 531412 154232 531464 154284
rect 27528 154164 27580 154216
rect 150164 154164 150216 154216
rect 207480 154164 207532 154216
rect 283748 154164 283800 154216
rect 292764 154164 292816 154216
rect 345388 154164 345440 154216
rect 350172 154164 350224 154216
rect 353024 154164 353076 154216
rect 357624 154164 357676 154216
rect 394148 154164 394200 154216
rect 397460 154164 397512 154216
rect 424324 154164 424376 154216
rect 425060 154164 425112 154216
rect 444840 154164 444892 154216
rect 518716 154164 518768 154216
rect 524788 154164 524840 154216
rect 526444 154164 526496 154216
rect 532700 154164 532752 154216
rect 23756 154096 23808 154148
rect 147588 154096 147640 154148
rect 154488 154096 154540 154148
rect 158536 154096 158588 154148
rect 204168 154096 204220 154148
rect 281172 154096 281224 154148
rect 281448 154096 281500 154148
rect 335084 154096 335136 154148
rect 337200 154096 337252 154148
rect 20628 154028 20680 154080
rect 145012 154028 145064 154080
rect 200580 154028 200632 154080
rect 278596 154028 278648 154080
rect 285680 154028 285732 154080
rect 340236 154028 340288 154080
rect 340788 154096 340840 154148
rect 342168 154096 342220 154148
rect 378692 154096 378744 154148
rect 391296 154096 391348 154148
rect 419816 154096 419868 154148
rect 422484 154096 422536 154148
rect 442908 154096 442960 154148
rect 462136 154096 462188 154148
rect 464160 154096 464212 154148
rect 473176 154096 473228 154148
rect 476304 154096 476356 154148
rect 485504 154096 485556 154148
rect 487896 154096 487948 154148
rect 491208 154096 491260 154148
rect 492404 154096 492456 154148
rect 517428 154096 517480 154148
rect 523040 154096 523092 154148
rect 523868 154096 523920 154148
rect 531320 154096 531372 154148
rect 343548 154028 343600 154080
rect 383200 154028 383252 154080
rect 390376 154028 390428 154080
rect 419172 154028 419224 154080
rect 419264 154028 419316 154080
rect 440332 154028 440384 154080
rect 442816 154028 442868 154080
rect 452568 154028 452620 154080
rect 469312 154028 469364 154080
rect 473728 154028 473780 154080
rect 523224 154028 523276 154080
rect 527180 154028 527232 154080
rect 16856 153960 16908 154012
rect 142436 153960 142488 154012
rect 187608 153960 187660 154012
rect 268292 153960 268344 154012
rect 269948 153960 270000 154012
rect 329932 153960 329984 154012
rect 332324 153960 332376 154012
rect 376208 153960 376260 154012
rect 379428 153960 379480 154012
rect 409512 153960 409564 154012
rect 411260 153960 411312 154012
rect 434628 153960 434680 154012
rect 436376 153960 436428 154012
rect 13728 153892 13780 153944
rect 139860 153892 139912 153944
rect 179788 153892 179840 153944
rect 263140 153892 263192 153944
rect 263232 153892 263284 153944
rect 324780 153892 324832 153944
rect 325424 153892 325476 153944
rect 371056 153892 371108 153944
rect 383476 153892 383528 153944
rect 414020 153892 414072 153944
rect 414756 153892 414808 153944
rect 437204 153892 437256 153944
rect 449992 153960 450044 154012
rect 474740 153960 474792 154012
rect 477592 153960 477644 154012
rect 482008 153960 482060 154012
rect 483388 153960 483440 154012
rect 529664 153960 529716 154012
rect 453212 153892 453264 153944
rect 529020 153892 529072 153944
rect 9864 153824 9916 153876
rect 137284 153824 137336 153876
rect 154396 153824 154448 153876
rect 163596 153824 163648 153876
rect 169484 153824 169536 153876
rect 255412 153824 255464 153876
rect 256056 153824 256108 153876
rect 319628 153824 319680 153876
rect 321744 153824 321796 153876
rect 367836 153824 367888 153876
rect 370504 153824 370556 153876
rect 404452 153824 404504 153876
rect 408500 153824 408552 153876
rect 410800 153824 410852 153876
rect 242164 153756 242216 153808
rect 309416 153756 309468 153808
rect 316224 153756 316276 153808
rect 327356 153756 327408 153808
rect 330760 153756 330812 153808
rect 372988 153756 373040 153808
rect 405188 153756 405240 153808
rect 430120 153824 430172 153876
rect 433248 153824 433300 153876
rect 450636 153824 450688 153876
rect 451740 153824 451792 153876
rect 460940 153824 460992 153876
rect 463700 153824 463752 153876
rect 466092 153824 466144 153876
rect 469220 153824 469272 153876
rect 474372 153824 474424 153876
rect 527088 153824 527140 153876
rect 535552 153824 535604 153876
rect 249156 153688 249208 153740
rect 314568 153688 314620 153740
rect 324320 153688 324372 153740
rect 365904 153688 365956 153740
rect 415216 153688 415268 153740
rect 416596 153688 416648 153740
rect 280988 153620 281040 153672
rect 293960 153620 294012 153672
rect 306840 153620 306892 153672
rect 311900 153620 311952 153672
rect 322204 153620 322256 153672
rect 328368 153620 328420 153672
rect 332508 153620 332560 153672
rect 351920 153620 351972 153672
rect 378048 153620 378100 153672
rect 462872 153552 462924 153604
rect 464804 153552 464856 153604
rect 481088 153552 481140 153604
rect 482100 153552 482152 153604
rect 515496 153552 515548 153604
rect 520188 153552 520240 153604
rect 520648 153552 520700 153604
rect 527364 153552 527416 153604
rect 43812 153484 43864 153536
rect 118056 153484 118108 153536
rect 387800 153484 387852 153536
rect 390928 153484 390980 153536
rect 95148 153416 95200 153468
rect 126704 153416 126756 153468
rect 463792 153416 463844 153468
rect 465448 153416 465500 153468
rect 466828 153416 466880 153468
rect 471796 153416 471848 153468
rect 488264 153416 488316 153468
rect 490472 153416 490524 153468
rect 514852 153416 514904 153468
rect 518900 153416 518952 153468
rect 50620 153348 50672 153400
rect 115296 153348 115348 153400
rect 459560 153348 459612 153400
rect 462872 153348 462924 153400
rect 468116 153348 468168 153400
rect 473084 153348 473136 153400
rect 488540 153348 488592 153400
rect 491760 153348 491812 153400
rect 516140 153348 516192 153400
rect 520740 153348 520792 153400
rect 522580 153348 522632 153400
rect 529940 153348 529992 153400
rect 46756 153280 46808 153332
rect 117228 153280 117280 153332
rect 379520 153280 379572 153332
rect 385776 153280 385828 153332
rect 459836 153280 459888 153332
rect 462228 153280 462280 153332
rect 468208 153280 468260 153332
rect 472440 153280 472492 153332
rect 478880 153280 478932 153332
rect 481456 153280 481508 153332
rect 521936 153280 521988 153332
rect 528560 153280 528612 153332
rect 108948 153212 109000 153264
rect 119896 153212 119948 153264
rect 114652 153144 114704 153196
rect 182916 153144 182968 153196
rect 184112 153144 184164 153196
rect 266360 153144 266412 153196
rect 274548 153144 274600 153196
rect 310244 153212 310296 153264
rect 317052 153212 317104 153264
rect 382280 153212 382332 153264
rect 383844 153212 383896 153264
rect 420920 153212 420972 153264
rect 422392 153212 422444 153264
rect 429200 153212 429252 153264
rect 433984 153212 434036 153264
rect 440240 153212 440292 153264
rect 441620 153212 441672 153264
rect 449900 153212 449952 153264
rect 451924 153212 451976 153264
rect 458180 153212 458232 153264
rect 461584 153212 461636 153264
rect 476396 153212 476448 153264
rect 478972 153212 479024 153264
rect 480812 153212 480864 153264
rect 488632 153212 488684 153264
rect 491116 153212 491168 153264
rect 516784 153212 516836 153264
rect 520556 153212 520608 153264
rect 333152 153144 333204 153196
rect 478880 153144 478932 153196
rect 118700 153076 118752 153128
rect 175832 153076 175884 153128
rect 177212 153076 177264 153128
rect 261208 153076 261260 153128
rect 324136 153076 324188 153128
rect 62120 153008 62172 153060
rect 146300 153008 146352 153060
rect 143264 152940 143316 152992
rect 235540 152940 235592 152992
rect 236092 152940 236144 152992
rect 304908 152940 304960 152992
rect 222292 152872 222344 152924
rect 125508 152804 125560 152856
rect 222660 152804 222712 152856
rect 229192 152872 229244 152924
rect 299756 152872 299808 152924
rect 308772 152872 308824 152924
rect 294604 152804 294656 152856
rect 118608 152736 118660 152788
rect 217600 152736 217652 152788
rect 218796 152736 218848 152788
rect 292028 152736 292080 152788
rect 111708 152668 111760 152720
rect 212448 152668 212500 152720
rect 215300 152668 215352 152720
rect 289452 152668 289504 152720
rect 93952 152600 94004 152652
rect 199568 152600 199620 152652
rect 208400 152600 208452 152652
rect 284300 152600 284352 152652
rect 87052 152532 87104 152584
rect 194416 152532 194468 152584
rect 198004 152532 198056 152584
rect 276664 152532 276716 152584
rect 279424 152532 279476 152584
rect 337016 152532 337068 152584
rect 2964 152464 3016 152516
rect 132132 152464 132184 152516
rect 227720 152464 227772 152516
rect 298468 152464 298520 152516
rect 152004 152396 152056 152448
rect 242624 152396 242676 152448
rect 262220 152396 262272 152448
rect 132960 152328 133012 152380
rect 228456 152328 228508 152380
rect 241520 152328 241572 152380
rect 16212 152260 16264 152312
rect 124864 152260 124916 152312
rect 135536 152260 135588 152312
rect 230388 152260 230440 152312
rect 101910 152192 101962 152244
rect 118608 152192 118660 152244
rect 91606 152124 91658 152176
rect 116584 152124 116636 152176
rect 39994 152056 40046 152108
rect 115204 152056 115256 152108
rect 36912 151988 36964 152040
rect 120816 151988 120868 152040
rect 30012 151920 30064 151972
rect 122196 151920 122248 151972
rect 19708 151852 19760 151904
rect 123484 151852 123536 151904
rect 105636 151784 105688 151836
rect 114560 151784 114612 151836
rect 531596 151512 531648 151564
rect 534724 151512 534776 151564
rect 60832 151419 60884 151428
rect 60832 151385 60841 151419
rect 60841 151385 60875 151419
rect 60875 151385 60884 151419
rect 60832 151376 60884 151385
rect 64420 151419 64472 151428
rect 64420 151385 64429 151419
rect 64429 151385 64463 151419
rect 64463 151385 64472 151419
rect 64420 151376 64472 151385
rect 53932 151308 53984 151360
rect 57520 151308 57572 151360
rect 67640 151351 67692 151360
rect 67640 151317 67649 151351
rect 67649 151317 67683 151351
rect 67683 151317 67692 151351
rect 67640 151308 67692 151317
rect 71320 151351 71372 151360
rect 71320 151317 71329 151351
rect 71329 151317 71363 151351
rect 71363 151317 71372 151351
rect 71320 151308 71372 151317
rect 74540 151351 74592 151360
rect 74540 151317 74549 151351
rect 74549 151317 74583 151351
rect 74583 151317 74592 151351
rect 78128 151351 78180 151360
rect 74540 151308 74592 151317
rect 78128 151317 78137 151351
rect 78137 151317 78171 151351
rect 78171 151317 78180 151351
rect 78128 151308 78180 151317
rect 81440 151351 81492 151360
rect 81440 151317 81449 151351
rect 81449 151317 81483 151351
rect 81483 151317 81492 151351
rect 81440 151308 81492 151317
rect 85028 151351 85080 151360
rect 85028 151317 85037 151351
rect 85037 151317 85071 151351
rect 85071 151317 85080 151351
rect 85028 151308 85080 151317
rect 88340 151351 88392 151360
rect 88340 151317 88349 151351
rect 88349 151317 88383 151351
rect 88383 151317 88392 151351
rect 88340 151308 88392 151317
rect 98828 151351 98880 151360
rect 98828 151317 98837 151351
rect 98837 151317 98871 151351
rect 98871 151317 98880 151351
rect 98828 151308 98880 151317
rect 116860 151240 116912 151292
rect 123576 151172 123628 151224
rect 115388 151104 115440 151156
rect 120724 151104 120776 151156
rect 127624 151104 127676 151156
rect 123668 151036 123720 151088
rect 122288 150968 122340 151020
rect 119528 150900 119580 150952
rect 116768 150832 116820 150884
rect 118148 150764 118200 150816
rect 120908 150696 120960 150748
rect 112536 150628 112588 150680
rect 126980 150628 127032 150680
rect 126336 150560 126388 150612
rect 124956 150492 125008 150544
rect 124588 150424 124640 150476
rect 126704 150424 126756 150476
rect 127900 150424 127952 150476
rect 532608 149880 532660 149932
rect 536104 149880 536156 149932
rect 117228 149676 117280 149728
rect 127716 149676 127768 149728
rect 119896 148996 119948 149048
rect 126980 148996 127032 149048
rect 532332 148996 532384 149048
rect 536196 148996 536248 149048
rect 114560 147568 114612 147620
rect 126980 147568 127032 147620
rect 118608 146208 118660 146260
rect 126980 146208 127032 146260
rect 532148 146072 532200 146124
rect 535368 146072 535420 146124
rect 116676 145188 116728 145240
rect 120724 145188 120776 145240
rect 531780 144848 531832 144900
rect 536288 144848 536340 144900
rect 124588 143488 124640 143540
rect 126980 143488 127032 143540
rect 531688 143216 531740 143268
rect 535276 143216 535328 143268
rect 531964 141856 532016 141908
rect 534908 141856 534960 141908
rect 116584 140700 116636 140752
rect 126980 140700 127032 140752
rect 531964 140700 532016 140752
rect 535184 140700 535236 140752
rect 531596 139340 531648 139392
rect 534724 139340 534776 139392
rect 115388 137912 115440 137964
rect 126980 137912 127032 137964
rect 531412 137912 531464 137964
rect 534816 137912 534868 137964
rect 123668 136552 123720 136604
rect 126980 136552 127032 136604
rect 532148 136348 532200 136400
rect 535092 136348 535144 136400
rect 531780 134852 531832 134904
rect 535000 134852 535052 134904
rect 122288 133832 122340 133884
rect 126980 133832 127032 133884
rect 531780 133492 531832 133544
rect 536196 133492 536248 133544
rect 119528 132404 119580 132456
rect 126980 132404 127032 132456
rect 531412 131996 531464 132048
rect 536012 131996 536064 132048
rect 116676 131044 116728 131096
rect 126980 131044 127032 131096
rect 532608 130636 532660 130688
rect 536748 130636 536800 130688
rect 531596 129412 531648 129464
rect 536656 129412 536708 129464
rect 118148 128256 118200 128308
rect 126980 128256 127032 128308
rect 531964 128052 532016 128104
rect 536564 128052 536616 128104
rect 120908 126896 120960 126948
rect 126980 126896 127032 126948
rect 531872 126556 531924 126608
rect 536472 126556 536524 126608
rect 532608 125196 532660 125248
rect 536380 125196 536432 125248
rect 531780 123836 531832 123888
rect 536104 123836 536156 123888
rect 532608 122476 532660 122528
rect 536288 122476 536340 122528
rect 124956 122408 125008 122460
rect 126980 122408 127032 122460
rect 116768 121388 116820 121440
rect 126980 121388 127032 121440
rect 532148 121116 532200 121168
rect 536196 121116 536248 121168
rect 532516 119892 532568 119944
rect 536656 119892 536708 119944
rect 123576 118600 123628 118652
rect 126980 118600 127032 118652
rect 532608 118396 532660 118448
rect 536748 118396 536800 118448
rect 115296 117240 115348 117292
rect 126980 117240 127032 117292
rect 532332 117036 532384 117088
rect 535460 117036 535512 117088
rect 532608 115676 532660 115728
rect 536380 115676 536432 115728
rect 531688 114316 531740 114368
rect 535644 114316 535696 114368
rect 118056 113092 118108 113144
rect 126980 113092 127032 113144
rect 531780 112888 531832 112940
rect 536288 112888 536340 112940
rect 532516 111800 532568 111852
rect 535460 111800 535512 111852
rect 115204 111732 115256 111784
rect 126980 111732 127032 111784
rect 532608 111460 532660 111512
rect 536472 111460 536524 111512
rect 532608 110440 532660 110492
rect 535460 110440 535512 110492
rect 531964 110100 532016 110152
rect 536196 110100 536248 110152
rect 532424 109012 532476 109064
rect 535460 109012 535512 109064
rect 120816 108944 120868 108996
rect 126980 108944 127032 108996
rect 531780 108876 531832 108928
rect 536656 108876 536708 108928
rect 532240 107652 532292 107704
rect 535460 107652 535512 107704
rect 119436 107584 119488 107636
rect 126980 107584 127032 107636
rect 531780 107380 531832 107432
rect 535552 107380 535604 107432
rect 532148 106292 532200 106344
rect 535460 106292 535512 106344
rect 532516 104864 532568 104916
rect 535460 104864 535512 104916
rect 122196 104796 122248 104848
rect 126980 104796 127032 104848
rect 532608 103708 532660 103760
rect 535460 103708 535512 103760
rect 117964 103436 118016 103488
rect 126980 103436 127032 103488
rect 532056 102144 532108 102196
rect 535460 102144 535512 102196
rect 122104 102076 122156 102128
rect 126980 102076 127032 102128
rect 532608 100716 532660 100768
rect 535460 100716 535512 100768
rect 116952 99424 117004 99476
rect 122104 99424 122156 99476
rect 123484 99288 123536 99340
rect 126980 99288 127032 99340
rect 532240 97996 532292 98048
rect 535460 97996 535512 98048
rect 124864 97928 124916 97980
rect 126980 97928 127032 97980
rect 532148 96636 532200 96688
rect 535460 96636 535512 96688
rect 119344 96568 119396 96620
rect 126980 96568 127032 96620
rect 532056 95208 532108 95260
rect 535460 95208 535512 95260
rect 532516 94188 532568 94240
rect 535460 94188 535512 94240
rect 532424 92488 532476 92540
rect 535460 92488 535512 92540
rect 531964 91060 532016 91112
rect 535460 91060 535512 91112
rect 532608 89700 532660 89752
rect 535460 89700 535512 89752
rect 120724 89632 120776 89684
rect 126980 89632 127032 89684
rect 115940 88544 115992 88596
rect 117964 88544 118016 88596
rect 532056 88340 532108 88392
rect 535460 88340 535512 88392
rect 116584 88272 116636 88324
rect 126980 88272 127032 88324
rect 532332 86980 532384 87032
rect 535460 86980 535512 87032
rect 116676 86912 116728 86964
rect 126980 86912 127032 86964
rect 532516 85552 532568 85604
rect 535460 85552 535512 85604
rect 532608 84192 532660 84244
rect 535460 84192 535512 84244
rect 116768 84124 116820 84176
rect 126980 84124 127032 84176
rect 122104 82764 122156 82816
rect 126980 82764 127032 82816
rect 117964 79976 118016 80028
rect 126980 79976 127032 80028
rect 532148 78684 532200 78736
rect 535644 78684 535696 78736
rect 116124 77936 116176 77988
rect 126980 77936 127032 77988
rect 532608 77188 532660 77240
rect 535552 77188 535604 77240
rect 116584 75896 116636 75948
rect 126980 75896 127032 75948
rect 532608 75828 532660 75880
rect 535460 75828 535512 75880
rect 532608 74468 532660 74520
rect 536288 74468 536340 74520
rect 116768 73176 116820 73228
rect 126980 73176 127032 73228
rect 532424 73108 532476 73160
rect 535552 73108 535604 73160
rect 116676 71748 116728 71800
rect 126980 71748 127032 71800
rect 532424 71680 532476 71732
rect 535644 71680 535696 71732
rect 531780 70524 531832 70576
rect 535736 70524 535788 70576
rect 531964 69776 532016 69828
rect 535552 69776 535604 69828
rect 120816 69028 120868 69080
rect 126980 69028 127032 69080
rect 531964 68144 532016 68196
rect 535460 68144 535512 68196
rect 118056 67600 118108 67652
rect 126980 67600 127032 67652
rect 531964 67532 532016 67584
rect 535552 67532 535604 67584
rect 124864 66240 124916 66292
rect 127440 66240 127492 66292
rect 532148 66172 532200 66224
rect 535460 66240 535512 66292
rect 531320 64812 531372 64864
rect 535460 64880 535512 64932
rect 119344 63520 119396 63572
rect 126980 63520 127032 63572
rect 532148 63452 532200 63504
rect 535460 63520 535512 63572
rect 115204 62092 115256 62144
rect 126980 62092 127032 62144
rect 532332 62024 532384 62076
rect 535460 62092 535512 62144
rect 532516 60664 532568 60716
rect 535460 60732 535512 60784
rect 532608 59304 532660 59356
rect 535460 59372 535512 59424
rect 532424 57876 532476 57928
rect 535460 57944 535512 57996
rect 115296 57196 115348 57248
rect 126980 57196 127032 57248
rect 532608 56516 532660 56568
rect 535460 56584 535512 56636
rect 531320 55156 531372 55208
rect 535460 55224 535512 55276
rect 116584 53796 116636 53848
rect 126980 53796 127032 53848
rect 117964 53048 118016 53100
rect 127808 53048 127860 53100
rect 532148 52980 532200 53032
rect 535460 52980 535512 53032
rect 532608 51280 532660 51332
rect 535460 51280 535512 51332
rect 120724 51076 120776 51128
rect 126980 51076 127032 51128
rect 532516 49988 532568 50040
rect 535460 49988 535512 50040
rect 531964 48628 532016 48680
rect 535460 48628 535512 48680
rect 532608 47404 532660 47456
rect 535460 47404 535512 47456
rect 123484 46928 123536 46980
rect 126980 46928 127032 46980
rect 532608 45772 532660 45824
rect 535460 45772 535512 45824
rect 532516 44548 532568 44600
rect 535460 44548 535512 44600
rect 122104 44140 122156 44192
rect 126980 44140 127032 44192
rect 532608 43052 532660 43104
rect 535460 43052 535512 43104
rect 119436 42780 119488 42832
rect 126980 42780 127032 42832
rect 532608 41692 532660 41744
rect 535460 41692 535512 41744
rect 124956 41420 125008 41472
rect 126980 41420 127032 41472
rect 532608 40128 532660 40180
rect 535460 40128 535512 40180
rect 532608 38768 532660 38820
rect 535460 38768 535512 38820
rect 118148 38632 118200 38684
rect 126980 38632 127032 38684
rect 532608 37408 532660 37460
rect 535368 37408 535420 37460
rect 116676 37272 116728 37324
rect 126980 37272 127032 37324
rect 532332 36048 532384 36100
rect 535368 36048 535420 36100
rect 532608 34688 532660 34740
rect 535368 34688 535420 34740
rect 116860 33328 116912 33380
rect 120816 33328 120868 33380
rect 531964 33328 532016 33380
rect 535368 33328 535420 33380
rect 123576 33124 123628 33176
rect 126980 33124 127032 33176
rect 532608 31968 532660 32020
rect 535368 31968 535420 32020
rect 122196 31764 122248 31816
rect 126980 31764 127032 31816
rect 532608 30608 532660 30660
rect 535368 30608 535420 30660
rect 532608 29248 532660 29300
rect 535368 29248 535420 29300
rect 120816 28976 120868 29028
rect 126980 28976 127032 29028
rect 119528 27616 119580 27668
rect 126980 27616 127032 27668
rect 532608 27616 532660 27668
rect 535460 27548 535512 27600
rect 532332 26528 532384 26580
rect 535368 26528 535420 26580
rect 116768 24828 116820 24880
rect 126980 24828 127032 24880
rect 532608 24828 532660 24880
rect 535368 24828 535420 24880
rect 532056 23672 532108 23724
rect 535276 23672 535328 23724
rect 531964 22312 532016 22364
rect 535368 22312 535420 22364
rect 123668 22108 123720 22160
rect 126980 22108 127032 22160
rect 115940 21088 115992 21140
rect 118056 21088 118108 21140
rect 531964 20952 532016 21004
rect 535276 20952 535328 21004
rect 531964 19592 532016 19644
rect 535184 19592 535236 19644
rect 122288 19320 122340 19372
rect 126980 19320 127032 19372
rect 120908 17960 120960 18012
rect 126980 17960 127032 18012
rect 532332 17960 532384 18012
rect 535368 17960 535420 18012
rect 532240 16872 532292 16924
rect 535276 16872 535328 16924
rect 532608 15512 532660 15564
rect 535368 15512 535420 15564
rect 532148 14152 532200 14204
rect 535276 14152 535328 14204
rect 118056 13812 118108 13864
rect 126980 13812 127032 13864
rect 531596 12656 531648 12708
rect 535368 12656 535420 12708
rect 115388 12452 115440 12504
rect 126980 12452 127032 12504
rect 531964 11296 532016 11348
rect 535184 11296 535236 11348
rect 125048 10888 125100 10940
rect 127716 10888 127768 10940
rect 531780 9664 531832 9716
rect 535000 9664 535052 9716
rect 117228 9052 117280 9104
rect 124864 9052 124916 9104
rect 124312 8984 124364 9036
rect 127256 8984 127308 9036
rect 532240 8304 532292 8356
rect 535276 8304 535328 8356
rect 531964 7080 532016 7132
rect 535184 7080 535236 7132
rect 531596 5856 531648 5908
rect 535368 5856 535420 5908
rect 124864 5516 124916 5568
rect 126980 5516 127032 5568
rect 116584 5312 116636 5364
rect 123484 5244 123536 5296
rect 122104 5176 122156 5228
rect 119436 5108 119488 5160
rect 116676 5040 116728 5092
rect 126336 4972 126388 5024
rect 123576 4904 123628 4956
rect 120816 4836 120868 4888
rect 9312 4632 9364 4684
rect 124864 4768 124916 4820
rect 49332 4632 49384 4684
rect 55956 4675 56008 4684
rect 55956 4641 55965 4675
rect 55965 4641 55999 4675
rect 55999 4641 56008 4675
rect 55956 4632 56008 4641
rect 62672 4675 62724 4684
rect 62672 4641 62681 4675
rect 62681 4641 62715 4675
rect 62715 4641 62724 4675
rect 62672 4632 62724 4641
rect 65984 4675 66036 4684
rect 65984 4641 65993 4675
rect 65993 4641 66027 4675
rect 66027 4641 66036 4675
rect 65984 4632 66036 4641
rect 75828 4675 75880 4684
rect 75828 4641 75837 4675
rect 75837 4641 75871 4675
rect 75871 4641 75880 4675
rect 75828 4632 75880 4641
rect 79324 4675 79376 4684
rect 79324 4641 79333 4675
rect 79333 4641 79367 4675
rect 79367 4641 79376 4675
rect 79324 4632 79376 4641
rect 82636 4675 82688 4684
rect 82636 4641 82645 4675
rect 82645 4641 82679 4675
rect 82679 4641 82688 4675
rect 82636 4632 82688 4641
rect 95976 4675 96028 4684
rect 95976 4641 95985 4675
rect 95985 4641 96019 4675
rect 96019 4641 96028 4675
rect 95976 4632 96028 4641
rect 532608 4496 532660 4548
rect 535460 4496 535512 4548
rect 117228 4156 117280 4208
rect 126980 4156 127032 4208
rect 6000 3544 6052 3596
rect 117228 3544 117280 3596
rect 105636 3476 105688 3528
rect 127624 3476 127676 3528
rect 91100 3408 91152 3460
rect 127808 3408 127860 3460
rect 33692 3340 33744 3392
rect 128360 3340 128412 3392
rect 89352 3272 89404 3324
rect 120724 3272 120776 3324
rect 68928 3204 68980 3256
rect 118148 3204 118200 3256
rect 52368 3136 52420 3188
rect 122196 3136 122248 3188
rect 45928 3068 45980 3120
rect 119528 3068 119580 3120
rect 42616 3000 42668 3052
rect 116768 3000 116820 3052
rect 39304 2932 39356 2984
rect 126428 2932 126480 2984
rect 101128 2864 101180 2916
rect 15936 2796 15988 2848
rect 127716 2796 127768 2848
rect 12348 2728 12400 2780
rect 91100 2728 91152 2780
rect 99288 2728 99340 2780
rect 105636 2728 105688 2780
rect 102692 2660 102744 2712
rect 117964 2728 118016 2780
rect 313280 2864 313332 2916
rect 371148 2864 371200 2916
rect 236184 2796 236236 2848
rect 179972 2728 180024 2780
rect 279976 2796 280028 2848
rect 303712 2796 303764 2848
rect 346676 2796 346728 2848
rect 438676 2796 438728 2848
rect 246672 2728 246724 2780
rect 108948 2660 109000 2712
rect 115204 2660 115256 2712
rect 128360 2660 128412 2712
rect 146668 2660 146720 2712
rect 112628 2592 112680 2644
rect 119344 2592 119396 2644
rect 28908 2524 28960 2576
rect 120908 2524 120960 2576
rect 32588 2456 32640 2508
rect 122288 2456 122340 2508
rect 35808 2388 35860 2440
rect 123668 2388 123720 2440
rect 92388 2320 92440 2372
rect 125048 2320 125100 2372
rect 72608 2252 72660 2304
rect 124956 2252 125008 2304
rect 85948 2184 86000 2236
rect 126244 2184 126296 2236
rect 19248 2116 19300 2168
rect 115388 2116 115440 2168
rect 168656 2116 168708 2168
rect 213276 2116 213328 2168
rect 25964 2048 26016 2100
rect 124312 2048 124364 2100
rect 183468 2048 183520 2100
rect 379980 2048 380032 2100
rect 506204 2048 506256 2100
rect 22652 1980 22704 2032
rect 118056 1980 118108 2032
rect 106004 1912 106056 1964
rect 115296 1912 115348 1964
rect 59268 1300 59320 1352
rect 183468 1300 183520 1352
<< metal2 >>
rect 386 163200 442 164000
rect 1214 163200 1270 164000
rect 2042 163200 2098 164000
rect 2962 163200 3018 164000
rect 3790 163200 3846 164000
rect 4710 163200 4766 164000
rect 5538 163200 5594 164000
rect 6366 163200 6422 164000
rect 7286 163200 7342 164000
rect 8114 163200 8170 164000
rect 9034 163200 9090 164000
rect 9862 163200 9918 164000
rect 10782 163200 10838 164000
rect 11610 163200 11666 164000
rect 12438 163200 12494 164000
rect 13358 163200 13414 164000
rect 13464 163254 13768 163282
rect 400 159458 428 163200
rect 1228 159526 1256 163200
rect 1216 159520 1268 159526
rect 1216 159462 1268 159468
rect 388 159452 440 159458
rect 388 159394 440 159400
rect 2056 156670 2084 163200
rect 2044 156664 2096 156670
rect 2044 156606 2096 156612
rect 2976 152522 3004 163200
rect 3804 159390 3832 163200
rect 4724 160750 4752 163200
rect 4712 160744 4764 160750
rect 4712 160686 4764 160692
rect 5552 159594 5580 163200
rect 5540 159588 5592 159594
rect 5540 159530 5592 159536
rect 3792 159384 3844 159390
rect 3792 159326 3844 159332
rect 6380 156738 6408 163200
rect 7300 158030 7328 163200
rect 8128 160721 8156 163200
rect 8114 160712 8170 160721
rect 8114 160647 8170 160656
rect 7288 158024 7340 158030
rect 7288 157966 7340 157972
rect 6368 156732 6420 156738
rect 6368 156674 6420 156680
rect 9048 155281 9076 163200
rect 9034 155272 9090 155281
rect 9034 155207 9090 155216
rect 9876 153882 9904 163200
rect 10796 158098 10824 163200
rect 11624 160818 11652 163200
rect 11612 160812 11664 160818
rect 11612 160754 11664 160760
rect 12452 159186 12480 163200
rect 13372 163146 13400 163200
rect 13464 163146 13492 163254
rect 13372 163118 13492 163146
rect 12440 159180 12492 159186
rect 12440 159122 12492 159128
rect 10784 158092 10836 158098
rect 10784 158034 10836 158040
rect 13740 153950 13768 163254
rect 14186 163200 14242 164000
rect 15106 163200 15162 164000
rect 15934 163200 15990 164000
rect 16854 163200 16910 164000
rect 17682 163200 17738 164000
rect 18510 163200 18566 164000
rect 19430 163200 19486 164000
rect 20258 163200 20314 164000
rect 20364 163254 20668 163282
rect 14200 161498 14228 163200
rect 14188 161492 14240 161498
rect 14188 161434 14240 161440
rect 13820 159180 13872 159186
rect 13820 159122 13872 159128
rect 13832 155242 13860 159122
rect 15120 158166 15148 163200
rect 15108 158160 15160 158166
rect 15108 158102 15160 158108
rect 15948 155417 15976 163200
rect 15934 155408 15990 155417
rect 15934 155343 15990 155352
rect 13820 155236 13872 155242
rect 13820 155178 13872 155184
rect 16868 154018 16896 163200
rect 17696 161566 17724 163200
rect 17684 161560 17736 161566
rect 17684 161502 17736 161508
rect 18524 160886 18552 163200
rect 18512 160880 18564 160886
rect 18512 160822 18564 160828
rect 19444 159798 19472 163200
rect 20272 163146 20300 163200
rect 20364 163146 20392 163254
rect 20272 163118 20392 163146
rect 19432 159792 19484 159798
rect 19432 159734 19484 159740
rect 20640 154086 20668 163254
rect 21178 163200 21234 164000
rect 22006 163200 22062 164000
rect 22834 163200 22890 164000
rect 23754 163200 23810 164000
rect 24582 163200 24638 164000
rect 25502 163200 25558 164000
rect 26330 163200 26386 164000
rect 27250 163200 27306 164000
rect 27356 163254 27568 163282
rect 21192 161634 21220 163200
rect 21180 161628 21232 161634
rect 21180 161570 21232 161576
rect 22020 159662 22048 163200
rect 22008 159656 22060 159662
rect 22008 159598 22060 159604
rect 22848 156806 22876 163200
rect 22836 156800 22888 156806
rect 22836 156742 22888 156748
rect 23768 154154 23796 163200
rect 24596 161702 24624 163200
rect 24584 161696 24636 161702
rect 24584 161638 24636 161644
rect 25516 155310 25544 163200
rect 26344 160954 26372 163200
rect 27264 163146 27292 163200
rect 27356 163146 27384 163254
rect 27264 163118 27384 163146
rect 26332 160948 26384 160954
rect 26332 160890 26384 160896
rect 25504 155304 25556 155310
rect 25504 155246 25556 155252
rect 27540 154222 27568 163254
rect 28078 163200 28134 164000
rect 28906 163200 28962 164000
rect 29826 163200 29882 164000
rect 30654 163200 30710 164000
rect 31574 163200 31630 164000
rect 32402 163200 32458 164000
rect 33322 163200 33378 164000
rect 34150 163200 34206 164000
rect 34256 163254 34468 163282
rect 28092 161770 28120 163200
rect 28080 161764 28132 161770
rect 28080 161706 28132 161712
rect 28920 160138 28948 163200
rect 28908 160132 28960 160138
rect 28908 160074 28960 160080
rect 28908 159588 28960 159594
rect 28908 159530 28960 159536
rect 28920 157146 28948 159530
rect 28908 157140 28960 157146
rect 28908 157082 28960 157088
rect 29840 155378 29868 163200
rect 29828 155372 29880 155378
rect 29828 155314 29880 155320
rect 30668 154290 30696 163200
rect 31588 161838 31616 163200
rect 31576 161832 31628 161838
rect 31576 161774 31628 161780
rect 32416 159730 32444 163200
rect 33336 159866 33364 163200
rect 34164 163146 34192 163200
rect 34256 163146 34284 163254
rect 34164 163118 34284 163146
rect 33324 159860 33376 159866
rect 33324 159802 33376 159808
rect 32404 159724 32456 159730
rect 32404 159666 32456 159672
rect 34440 154358 34468 163254
rect 34978 163200 35034 164000
rect 35898 163200 35954 164000
rect 35992 163532 36044 163538
rect 35992 163474 36044 163480
rect 34992 159594 35020 163200
rect 35912 163146 35940 163200
rect 36004 163146 36032 163474
rect 36726 163200 36782 164000
rect 37646 163200 37702 164000
rect 38474 163200 38530 164000
rect 39302 163200 39358 164000
rect 39396 163464 39448 163470
rect 39396 163406 39448 163412
rect 35912 163118 36032 163146
rect 34980 159588 35032 159594
rect 34980 159530 35032 159536
rect 34520 159384 34572 159390
rect 34520 159326 34572 159332
rect 34532 158642 34560 159326
rect 34520 158636 34572 158642
rect 34520 158578 34572 158584
rect 36740 156641 36768 163200
rect 37660 161022 37688 163200
rect 37648 161016 37700 161022
rect 37648 160958 37700 160964
rect 38488 159390 38516 163200
rect 39316 163146 39344 163200
rect 39408 163146 39436 163406
rect 40222 163200 40278 164000
rect 41050 163200 41106 164000
rect 41970 163200 42026 164000
rect 42798 163200 42854 164000
rect 42892 163668 42944 163674
rect 42892 163610 42944 163616
rect 39316 163118 39436 163146
rect 39948 159452 40000 159458
rect 39948 159394 40000 159400
rect 38476 159384 38528 159390
rect 38476 159326 38528 159332
rect 39960 157962 39988 159394
rect 39948 157956 40000 157962
rect 39948 157898 40000 157904
rect 40236 156777 40264 163200
rect 41064 159934 41092 163200
rect 41052 159928 41104 159934
rect 41052 159870 41104 159876
rect 41420 159792 41472 159798
rect 41420 159734 41472 159740
rect 40222 156768 40278 156777
rect 40222 156703 40278 156712
rect 36726 156632 36782 156641
rect 36726 156567 36782 156576
rect 41432 155786 41460 159734
rect 41984 158778 42012 163200
rect 42812 163146 42840 163200
rect 42904 163146 42932 163610
rect 43718 163200 43774 164000
rect 44546 163200 44602 164000
rect 45374 163200 45430 164000
rect 46294 163200 46350 164000
rect 46388 163600 46440 163606
rect 46388 163542 46440 163548
rect 42812 163118 42932 163146
rect 41972 158772 42024 158778
rect 41972 158714 42024 158720
rect 43732 156913 43760 163200
rect 43718 156904 43774 156913
rect 43718 156839 43774 156848
rect 41420 155780 41472 155786
rect 41420 155722 41472 155728
rect 44560 155446 44588 163200
rect 45388 159458 45416 163200
rect 46308 163146 46336 163200
rect 46400 163146 46428 163542
rect 47122 163200 47178 164000
rect 48042 163200 48098 164000
rect 48870 163200 48926 164000
rect 49790 163200 49846 164000
rect 49884 163736 49936 163742
rect 49884 163678 49936 163684
rect 46308 163118 46428 163146
rect 47136 159798 47164 163200
rect 47124 159792 47176 159798
rect 47124 159734 47176 159740
rect 45376 159452 45428 159458
rect 45376 159394 45428 159400
rect 48056 159322 48084 163200
rect 48044 159316 48096 159322
rect 48044 159258 48096 159264
rect 48884 158817 48912 163200
rect 49804 163146 49832 163200
rect 49896 163146 49924 163678
rect 50618 163200 50674 164000
rect 51446 163200 51502 164000
rect 52366 163200 52422 164000
rect 53194 163200 53250 164000
rect 53288 163804 53340 163810
rect 53288 163746 53340 163752
rect 49804 163118 49924 163146
rect 50632 160206 50660 163200
rect 50620 160200 50672 160206
rect 50620 160142 50672 160148
rect 49608 159860 49660 159866
rect 49608 159802 49660 159808
rect 48870 158808 48926 158817
rect 46388 158772 46440 158778
rect 48870 158743 48926 158752
rect 46388 158714 46440 158720
rect 46400 158001 46428 158714
rect 46386 157992 46442 158001
rect 46386 157927 46442 157936
rect 44548 155440 44600 155446
rect 44548 155382 44600 155388
rect 34428 154352 34480 154358
rect 34428 154294 34480 154300
rect 30656 154284 30708 154290
rect 30656 154226 30708 154232
rect 27528 154216 27580 154222
rect 27528 154158 27580 154164
rect 23756 154148 23808 154154
rect 23756 154090 23808 154096
rect 20628 154080 20680 154086
rect 20628 154022 20680 154028
rect 16856 154012 16908 154018
rect 16856 153954 16908 153960
rect 13728 153944 13780 153950
rect 13728 153886 13780 153892
rect 9864 153876 9916 153882
rect 9864 153818 9916 153824
rect 43812 153536 43864 153542
rect 43812 153478 43864 153484
rect 26606 153368 26662 153377
rect 26606 153303 26662 153312
rect 5998 153232 6054 153241
rect 5998 153167 6054 153176
rect 2964 152516 3016 152522
rect 2964 152458 3016 152464
rect 6012 151994 6040 153167
rect 16212 152312 16264 152318
rect 16212 152254 16264 152260
rect 16224 151994 16252 152254
rect 26620 151994 26648 153303
rect 39994 152108 40046 152114
rect 39994 152050 40046 152056
rect 36912 152040 36964 152046
rect 5704 151966 6040 151994
rect 16008 151966 16252 151994
rect 26312 151966 26648 151994
rect 29716 151978 30052 151994
rect 36616 151988 36912 151994
rect 36616 151982 36964 151988
rect 29716 151972 30064 151978
rect 29716 151966 30012 151972
rect 36616 151966 36952 151982
rect 40006 151980 40034 152050
rect 43824 151994 43852 153478
rect 46756 153332 46808 153338
rect 46756 153274 46808 153280
rect 43516 151966 43852 151994
rect 30012 151914 30064 151920
rect 19708 151904 19760 151910
rect 12806 151872 12862 151881
rect 12512 151830 12806 151858
rect 19412 151852 19708 151858
rect 19412 151846 19760 151852
rect 46768 151858 46796 153274
rect 49620 152425 49648 159802
rect 51460 158302 51488 163200
rect 52380 159882 52408 163200
rect 53208 163146 53236 163200
rect 53300 163146 53328 163746
rect 54114 163200 54170 164000
rect 54942 163200 54998 164000
rect 55862 163200 55918 164000
rect 56690 163200 56746 164000
rect 56784 163872 56836 163878
rect 56784 163814 56836 163820
rect 53208 163118 53328 163146
rect 52380 159854 52500 159882
rect 51448 158296 51500 158302
rect 51448 158238 51500 158244
rect 52472 158234 52500 159854
rect 52460 158228 52512 158234
rect 52460 158170 52512 158176
rect 54128 157185 54156 163200
rect 54114 157176 54170 157185
rect 54114 157111 54170 157120
rect 54956 157049 54984 163200
rect 55876 159361 55904 163200
rect 56704 163146 56732 163200
rect 56796 163146 56824 163814
rect 57518 163200 57574 164000
rect 58438 163200 58494 164000
rect 59266 163200 59322 164000
rect 60186 163200 60242 164000
rect 60464 163940 60516 163946
rect 60464 163882 60516 163888
rect 60476 163282 60504 163882
rect 60292 163254 60504 163282
rect 56704 163118 56824 163146
rect 56508 159928 56560 159934
rect 56508 159870 56560 159876
rect 55862 159352 55918 159361
rect 55862 159287 55918 159296
rect 54942 157040 54998 157049
rect 54942 156975 54998 156984
rect 50620 153400 50672 153406
rect 50620 153342 50672 153348
rect 49606 152416 49662 152425
rect 49606 152351 49662 152360
rect 50632 151994 50660 153342
rect 56520 152697 56548 159870
rect 57532 155514 57560 163200
rect 58452 162450 58480 163200
rect 58440 162444 58492 162450
rect 58440 162386 58492 162392
rect 59280 159882 59308 163200
rect 60200 163146 60228 163200
rect 60292 163146 60320 163254
rect 61014 163200 61070 164000
rect 61842 163200 61898 164000
rect 62762 163200 62818 164000
rect 63590 163200 63646 164000
rect 63868 163940 63920 163946
rect 63868 163882 63920 163888
rect 63880 163282 63908 163882
rect 63696 163254 63908 163282
rect 60200 163118 60320 163146
rect 59280 159854 59400 159882
rect 59372 158370 59400 159854
rect 59360 158364 59412 158370
rect 59360 158306 59412 158312
rect 61028 156874 61056 163200
rect 61856 160002 61884 163200
rect 61844 159996 61896 160002
rect 61844 159938 61896 159944
rect 62120 159656 62172 159662
rect 62776 159633 62804 163200
rect 63604 163146 63632 163200
rect 63696 163146 63724 163254
rect 64510 163200 64566 164000
rect 65338 163200 65394 164000
rect 66258 163200 66314 164000
rect 67086 163200 67142 164000
rect 67914 163200 67970 164000
rect 68834 163200 68890 164000
rect 69662 163200 69718 164000
rect 70582 163200 70638 164000
rect 71410 163200 71466 164000
rect 72330 163200 72386 164000
rect 73158 163200 73214 164000
rect 73986 163200 74042 164000
rect 74906 163200 74962 164000
rect 75734 163200 75790 164000
rect 76654 163200 76710 164000
rect 77482 163200 77538 164000
rect 78310 163200 78366 164000
rect 79230 163200 79286 164000
rect 80058 163200 80114 164000
rect 80978 163200 81034 164000
rect 81806 163200 81862 164000
rect 82726 163200 82782 164000
rect 83554 163200 83610 164000
rect 84382 163200 84438 164000
rect 85302 163200 85358 164000
rect 86130 163200 86186 164000
rect 87050 163200 87106 164000
rect 87878 163200 87934 164000
rect 88798 163200 88854 164000
rect 89626 163200 89682 164000
rect 90454 163200 90510 164000
rect 91374 163200 91430 164000
rect 92202 163200 92258 164000
rect 93122 163200 93178 164000
rect 93950 163200 94006 164000
rect 94870 163200 94926 164000
rect 95698 163200 95754 164000
rect 96526 163200 96582 164000
rect 97446 163200 97502 164000
rect 98274 163200 98330 164000
rect 99194 163200 99250 164000
rect 100022 163200 100078 164000
rect 100850 163200 100906 164000
rect 101770 163200 101826 164000
rect 102598 163200 102654 164000
rect 103518 163200 103574 164000
rect 104346 163200 104402 164000
rect 105266 163200 105322 164000
rect 106094 163200 106150 164000
rect 106922 163200 106978 164000
rect 107842 163200 107898 164000
rect 108670 163200 108726 164000
rect 109590 163200 109646 164000
rect 110418 163200 110474 164000
rect 110512 163260 110564 163266
rect 110512 163202 110564 163208
rect 63604 163118 63724 163146
rect 62120 159598 62172 159604
rect 62762 159624 62818 159633
rect 61016 156868 61068 156874
rect 61016 156810 61068 156816
rect 57520 155508 57572 155514
rect 57520 155450 57572 155456
rect 62132 153066 62160 159598
rect 62762 159559 62818 159568
rect 64524 155553 64552 163200
rect 65352 155689 65380 163200
rect 66272 161090 66300 163200
rect 67100 162518 67128 163200
rect 67088 162512 67140 162518
rect 67088 162454 67140 162460
rect 66260 161084 66312 161090
rect 66260 161026 66312 161032
rect 65338 155680 65394 155689
rect 65338 155615 65394 155624
rect 67928 155582 67956 163200
rect 68848 159497 68876 163200
rect 69676 160993 69704 163200
rect 70596 162654 70624 163200
rect 70584 162648 70636 162654
rect 70584 162590 70636 162596
rect 69662 160984 69718 160993
rect 69662 160919 69718 160928
rect 71424 159866 71452 163200
rect 72344 160857 72372 163200
rect 72330 160848 72386 160857
rect 72330 160783 72386 160792
rect 71412 159860 71464 159866
rect 71412 159802 71464 159808
rect 73172 159769 73200 163200
rect 74000 162722 74028 163200
rect 73988 162716 74040 162722
rect 73988 162658 74040 162664
rect 73158 159760 73214 159769
rect 69664 159724 69716 159730
rect 73158 159695 73214 159704
rect 69664 159666 69716 159672
rect 68834 159488 68890 159497
rect 68834 159423 68890 159432
rect 67916 155576 67968 155582
rect 64510 155544 64566 155553
rect 67916 155518 67968 155524
rect 64510 155479 64566 155488
rect 69676 153105 69704 159666
rect 74920 157010 74948 163200
rect 75748 160041 75776 163200
rect 75734 160032 75790 160041
rect 75734 159967 75790 159976
rect 76668 158438 76696 163200
rect 77496 162858 77524 163200
rect 77484 162852 77536 162858
rect 77484 162794 77536 162800
rect 76656 158432 76708 158438
rect 76656 158374 76708 158380
rect 74908 157004 74960 157010
rect 74908 156946 74960 156952
rect 78324 156942 78352 163200
rect 79244 162790 79272 163200
rect 79232 162784 79284 162790
rect 79232 162726 79284 162732
rect 80072 161158 80100 163200
rect 80992 162926 81020 163200
rect 80980 162920 81032 162926
rect 80980 162862 81032 162868
rect 80060 161152 80112 161158
rect 80060 161094 80112 161100
rect 80060 159588 80112 159594
rect 80060 159530 80112 159536
rect 80072 157894 80100 159530
rect 80060 157888 80112 157894
rect 80060 157830 80112 157836
rect 81820 157078 81848 163200
rect 82740 159730 82768 163200
rect 83568 161129 83596 163200
rect 84396 163062 84424 163200
rect 84384 163056 84436 163062
rect 84384 162998 84436 163004
rect 83554 161120 83610 161129
rect 83554 161055 83610 161064
rect 82728 159724 82780 159730
rect 82728 159666 82780 159672
rect 81808 157072 81860 157078
rect 81808 157014 81860 157020
rect 78312 156936 78364 156942
rect 78312 156878 78364 156884
rect 85316 155650 85344 163200
rect 86144 158137 86172 163200
rect 86130 158128 86186 158137
rect 86130 158063 86186 158072
rect 85304 155644 85356 155650
rect 85304 155586 85356 155592
rect 69662 153096 69718 153105
rect 62120 153060 62172 153066
rect 69662 153031 69718 153040
rect 62120 153002 62172 153008
rect 56506 152688 56562 152697
rect 56506 152623 56562 152632
rect 87064 152590 87092 163200
rect 87892 163130 87920 163200
rect 87880 163124 87932 163130
rect 87880 163066 87932 163072
rect 88812 162994 88840 163200
rect 88800 162988 88852 162994
rect 88800 162930 88852 162936
rect 89640 159934 89668 163200
rect 90468 161226 90496 163200
rect 90456 161220 90508 161226
rect 90456 161162 90508 161168
rect 89628 159928 89680 159934
rect 89628 159870 89680 159876
rect 91388 159526 91416 163200
rect 89720 159520 89772 159526
rect 89720 159462 89772 159468
rect 91376 159520 91428 159526
rect 91376 159462 91428 159468
rect 89732 157865 89760 159462
rect 89718 157856 89774 157865
rect 89718 157791 89774 157800
rect 92216 155718 92244 163200
rect 92204 155712 92256 155718
rect 92204 155654 92256 155660
rect 87052 152584 87104 152590
rect 93136 152561 93164 163200
rect 93964 152658 93992 163200
rect 94884 158846 94912 163200
rect 94872 158840 94924 158846
rect 94872 158782 94924 158788
rect 95712 155825 95740 163200
rect 96540 159905 96568 163200
rect 97460 161265 97488 163200
rect 98288 163146 98316 163200
rect 98368 163192 98420 163198
rect 98288 163140 98368 163146
rect 98288 163134 98420 163140
rect 98288 163118 98408 163134
rect 97446 161256 97502 161265
rect 97446 161191 97502 161200
rect 96526 159896 96582 159905
rect 96526 159831 96582 159840
rect 99208 159254 99236 163200
rect 99380 159520 99432 159526
rect 99380 159462 99432 159468
rect 99196 159248 99248 159254
rect 99196 159190 99248 159196
rect 97816 158840 97868 158846
rect 97816 158782 97868 158788
rect 97828 155961 97856 158782
rect 99392 156602 99420 159462
rect 100036 159225 100064 163200
rect 100760 159792 100812 159798
rect 100760 159734 100812 159740
rect 100022 159216 100078 159225
rect 100022 159151 100078 159160
rect 100772 158681 100800 159734
rect 100864 159594 100892 163200
rect 100944 160268 100996 160274
rect 100944 160210 100996 160216
rect 100852 159588 100904 159594
rect 100852 159530 100904 159536
rect 100956 159322 100984 160210
rect 101784 159662 101812 163200
rect 101772 159656 101824 159662
rect 101772 159598 101824 159604
rect 100944 159316 100996 159322
rect 100944 159258 100996 159264
rect 100758 158672 100814 158681
rect 100758 158607 100814 158616
rect 102612 158506 102640 163200
rect 102600 158500 102652 158506
rect 102600 158442 102652 158448
rect 103532 157282 103560 163200
rect 104360 159526 104388 163200
rect 105280 161294 105308 163200
rect 105268 161288 105320 161294
rect 105268 161230 105320 161236
rect 104348 159520 104400 159526
rect 104348 159462 104400 159468
rect 103520 157276 103572 157282
rect 103520 157218 103572 157224
rect 106108 157214 106136 163200
rect 106936 159322 106964 163200
rect 106924 159316 106976 159322
rect 106924 159258 106976 159264
rect 107856 158273 107884 163200
rect 107842 158264 107898 158273
rect 107842 158199 107898 158208
rect 108684 157350 108712 163200
rect 108672 157344 108724 157350
rect 109604 157321 109632 163200
rect 110432 163146 110460 163200
rect 110524 163146 110552 163202
rect 111338 163200 111394 164000
rect 111444 163254 111748 163282
rect 110432 163118 110552 163146
rect 111352 163146 111380 163200
rect 111444 163146 111472 163254
rect 111352 163118 111472 163146
rect 108672 157286 108724 157292
rect 109590 157312 109646 157321
rect 109590 157247 109646 157256
rect 106096 157208 106148 157214
rect 106096 157150 106148 157156
rect 99380 156596 99432 156602
rect 99380 156538 99432 156544
rect 97814 155952 97870 155961
rect 97814 155887 97870 155896
rect 95698 155816 95754 155825
rect 95698 155751 95754 155760
rect 95148 153468 95200 153474
rect 95148 153410 95200 153416
rect 93952 152652 94004 152658
rect 93952 152594 94004 152600
rect 87052 152526 87104 152532
rect 93122 152552 93178 152561
rect 93122 152487 93178 152496
rect 91606 152176 91658 152182
rect 91606 152118 91658 152124
rect 50324 151966 50660 151994
rect 91618 151980 91646 152118
rect 95160 151994 95188 153410
rect 108948 153264 109000 153270
rect 108948 153206 109000 153212
rect 101910 152244 101962 152250
rect 101910 152186 101962 152192
rect 95036 151966 95188 151994
rect 101922 151980 101950 152186
rect 108960 151994 108988 153206
rect 111720 152726 111748 163254
rect 112166 163200 112222 164000
rect 112260 163328 112312 163334
rect 112260 163270 112312 163276
rect 112180 163146 112208 163200
rect 112272 163146 112300 163270
rect 112994 163200 113050 164000
rect 113914 163200 113970 164000
rect 114742 163200 114798 164000
rect 114836 163396 114888 163402
rect 114836 163338 114888 163344
rect 112180 163118 112300 163146
rect 113008 158409 113036 163200
rect 113928 159798 113956 163200
rect 114756 163146 114784 163200
rect 114848 163146 114876 163338
rect 115662 163200 115718 164000
rect 116490 163200 116546 164000
rect 117318 163200 117374 164000
rect 118238 163200 118294 164000
rect 118344 163254 118648 163282
rect 114756 163118 114876 163146
rect 114652 159860 114704 159866
rect 114652 159802 114704 159808
rect 113916 159792 113968 159798
rect 113916 159734 113968 159740
rect 112994 158400 113050 158409
rect 112994 158335 113050 158344
rect 114664 153202 114692 159802
rect 115676 155145 115704 163200
rect 115662 155136 115718 155145
rect 115662 155071 115718 155080
rect 116504 155038 116532 163200
rect 117332 161401 117360 163200
rect 118252 163146 118280 163200
rect 118344 163146 118372 163254
rect 118252 163118 118372 163146
rect 117318 161392 117374 161401
rect 117318 161327 117374 161336
rect 116492 155032 116544 155038
rect 116492 154974 116544 154980
rect 118056 153536 118108 153542
rect 118056 153478 118108 153484
rect 115296 153400 115348 153406
rect 115296 153342 115348 153348
rect 117962 153368 118018 153377
rect 114652 153196 114704 153202
rect 114652 153138 114704 153144
rect 111708 152720 111760 152726
rect 111708 152662 111760 152668
rect 115204 152108 115256 152114
rect 115204 152050 115256 152056
rect 108836 151966 108988 151994
rect 19412 151830 19748 151846
rect 46768 151830 46920 151858
rect 105340 151842 105676 151858
rect 105340 151836 105688 151842
rect 105340 151830 105636 151836
rect 12806 151807 12862 151816
rect 105636 151778 105688 151784
rect 114560 151836 114612 151842
rect 114560 151778 114612 151784
rect 60720 151434 60872 151450
rect 64124 151434 64460 151450
rect 60720 151428 60884 151434
rect 60720 151422 60832 151428
rect 64124 151428 64472 151434
rect 64124 151422 64420 151428
rect 60832 151370 60884 151376
rect 64420 151370 64472 151376
rect 53932 151360 53984 151366
rect 9402 151328 9458 151337
rect 9108 151286 9402 151314
rect 23110 151328 23166 151337
rect 22816 151286 23110 151314
rect 9402 151263 9458 151272
rect 33506 151328 33562 151337
rect 33212 151286 33506 151314
rect 23110 151263 23166 151272
rect 53820 151308 53932 151314
rect 57520 151360 57572 151366
rect 53820 151302 53984 151308
rect 57224 151308 57520 151314
rect 67640 151360 67692 151366
rect 57224 151302 57572 151308
rect 67528 151308 67640 151314
rect 71320 151360 71372 151366
rect 67528 151302 67692 151308
rect 71024 151308 71320 151314
rect 74540 151360 74592 151366
rect 71024 151302 71372 151308
rect 74428 151308 74540 151314
rect 78128 151360 78180 151366
rect 74428 151302 74592 151308
rect 77832 151308 78128 151314
rect 81440 151360 81492 151366
rect 77832 151302 78180 151308
rect 81328 151308 81440 151314
rect 85028 151360 85080 151366
rect 81328 151302 81492 151308
rect 84732 151308 85028 151314
rect 88340 151360 88392 151366
rect 84732 151302 85080 151308
rect 88228 151308 88340 151314
rect 98828 151360 98880 151366
rect 88228 151302 88392 151308
rect 98532 151308 98828 151314
rect 98532 151302 98880 151308
rect 53820 151286 53972 151302
rect 57224 151286 57560 151302
rect 67528 151286 67680 151302
rect 71024 151286 71360 151302
rect 74428 151286 74580 151302
rect 77832 151286 78168 151302
rect 81328 151286 81480 151302
rect 84732 151286 85068 151302
rect 88228 151286 88380 151302
rect 98532 151286 98868 151302
rect 112240 151286 112576 151314
rect 33506 151263 33562 151272
rect 112548 150686 112576 151286
rect 112536 150680 112588 150686
rect 112536 150622 112588 150628
rect 114572 147626 114600 151778
rect 114560 147620 114612 147626
rect 114560 147562 114612 147568
rect 115216 111790 115244 152050
rect 115308 117298 115336 153342
rect 117228 153332 117280 153338
rect 117962 153303 118018 153312
rect 117228 153274 117280 153280
rect 116584 152176 116636 152182
rect 116584 152118 116636 152124
rect 115388 151156 115440 151162
rect 115388 151098 115440 151104
rect 115400 137970 115428 151098
rect 116596 140758 116624 152118
rect 116860 151292 116912 151298
rect 116860 151234 116912 151240
rect 116768 150884 116820 150890
rect 116768 150826 116820 150832
rect 116674 146160 116730 146169
rect 116674 146095 116730 146104
rect 116688 145246 116716 146095
rect 116676 145240 116728 145246
rect 116676 145182 116728 145188
rect 116780 145058 116808 150826
rect 116688 145030 116808 145058
rect 116584 140752 116636 140758
rect 116584 140694 116636 140700
rect 115388 137964 115440 137970
rect 115388 137906 115440 137912
rect 116582 134736 116638 134745
rect 116582 134671 116638 134680
rect 115296 117292 115348 117298
rect 115296 117234 115348 117240
rect 115204 111784 115256 111790
rect 115204 111726 115256 111732
rect 115938 89176 115994 89185
rect 115938 89111 115994 89120
rect 115952 88602 115980 89111
rect 115940 88596 115992 88602
rect 115940 88538 115992 88544
rect 116596 88330 116624 134671
rect 116688 131102 116716 145030
rect 116872 142154 116900 151234
rect 117240 149734 117268 153274
rect 117228 149728 117280 149734
rect 117228 149670 117280 149676
rect 116780 142126 116900 142154
rect 116676 131096 116728 131102
rect 116676 131038 116728 131044
rect 116674 123312 116730 123321
rect 116674 123247 116730 123256
rect 116584 88324 116636 88330
rect 116584 88266 116636 88272
rect 116688 86970 116716 123247
rect 116780 121446 116808 142126
rect 116768 121440 116820 121446
rect 116768 121382 116820 121388
rect 116766 112024 116822 112033
rect 116766 111959 116822 111968
rect 116676 86964 116728 86970
rect 116676 86906 116728 86912
rect 116780 84182 116808 111959
rect 117976 103494 118004 153303
rect 118068 113150 118096 153478
rect 118620 152794 118648 163254
rect 119066 163200 119122 164000
rect 119986 163200 120042 164000
rect 120814 163200 120870 164000
rect 121734 163200 121790 164000
rect 122562 163200 122618 164000
rect 123390 163200 123446 164000
rect 124310 163200 124366 164000
rect 125138 163200 125194 164000
rect 125244 163254 125548 163282
rect 118700 159996 118752 160002
rect 118700 159938 118752 159944
rect 118712 153134 118740 159938
rect 119080 159866 119108 163200
rect 119068 159860 119120 159866
rect 119068 159802 119120 159808
rect 120000 158574 120028 163200
rect 119988 158568 120040 158574
rect 119988 158510 120040 158516
rect 120828 155922 120856 163200
rect 121748 161362 121776 163200
rect 121736 161356 121788 161362
rect 121736 161298 121788 161304
rect 120816 155916 120868 155922
rect 120816 155858 120868 155864
rect 122576 155854 122604 163200
rect 123404 156534 123432 163200
rect 124324 161974 124352 163200
rect 125152 163146 125180 163200
rect 125244 163146 125272 163254
rect 125152 163118 125272 163146
rect 124312 161968 124364 161974
rect 124312 161910 124364 161916
rect 123392 156528 123444 156534
rect 123392 156470 123444 156476
rect 122564 155848 122616 155854
rect 122564 155790 122616 155796
rect 119896 153264 119948 153270
rect 119896 153206 119948 153212
rect 120722 153232 120778 153241
rect 118700 153128 118752 153134
rect 118700 153070 118752 153076
rect 118608 152788 118660 152794
rect 118608 152730 118660 152736
rect 118608 152244 118660 152250
rect 118608 152186 118660 152192
rect 118148 150816 118200 150822
rect 118148 150758 118200 150764
rect 118160 128314 118188 150758
rect 118620 146266 118648 152186
rect 119342 151872 119398 151881
rect 119342 151807 119398 151816
rect 118608 146260 118660 146266
rect 118608 146202 118660 146208
rect 118148 128308 118200 128314
rect 118148 128250 118200 128256
rect 118056 113144 118108 113150
rect 118056 113086 118108 113092
rect 117964 103488 118016 103494
rect 117964 103430 118016 103436
rect 116950 100600 117006 100609
rect 116950 100535 117006 100544
rect 116964 99482 116992 100535
rect 116952 99476 117004 99482
rect 116952 99418 117004 99424
rect 119356 96626 119384 151807
rect 119528 150952 119580 150958
rect 119528 150894 119580 150900
rect 119434 150784 119490 150793
rect 119434 150719 119490 150728
rect 119448 107642 119476 150719
rect 119540 132462 119568 150894
rect 119908 149054 119936 153206
rect 120722 153167 120778 153176
rect 120736 151162 120764 153167
rect 125520 152862 125548 163254
rect 126058 163200 126114 164000
rect 126886 163200 126942 164000
rect 127806 163200 127862 164000
rect 128634 163200 128690 164000
rect 129462 163200 129518 164000
rect 130382 163200 130438 164000
rect 131210 163200 131266 164000
rect 132130 163200 132186 164000
rect 132236 163254 132448 163282
rect 126072 161906 126100 163200
rect 126060 161900 126112 161906
rect 126060 161842 126112 161848
rect 126900 158545 126928 163200
rect 127820 158710 127848 163200
rect 127808 158704 127860 158710
rect 127808 158646 127860 158652
rect 126886 158536 126942 158545
rect 126886 158471 126942 158480
rect 126704 153468 126756 153474
rect 126704 153410 126756 153416
rect 125508 152856 125560 152862
rect 125508 152798 125560 152804
rect 124864 152312 124916 152318
rect 124864 152254 124916 152260
rect 120816 152040 120868 152046
rect 120816 151982 120868 151988
rect 120724 151156 120776 151162
rect 120724 151098 120776 151104
rect 119896 149048 119948 149054
rect 119896 148990 119948 148996
rect 120724 145240 120776 145246
rect 120724 145182 120776 145188
rect 119528 132456 119580 132462
rect 119528 132398 119580 132404
rect 119436 107636 119488 107642
rect 119436 107578 119488 107584
rect 119344 96620 119396 96626
rect 119344 96562 119396 96568
rect 120736 89690 120764 145182
rect 120828 109002 120856 151982
rect 122196 151972 122248 151978
rect 122196 151914 122248 151920
rect 120908 150748 120960 150754
rect 120908 150690 120960 150696
rect 120920 126954 120948 150690
rect 122102 150648 122158 150657
rect 122102 150583 122158 150592
rect 120908 126948 120960 126954
rect 120908 126890 120960 126896
rect 120816 108996 120868 109002
rect 120816 108938 120868 108944
rect 122116 102134 122144 150583
rect 122208 104854 122236 151914
rect 123484 151904 123536 151910
rect 123484 151846 123536 151852
rect 122288 151020 122340 151026
rect 122288 150962 122340 150968
rect 122300 133890 122328 150962
rect 122288 133884 122340 133890
rect 122288 133826 122340 133832
rect 122196 104848 122248 104854
rect 122196 104790 122248 104796
rect 122104 102128 122156 102134
rect 122104 102070 122156 102076
rect 122104 99476 122156 99482
rect 122104 99418 122156 99424
rect 120724 89684 120776 89690
rect 120724 89626 120776 89632
rect 117964 88596 118016 88602
rect 117964 88538 118016 88544
rect 116768 84176 116820 84182
rect 116768 84118 116820 84124
rect 117976 80034 118004 88538
rect 122116 82822 122144 99418
rect 123496 99346 123524 151846
rect 123576 151224 123628 151230
rect 123576 151166 123628 151172
rect 123588 118658 123616 151166
rect 123668 151088 123720 151094
rect 123668 151030 123720 151036
rect 123680 136610 123708 151030
rect 124588 150476 124640 150482
rect 124588 150418 124640 150424
rect 124600 143546 124628 150418
rect 124588 143540 124640 143546
rect 124588 143482 124640 143488
rect 123668 136604 123720 136610
rect 123668 136546 123720 136552
rect 123576 118652 123628 118658
rect 123576 118594 123628 118600
rect 123484 99340 123536 99346
rect 123484 99282 123536 99288
rect 124876 97986 124904 152254
rect 126336 150612 126388 150618
rect 126336 150554 126388 150560
rect 124956 150544 125008 150550
rect 124956 150486 125008 150492
rect 126242 150512 126298 150521
rect 124968 122466 124996 150486
rect 126242 150447 126298 150456
rect 124956 122460 125008 122466
rect 124956 122402 125008 122408
rect 124864 97980 124916 97986
rect 124864 97922 124916 97928
rect 126256 93265 126284 150447
rect 126348 124137 126376 150554
rect 126716 150482 126744 153410
rect 128648 152969 128676 163200
rect 129476 155174 129504 163200
rect 130396 157962 130424 163200
rect 131224 160002 131252 163200
rect 132144 163146 132172 163200
rect 132236 163146 132264 163254
rect 132144 163118 132264 163146
rect 131212 159996 131264 160002
rect 131212 159938 131264 159944
rect 130292 157956 130344 157962
rect 130292 157898 130344 157904
rect 130384 157956 130436 157962
rect 130384 157898 130436 157904
rect 129464 155168 129516 155174
rect 129464 155110 129516 155116
rect 128634 152960 128690 152969
rect 128634 152895 128690 152904
rect 130304 151980 130332 157898
rect 130842 157856 130898 157865
rect 130842 157791 130898 157800
rect 130856 151980 130884 157791
rect 131488 156664 131540 156670
rect 131488 156606 131540 156612
rect 131500 151980 131528 156606
rect 132420 152833 132448 163254
rect 132958 163200 133014 164000
rect 133878 163200 133934 164000
rect 134706 163200 134762 164000
rect 135534 163200 135590 164000
rect 136454 163200 136510 164000
rect 137282 163200 137338 164000
rect 138202 163200 138258 164000
rect 139030 163200 139086 164000
rect 139858 163200 139914 164000
rect 140778 163200 140834 164000
rect 141606 163200 141662 164000
rect 142526 163200 142582 164000
rect 143354 163200 143410 164000
rect 144274 163200 144330 164000
rect 145102 163200 145158 164000
rect 145930 163200 145986 164000
rect 146850 163200 146906 164000
rect 147678 163200 147734 164000
rect 148598 163200 148654 164000
rect 149426 163200 149482 164000
rect 150346 163200 150402 164000
rect 151174 163200 151230 164000
rect 152002 163200 152058 164000
rect 152922 163200 152978 164000
rect 153750 163200 153806 164000
rect 154670 163200 154726 164000
rect 155498 163200 155554 164000
rect 156236 163532 156288 163538
rect 156236 163474 156288 163480
rect 132776 158636 132828 158642
rect 132776 158578 132828 158584
rect 132406 152824 132462 152833
rect 132406 152759 132462 152768
rect 132132 152516 132184 152522
rect 132132 152458 132184 152464
rect 132144 151980 132172 152458
rect 132788 151980 132816 158578
rect 132972 152386 133000 163200
rect 133420 160744 133472 160750
rect 133420 160686 133472 160692
rect 132960 152380 133012 152386
rect 132960 152322 133012 152328
rect 133432 151980 133460 160686
rect 133892 158642 133920 163200
rect 134720 161474 134748 163200
rect 134720 161446 134840 161474
rect 133880 158636 133932 158642
rect 133880 158578 133932 158584
rect 134064 157140 134116 157146
rect 134064 157082 134116 157088
rect 134076 151980 134104 157082
rect 134708 156732 134760 156738
rect 134708 156674 134760 156680
rect 134720 151980 134748 156674
rect 134812 156505 134840 161446
rect 135352 158024 135404 158030
rect 135352 157966 135404 157972
rect 134798 156496 134854 156505
rect 134798 156431 134854 156440
rect 135364 151980 135392 157966
rect 135548 152318 135576 163200
rect 135994 160712 136050 160721
rect 135994 160647 136050 160656
rect 135536 152312 135588 152318
rect 135536 152254 135588 152260
rect 136008 151980 136036 160647
rect 136468 156670 136496 163200
rect 137296 157146 137324 163200
rect 138216 160070 138244 163200
rect 138572 160812 138624 160818
rect 138572 160754 138624 160760
rect 138204 160064 138256 160070
rect 138204 160006 138256 160012
rect 138020 159248 138072 159254
rect 138020 159190 138072 159196
rect 137928 158092 137980 158098
rect 137928 158034 137980 158040
rect 137284 157140 137336 157146
rect 137284 157082 137336 157088
rect 136456 156664 136508 156670
rect 136456 156606 136508 156612
rect 136638 155272 136694 155281
rect 136638 155207 136694 155216
rect 136652 151980 136680 155207
rect 137284 153876 137336 153882
rect 137284 153818 137336 153824
rect 137296 151980 137324 153818
rect 137940 151980 137968 158034
rect 138032 155281 138060 159190
rect 138018 155272 138074 155281
rect 138018 155207 138074 155216
rect 138584 151980 138612 160754
rect 139044 160750 139072 163200
rect 139872 162042 139900 163200
rect 139860 162036 139912 162042
rect 139860 161978 139912 161984
rect 140504 161492 140556 161498
rect 140504 161434 140556 161440
rect 139032 160744 139084 160750
rect 139032 160686 139084 160692
rect 139216 155236 139268 155242
rect 139216 155178 139268 155184
rect 139228 151980 139256 155178
rect 139860 153944 139912 153950
rect 139860 153886 139912 153892
rect 139872 151980 139900 153886
rect 140516 151980 140544 161434
rect 140792 158030 140820 163200
rect 141620 162110 141648 163200
rect 141608 162104 141660 162110
rect 141608 162046 141660 162052
rect 142436 161560 142488 161566
rect 142436 161502 142488 161508
rect 141148 158160 141200 158166
rect 141148 158102 141200 158108
rect 140780 158024 140832 158030
rect 140780 157966 140832 157972
rect 141160 151980 141188 158102
rect 142448 156618 142476 161502
rect 142540 158778 142568 163200
rect 142528 158772 142580 158778
rect 142528 158714 142580 158720
rect 143264 158772 143316 158778
rect 143264 158714 143316 158720
rect 142448 156590 143120 156618
rect 141790 155408 141846 155417
rect 141790 155343 141846 155352
rect 141804 151980 141832 155343
rect 142436 154012 142488 154018
rect 142436 153954 142488 153960
rect 142448 151980 142476 153954
rect 143092 151980 143120 156590
rect 143276 152998 143304 158714
rect 143368 156738 143396 163200
rect 143724 160880 143776 160886
rect 143724 160822 143776 160828
rect 143356 156732 143408 156738
rect 143356 156674 143408 156680
rect 143264 152992 143316 152998
rect 143264 152934 143316 152940
rect 143736 151980 143764 160822
rect 144288 158098 144316 163200
rect 144276 158092 144328 158098
rect 144276 158034 144328 158040
rect 144368 155780 144420 155786
rect 144368 155722 144420 155728
rect 144380 151980 144408 155722
rect 145116 155242 145144 163200
rect 145656 161628 145708 161634
rect 145656 161570 145708 161576
rect 145104 155236 145156 155242
rect 145104 155178 145156 155184
rect 145012 154080 145064 154086
rect 145012 154022 145064 154028
rect 145024 151980 145052 154022
rect 145668 151980 145696 161570
rect 145944 160818 145972 163200
rect 146864 161498 146892 163200
rect 146852 161492 146904 161498
rect 146852 161434 146904 161440
rect 145932 160812 145984 160818
rect 145932 160754 145984 160760
rect 147692 158166 147720 163200
rect 148232 161696 148284 161702
rect 148232 161638 148284 161644
rect 147680 158160 147732 158166
rect 147680 158102 147732 158108
rect 146944 156800 146996 156806
rect 146944 156742 146996 156748
rect 146300 153060 146352 153066
rect 146300 153002 146352 153008
rect 146312 151980 146340 153002
rect 146956 151980 146984 156742
rect 147588 154148 147640 154154
rect 147588 154090 147640 154096
rect 147600 151980 147628 154090
rect 148244 151980 148272 161638
rect 148612 159254 148640 163200
rect 149440 162246 149468 163200
rect 149428 162240 149480 162246
rect 149428 162182 149480 162188
rect 149520 160948 149572 160954
rect 149520 160890 149572 160896
rect 148600 159248 148652 159254
rect 148600 159190 148652 159196
rect 148876 155304 148928 155310
rect 148876 155246 148928 155252
rect 148888 151980 148916 155246
rect 149532 151980 149560 160890
rect 150360 155786 150388 163200
rect 150808 161764 150860 161770
rect 150808 161706 150860 161712
rect 150348 155780 150400 155786
rect 150348 155722 150400 155728
rect 150164 154216 150216 154222
rect 150164 154158 150216 154164
rect 150176 151980 150204 154158
rect 150820 151980 150848 161706
rect 151188 155310 151216 163200
rect 151452 160132 151504 160138
rect 151452 160074 151504 160080
rect 151176 155304 151228 155310
rect 151176 155246 151228 155252
rect 151464 151980 151492 160074
rect 152016 152454 152044 163200
rect 152936 160886 152964 163200
rect 153764 162178 153792 163200
rect 153752 162172 153804 162178
rect 153752 162114 153804 162120
rect 153384 161832 153436 161838
rect 153384 161774 153436 161780
rect 152924 160880 152976 160886
rect 152924 160822 152976 160828
rect 152096 155372 152148 155378
rect 152096 155314 152148 155320
rect 152004 152448 152056 152454
rect 152004 152390 152056 152396
rect 152108 151980 152136 155314
rect 152740 154284 152792 154290
rect 152740 154226 152792 154232
rect 152752 151980 152780 154226
rect 153396 151980 153424 161774
rect 154396 159452 154448 159458
rect 154396 159394 154448 159400
rect 154408 153882 154436 159394
rect 154488 159384 154540 159390
rect 154488 159326 154540 159332
rect 154500 154154 154528 159326
rect 154684 156806 154712 163200
rect 155512 159390 155540 163200
rect 155500 159384 155552 159390
rect 155500 159326 155552 159332
rect 155960 157888 156012 157894
rect 155960 157830 156012 157836
rect 154672 156800 154724 156806
rect 154672 156742 154724 156748
rect 155316 154352 155368 154358
rect 155316 154294 155368 154300
rect 154488 154148 154540 154154
rect 154488 154090 154540 154096
rect 154396 153876 154448 153882
rect 154396 153818 154448 153824
rect 154026 153096 154082 153105
rect 154026 153031 154082 153040
rect 154040 151980 154068 153031
rect 154670 152416 154726 152425
rect 154670 152351 154726 152360
rect 154684 151980 154712 152351
rect 155328 151980 155356 154294
rect 155972 151980 156000 157830
rect 156248 156618 156276 163474
rect 156326 163200 156382 164000
rect 156432 163254 156736 163282
rect 156340 163146 156368 163200
rect 156432 163146 156460 163254
rect 156340 163118 156460 163146
rect 156248 156590 156644 156618
rect 156616 151980 156644 156590
rect 156708 152425 156736 163254
rect 157246 163200 157302 164000
rect 158074 163200 158130 164000
rect 158994 163200 159050 164000
rect 159180 163464 159232 163470
rect 159180 163406 159232 163412
rect 157260 161566 157288 163200
rect 157248 161560 157300 161566
rect 157248 161502 157300 161508
rect 157892 161016 157944 161022
rect 157892 160958 157944 160964
rect 157246 156632 157302 156641
rect 157246 156567 157302 156576
rect 156694 152416 156750 152425
rect 156694 152351 156750 152360
rect 157260 151980 157288 156567
rect 157904 151980 157932 160958
rect 158088 157894 158116 163200
rect 159008 161634 159036 163200
rect 158996 161628 159048 161634
rect 158996 161570 159048 161576
rect 158076 157888 158128 157894
rect 158076 157830 158128 157836
rect 158536 154148 158588 154154
rect 158536 154090 158588 154096
rect 158548 151980 158576 154090
rect 159192 151980 159220 163406
rect 159822 163200 159878 164000
rect 160742 163200 160798 164000
rect 161570 163200 161626 164000
rect 161664 163668 161716 163674
rect 161664 163610 161716 163616
rect 159836 160954 159864 163200
rect 160756 162382 160784 163200
rect 160744 162376 160796 162382
rect 160744 162318 160796 162324
rect 161584 161702 161612 163200
rect 161572 161696 161624 161702
rect 161572 161638 161624 161644
rect 159824 160948 159876 160954
rect 159824 160890 159876 160896
rect 161018 157992 161074 158001
rect 161018 157927 161074 157936
rect 159822 156768 159878 156777
rect 159822 156703 159878 156712
rect 159836 151980 159864 156703
rect 160466 152688 160522 152697
rect 160466 152623 160522 152632
rect 160480 151980 160508 152623
rect 161032 151980 161060 157927
rect 161676 151980 161704 163610
rect 162398 163200 162454 164000
rect 163318 163200 163374 164000
rect 164146 163200 164202 164000
rect 164240 163600 164292 163606
rect 164240 163542 164292 163548
rect 162412 159458 162440 163200
rect 163332 161430 163360 163200
rect 164160 162314 164188 163200
rect 164148 162308 164200 162314
rect 164148 162250 164200 162256
rect 163320 161424 163372 161430
rect 163320 161366 163372 161372
rect 162400 159452 162452 159458
rect 162400 159394 162452 159400
rect 162306 156904 162362 156913
rect 162306 156839 162362 156848
rect 162320 151980 162348 156839
rect 162952 155440 163004 155446
rect 162952 155382 163004 155388
rect 162964 151980 162992 155382
rect 163596 153876 163648 153882
rect 163596 153818 163648 153824
rect 163608 151980 163636 153818
rect 164252 151980 164280 163542
rect 165066 163200 165122 164000
rect 165620 163736 165672 163742
rect 165620 163678 165672 163684
rect 164882 158672 164938 158681
rect 164882 158607 164938 158616
rect 164896 151980 164924 158607
rect 165080 155378 165108 163200
rect 165528 160268 165580 160274
rect 165528 160210 165580 160216
rect 165068 155372 165120 155378
rect 165068 155314 165120 155320
rect 165540 151980 165568 160210
rect 165632 156466 165660 163678
rect 165894 163200 165950 164000
rect 166814 163200 166870 164000
rect 167642 163200 167698 164000
rect 167736 163464 167788 163470
rect 167736 163406 167788 163412
rect 165908 162586 165936 163200
rect 165896 162580 165948 162586
rect 165896 162522 165948 162528
rect 166828 161022 166856 163200
rect 167656 163146 167684 163200
rect 167748 163146 167776 163406
rect 168470 163200 168526 164000
rect 169300 163804 169352 163810
rect 169300 163746 169352 163752
rect 167656 163118 167776 163146
rect 166816 161016 166868 161022
rect 166816 160958 166868 160964
rect 167460 160200 167512 160206
rect 167460 160142 167512 160148
rect 166170 157448 166226 157457
rect 166170 157383 166226 157392
rect 165620 156460 165672 156466
rect 165620 156402 165672 156408
rect 166184 151980 166212 157383
rect 166816 156460 166868 156466
rect 166816 156402 166868 156408
rect 166828 151980 166856 156402
rect 167472 151980 167500 160142
rect 168104 158296 168156 158302
rect 168104 158238 168156 158244
rect 168116 151980 168144 158238
rect 168484 158234 168512 163200
rect 168748 158296 168800 158302
rect 168748 158238 168800 158244
rect 168472 158228 168524 158234
rect 168472 158170 168524 158176
rect 168760 151980 168788 158238
rect 169312 156618 169340 163746
rect 169390 163200 169446 164000
rect 170218 163200 170274 164000
rect 171138 163200 171194 164000
rect 171876 163872 171928 163878
rect 171876 163814 171928 163820
rect 169404 161474 169432 163200
rect 169404 161446 169524 161474
rect 169312 156590 169432 156618
rect 169404 151980 169432 156590
rect 169496 153882 169524 161446
rect 170232 160682 170260 163200
rect 170220 160676 170272 160682
rect 170220 160618 170272 160624
rect 171046 159352 171102 159361
rect 171046 159287 171102 159296
rect 171060 157298 171088 159287
rect 171152 158386 171180 163200
rect 171152 158358 171456 158386
rect 171060 157270 171364 157298
rect 170034 157176 170090 157185
rect 170034 157111 170090 157120
rect 169484 153876 169536 153882
rect 169484 153818 169536 153824
rect 170048 151980 170076 157111
rect 170678 157040 170734 157049
rect 170678 156975 170734 156984
rect 170692 151980 170720 156975
rect 171336 151980 171364 157270
rect 171428 155446 171456 158358
rect 171888 156618 171916 163814
rect 171966 163200 172022 164000
rect 172886 163200 172942 164000
rect 173714 163200 173770 164000
rect 174452 163940 174504 163946
rect 174452 163882 174504 163888
rect 171980 161474 172008 163200
rect 172796 162444 172848 162450
rect 172796 162386 172848 162392
rect 171980 161446 172100 161474
rect 172072 156641 172100 161446
rect 172058 156632 172114 156641
rect 171888 156590 172008 156618
rect 171416 155440 171468 155446
rect 171416 155382 171468 155388
rect 171980 151980 172008 156590
rect 172808 156618 172836 162386
rect 172900 158778 172928 163200
rect 173728 160614 173756 163200
rect 174464 161474 174492 163882
rect 174542 163200 174598 164000
rect 175462 163200 175518 164000
rect 176290 163200 176346 164000
rect 177120 163940 177172 163946
rect 177120 163882 177172 163888
rect 174556 162450 174584 163200
rect 174544 162444 174596 162450
rect 174544 162386 174596 162392
rect 174464 161446 174584 161474
rect 173716 160608 173768 160614
rect 173716 160550 173768 160556
rect 174082 159624 174138 159633
rect 174082 159559 174138 159568
rect 172888 158772 172940 158778
rect 172888 158714 172940 158720
rect 173348 158772 173400 158778
rect 173348 158714 173400 158720
rect 172808 156590 173296 156618
rect 172058 156567 172114 156576
rect 172612 155508 172664 155514
rect 172612 155450 172664 155456
rect 172624 151980 172652 155450
rect 173268 151980 173296 156590
rect 173360 153921 173388 158714
rect 173900 158364 173952 158370
rect 173900 158306 173952 158312
rect 173346 153912 173402 153921
rect 173346 153847 173402 153856
rect 173912 151980 173940 158306
rect 174096 155990 174124 159559
rect 174084 155984 174136 155990
rect 174084 155926 174136 155932
rect 174556 151980 174584 161446
rect 175476 158302 175504 163200
rect 175830 160032 175886 160041
rect 175830 159967 175886 159976
rect 175464 158296 175516 158302
rect 175464 158238 175516 158244
rect 175188 156868 175240 156874
rect 175188 156810 175240 156816
rect 175200 151980 175228 156810
rect 175844 155106 175872 159967
rect 175832 155100 175884 155106
rect 175832 155042 175884 155048
rect 176304 153785 176332 163200
rect 176476 155984 176528 155990
rect 176476 155926 176528 155932
rect 176290 153776 176346 153785
rect 176290 153711 176346 153720
rect 175832 153128 175884 153134
rect 175832 153070 175884 153076
rect 175844 151980 175872 153070
rect 176488 151980 176516 155926
rect 177132 151980 177160 163882
rect 177210 163200 177266 164000
rect 178038 163200 178094 164000
rect 178866 163200 178922 164000
rect 179786 163200 179842 164000
rect 180614 163200 180670 164000
rect 181534 163200 181590 164000
rect 182362 163200 182418 164000
rect 183282 163200 183338 164000
rect 184110 163200 184166 164000
rect 184938 163200 184994 164000
rect 185858 163200 185914 164000
rect 186686 163200 186742 164000
rect 187606 163200 187662 164000
rect 188434 163200 188490 164000
rect 189354 163200 189410 164000
rect 190182 163200 190238 164000
rect 191010 163200 191066 164000
rect 191930 163200 191986 164000
rect 192758 163200 192814 164000
rect 193678 163200 193734 164000
rect 194506 163200 194562 164000
rect 195334 163200 195390 164000
rect 196254 163200 196310 164000
rect 197082 163200 197138 164000
rect 198002 163200 198058 164000
rect 198830 163200 198886 164000
rect 199750 163200 199806 164000
rect 200578 163200 200634 164000
rect 201406 163200 201462 164000
rect 202326 163200 202382 164000
rect 203154 163200 203210 164000
rect 204074 163200 204130 164000
rect 204902 163200 204958 164000
rect 205822 163200 205878 164000
rect 206650 163200 206706 164000
rect 207478 163200 207534 164000
rect 208398 163200 208454 164000
rect 209226 163200 209282 164000
rect 210146 163200 210202 164000
rect 210974 163200 211030 164000
rect 211804 163260 211856 163266
rect 211804 163202 211856 163208
rect 177224 153134 177252 163200
rect 178052 161770 178080 163200
rect 178040 161764 178092 161770
rect 178040 161706 178092 161712
rect 178880 158370 178908 163200
rect 179696 162512 179748 162518
rect 179696 162454 179748 162460
rect 179052 161084 179104 161090
rect 179052 161026 179104 161032
rect 178868 158364 178920 158370
rect 178868 158306 178920 158312
rect 178406 155680 178462 155689
rect 178406 155615 178462 155624
rect 177762 155544 177818 155553
rect 177762 155479 177818 155488
rect 177212 153128 177264 153134
rect 177212 153070 177264 153076
rect 177776 151980 177804 155479
rect 178420 151980 178448 155615
rect 179064 151980 179092 161026
rect 179708 151980 179736 162454
rect 179800 153950 179828 163200
rect 180628 161090 180656 163200
rect 180616 161084 180668 161090
rect 180616 161026 180668 161032
rect 180982 159488 181038 159497
rect 180982 159423 181038 159432
rect 180340 155576 180392 155582
rect 180340 155518 180392 155524
rect 179788 153944 179840 153950
rect 179788 153886 179840 153892
rect 180352 151980 180380 155518
rect 180996 151980 181024 159423
rect 181548 155514 181576 163200
rect 182272 162648 182324 162654
rect 182272 162590 182324 162596
rect 181626 160984 181682 160993
rect 181626 160919 181682 160928
rect 181536 155508 181588 155514
rect 181536 155450 181588 155456
rect 181640 151980 181668 160919
rect 182284 151980 182312 162590
rect 182376 161838 182404 163200
rect 182364 161832 182416 161838
rect 182364 161774 182416 161780
rect 183296 154057 183324 163200
rect 183560 162716 183612 162722
rect 183560 162658 183612 162664
rect 183468 159724 183520 159730
rect 183468 159666 183520 159672
rect 183480 156466 183508 159666
rect 183572 156874 183600 162658
rect 183650 160848 183706 160857
rect 183650 160783 183706 160792
rect 183560 156868 183612 156874
rect 183560 156810 183612 156816
rect 183468 156460 183520 156466
rect 183468 156402 183520 156408
rect 183664 156346 183692 160783
rect 183572 156318 183692 156346
rect 183282 154048 183338 154057
rect 183282 153983 183338 153992
rect 182916 153196 182968 153202
rect 182916 153138 182968 153144
rect 182928 151980 182956 153138
rect 183572 151980 183600 156318
rect 184124 153202 184152 163200
rect 184952 162654 184980 163200
rect 184940 162648 184992 162654
rect 184940 162590 184992 162596
rect 184202 159760 184258 159769
rect 185872 159730 185900 163200
rect 186596 162852 186648 162858
rect 186596 162794 186648 162800
rect 186228 159928 186280 159934
rect 186228 159870 186280 159876
rect 184202 159695 184258 159704
rect 185860 159724 185912 159730
rect 184112 153196 184164 153202
rect 184112 153138 184164 153144
rect 184216 151980 184244 159695
rect 185860 159666 185912 159672
rect 185492 157004 185544 157010
rect 185492 156946 185544 156952
rect 184848 156868 184900 156874
rect 184848 156810 184900 156816
rect 184860 151980 184888 156810
rect 185504 151980 185532 156946
rect 186240 155106 186268 159870
rect 186504 158432 186556 158438
rect 186504 158374 186556 158380
rect 186516 155122 186544 158374
rect 186608 156618 186636 162794
rect 186700 158778 186728 163200
rect 187620 160721 187648 163200
rect 188344 162784 188396 162790
rect 188344 162726 188396 162732
rect 187606 160712 187662 160721
rect 187606 160647 187662 160656
rect 186688 158772 186740 158778
rect 186688 158714 186740 158720
rect 187608 158772 187660 158778
rect 187608 158714 187660 158720
rect 186608 156590 187464 156618
rect 186136 155100 186188 155106
rect 186136 155042 186188 155048
rect 186228 155100 186280 155106
rect 186516 155094 186820 155122
rect 186228 155042 186280 155048
rect 186148 151980 186176 155042
rect 186792 151980 186820 155094
rect 187436 151980 187464 156590
rect 187620 154018 187648 158714
rect 188068 156936 188120 156942
rect 188068 156878 188120 156884
rect 187608 154012 187660 154018
rect 187608 153954 187660 153960
rect 188080 151980 188108 156878
rect 188356 156618 188384 162726
rect 188448 156874 188476 163200
rect 189264 162920 189316 162926
rect 189264 162862 189316 162868
rect 189172 161152 189224 161158
rect 189172 161094 189224 161100
rect 188436 156868 188488 156874
rect 188436 156810 188488 156816
rect 188356 156590 188752 156618
rect 188724 151980 188752 156590
rect 189184 156482 189212 161094
rect 189276 156618 189304 162862
rect 189368 158438 189396 163200
rect 189356 158432 189408 158438
rect 189356 158374 189408 158380
rect 189276 156590 190040 156618
rect 189184 156454 189396 156482
rect 189368 151980 189396 156454
rect 190012 151980 190040 156590
rect 190196 154193 190224 163200
rect 191024 161158 191052 163200
rect 191012 161152 191064 161158
rect 191012 161094 191064 161100
rect 191838 161120 191894 161129
rect 191838 161055 191894 161064
rect 190644 157072 190696 157078
rect 190644 157014 190696 157020
rect 190182 154184 190238 154193
rect 190182 154119 190238 154128
rect 190656 151980 190684 157014
rect 191288 156460 191340 156466
rect 191288 156402 191340 156408
rect 191300 151980 191328 156402
rect 191852 151980 191880 161055
rect 191944 156942 191972 163200
rect 192484 163056 192536 163062
rect 192484 162998 192536 163004
rect 191932 156936 191984 156942
rect 191932 156878 191984 156884
rect 192496 151980 192524 162998
rect 192772 157010 192800 163200
rect 192760 157004 192812 157010
rect 192760 156946 192812 156952
rect 193128 155644 193180 155650
rect 193128 155586 193180 155592
rect 193140 151980 193168 155586
rect 193692 154329 193720 163200
rect 194520 159361 194548 163200
rect 195060 163124 195112 163130
rect 195060 163066 195112 163072
rect 194692 162988 194744 162994
rect 194692 162930 194744 162936
rect 194506 159352 194562 159361
rect 194506 159287 194562 159296
rect 193770 158128 193826 158137
rect 193770 158063 193826 158072
rect 193678 154320 193734 154329
rect 193678 154255 193734 154264
rect 193784 151980 193812 158063
rect 194704 156602 194732 162930
rect 194692 156596 194744 156602
rect 194692 156538 194744 156544
rect 194416 152584 194468 152590
rect 194416 152526 194468 152532
rect 194428 151980 194456 152526
rect 195072 151980 195100 163066
rect 195348 155582 195376 163200
rect 196268 159934 196296 163200
rect 196992 161220 197044 161226
rect 196992 161162 197044 161168
rect 196256 159928 196308 159934
rect 196256 159870 196308 159876
rect 195704 156596 195756 156602
rect 195704 156538 195756 156544
rect 195336 155576 195388 155582
rect 195336 155518 195388 155524
rect 195716 151980 195744 156538
rect 196348 155100 196400 155106
rect 196348 155042 196400 155048
rect 196360 151980 196388 155042
rect 197004 151980 197032 161162
rect 197096 154465 197124 163200
rect 197358 159216 197414 159225
rect 197358 159151 197414 159160
rect 197372 155650 197400 159151
rect 197636 156460 197688 156466
rect 197636 156402 197688 156408
rect 197360 155644 197412 155650
rect 197360 155586 197412 155592
rect 197082 154456 197138 154465
rect 197082 154391 197138 154400
rect 197648 151980 197676 156402
rect 198016 152590 198044 163200
rect 198740 159316 198792 159322
rect 198740 159258 198792 159264
rect 198752 155718 198780 159258
rect 198844 156602 198872 163200
rect 199764 161226 199792 163200
rect 199752 161220 199804 161226
rect 199752 161162 199804 161168
rect 198832 156596 198884 156602
rect 198832 156538 198884 156544
rect 200210 155952 200266 155961
rect 200210 155887 200266 155896
rect 198280 155712 198332 155718
rect 198280 155654 198332 155660
rect 198740 155712 198792 155718
rect 198740 155654 198792 155660
rect 198004 152584 198056 152590
rect 198004 152526 198056 152532
rect 198292 151980 198320 155654
rect 199568 152652 199620 152658
rect 199568 152594 199620 152600
rect 198922 152552 198978 152561
rect 198922 152487 198978 152496
rect 198936 151980 198964 152487
rect 199580 151980 199608 152594
rect 200224 151980 200252 155887
rect 200592 154086 200620 163200
rect 201314 159896 201370 159905
rect 201314 159831 201370 159840
rect 200854 155816 200910 155825
rect 201328 155802 201356 159831
rect 201420 159497 201448 163200
rect 202236 163192 202288 163198
rect 202236 163134 202288 163140
rect 202142 161256 202198 161265
rect 202142 161191 202198 161200
rect 201406 159488 201462 159497
rect 201406 159423 201462 159432
rect 201328 155774 201540 155802
rect 200854 155751 200910 155760
rect 200580 154080 200632 154086
rect 200580 154022 200632 154028
rect 200868 151980 200896 155751
rect 201512 151980 201540 155774
rect 202156 151980 202184 161191
rect 202248 156618 202276 163134
rect 202340 157078 202368 163200
rect 202328 157072 202380 157078
rect 202328 157014 202380 157020
rect 202248 156590 202828 156618
rect 202800 151980 202828 156590
rect 203168 155417 203196 163200
rect 204088 161474 204116 163200
rect 204088 161446 204208 161474
rect 204076 155644 204128 155650
rect 204076 155586 204128 155592
rect 203154 155408 203210 155417
rect 203154 155343 203210 155352
rect 203430 155272 203486 155281
rect 203430 155207 203486 155216
rect 203444 151980 203472 155207
rect 204088 151980 204116 155586
rect 204180 154154 204208 161446
rect 204720 159588 204772 159594
rect 204720 159530 204772 159536
rect 204168 154148 204220 154154
rect 204168 154090 204220 154096
rect 204732 151980 204760 159530
rect 204916 155650 204944 163200
rect 205364 159656 205416 159662
rect 205364 159598 205416 159604
rect 204904 155644 204956 155650
rect 204904 155586 204956 155592
rect 205376 151980 205404 159598
rect 205836 157282 205864 163200
rect 206664 158506 206692 163200
rect 207296 159520 207348 159526
rect 207296 159462 207348 159468
rect 206008 158500 206060 158506
rect 206008 158442 206060 158448
rect 206652 158500 206704 158506
rect 206652 158442 206704 158448
rect 205824 157276 205876 157282
rect 205824 157218 205876 157224
rect 206020 151980 206048 158442
rect 206652 157208 206704 157214
rect 206652 157150 206704 157156
rect 206664 151980 206692 157150
rect 207308 151980 207336 159462
rect 207492 154222 207520 163200
rect 207940 161288 207992 161294
rect 207940 161230 207992 161236
rect 207480 154216 207532 154222
rect 207480 154158 207532 154164
rect 207952 151980 207980 161230
rect 208412 152658 208440 163200
rect 209240 157214 209268 163200
rect 210160 159526 210188 163200
rect 210148 159520 210200 159526
rect 210148 159462 210200 159468
rect 209870 158264 209926 158273
rect 209870 158199 209926 158208
rect 209228 157208 209280 157214
rect 209228 157150 209280 157156
rect 208584 156460 208636 156466
rect 208584 156402 208636 156408
rect 208400 152652 208452 152658
rect 208400 152594 208452 152600
rect 208596 151980 208624 156402
rect 209228 155712 209280 155718
rect 209228 155654 209280 155660
rect 209240 151980 209268 155654
rect 209884 151980 209912 158199
rect 210516 157344 210568 157350
rect 210516 157286 210568 157292
rect 210528 151980 210556 157286
rect 210988 154290 211016 163200
rect 211158 157312 211214 157321
rect 211158 157247 211214 157256
rect 210976 154284 211028 154290
rect 210976 154226 211028 154232
rect 211172 151980 211200 157247
rect 211816 151980 211844 163202
rect 211894 163200 211950 164000
rect 212632 163328 212684 163334
rect 212632 163270 212684 163276
rect 211908 161294 211936 163200
rect 211896 161288 211948 161294
rect 211896 161230 211948 161236
rect 212644 156618 212672 163270
rect 212722 163200 212778 164000
rect 213550 163200 213606 164000
rect 214380 163396 214432 163402
rect 214380 163338 214432 163344
rect 212736 158778 212764 163200
rect 213564 159594 213592 163200
rect 214288 159792 214340 159798
rect 214288 159734 214340 159740
rect 213552 159588 213604 159594
rect 213552 159530 213604 159536
rect 212724 158772 212776 158778
rect 212724 158714 212776 158720
rect 213644 158772 213696 158778
rect 213644 158714 213696 158720
rect 212644 156590 213132 156618
rect 212448 152720 212500 152726
rect 212448 152662 212500 152668
rect 212460 151980 212488 152662
rect 213104 151980 213132 156590
rect 213656 155106 213684 158714
rect 213734 158400 213790 158409
rect 213734 158335 213790 158344
rect 213644 155100 213696 155106
rect 213644 155042 213696 155048
rect 213748 151980 213776 158335
rect 214300 155802 214328 159734
rect 214392 156618 214420 163338
rect 214470 163200 214526 164000
rect 215298 163200 215354 164000
rect 216218 163200 216274 164000
rect 217046 163200 217102 164000
rect 217874 163200 217930 164000
rect 218794 163200 218850 164000
rect 219622 163200 219678 164000
rect 220542 163200 220598 164000
rect 221370 163200 221426 164000
rect 222290 163200 222346 164000
rect 223118 163200 223174 164000
rect 223224 163254 223436 163282
rect 214484 158778 214512 163200
rect 214472 158772 214524 158778
rect 214472 158714 214524 158720
rect 215116 158772 215168 158778
rect 215116 158714 215168 158720
rect 214392 156590 215064 156618
rect 214300 155774 214420 155802
rect 214392 151980 214420 155774
rect 215036 151980 215064 156590
rect 215128 154358 215156 158714
rect 215116 154352 215168 154358
rect 215116 154294 215168 154300
rect 215312 152726 215340 163200
rect 216232 155718 216260 163200
rect 216954 161392 217010 161401
rect 216954 161327 217010 161336
rect 216220 155712 216272 155718
rect 216220 155654 216272 155660
rect 215666 155136 215722 155145
rect 215666 155071 215722 155080
rect 215300 152720 215352 152726
rect 215300 152662 215352 152668
rect 215680 151980 215708 155071
rect 216312 155032 216364 155038
rect 216312 154974 216364 154980
rect 216324 151980 216352 154974
rect 216968 151980 216996 161327
rect 217060 157350 217088 163200
rect 217048 157344 217100 157350
rect 217048 157286 217100 157292
rect 217888 154426 217916 163200
rect 218244 159860 218296 159866
rect 218244 159802 218296 159808
rect 217876 154420 217928 154426
rect 217876 154362 217928 154368
rect 217600 152788 217652 152794
rect 217600 152730 217652 152736
rect 217612 151980 217640 152730
rect 218256 151980 218284 159802
rect 218808 152794 218836 163200
rect 219636 158574 219664 163200
rect 220176 161356 220228 161362
rect 220176 161298 220228 161304
rect 218888 158568 218940 158574
rect 218888 158510 218940 158516
rect 219624 158568 219676 158574
rect 219624 158510 219676 158516
rect 218796 152788 218848 152794
rect 218796 152730 218848 152736
rect 218900 151980 218928 158510
rect 219532 155916 219584 155922
rect 219532 155858 219584 155864
rect 219544 151980 219572 155858
rect 220188 151980 220216 161298
rect 220556 158794 220584 163200
rect 221280 161968 221332 161974
rect 221280 161910 221332 161916
rect 220556 158766 220952 158794
rect 220924 155854 220952 158766
rect 221292 156618 221320 161910
rect 221384 159662 221412 163200
rect 221372 159656 221424 159662
rect 221372 159598 221424 159604
rect 221292 156590 222148 156618
rect 221464 156528 221516 156534
rect 221464 156470 221516 156476
rect 220820 155848 220872 155854
rect 220820 155790 220872 155796
rect 220912 155848 220964 155854
rect 220912 155790 220964 155796
rect 220832 151980 220860 155790
rect 221476 151980 221504 156470
rect 222120 151980 222148 156590
rect 222304 152930 222332 163200
rect 223132 163146 223160 163200
rect 223224 163146 223252 163254
rect 223132 163118 223252 163146
rect 223028 161900 223080 161906
rect 223028 161842 223080 161848
rect 223040 156618 223068 161842
rect 223040 156590 223344 156618
rect 222292 152924 222344 152930
rect 222292 152866 222344 152872
rect 222660 152856 222712 152862
rect 222660 152798 222712 152804
rect 222672 151980 222700 152798
rect 223316 151980 223344 156590
rect 223408 156534 223436 163254
rect 223946 163200 224002 164000
rect 224866 163200 224922 164000
rect 225694 163200 225750 164000
rect 226614 163200 226670 164000
rect 227442 163200 227498 164000
rect 228362 163200 228418 164000
rect 229190 163200 229246 164000
rect 230018 163200 230074 164000
rect 230938 163200 230994 164000
rect 231766 163200 231822 164000
rect 232686 163200 232742 164000
rect 233514 163200 233570 164000
rect 234342 163200 234398 164000
rect 235262 163200 235318 164000
rect 236090 163200 236146 164000
rect 237010 163200 237066 164000
rect 237838 163200 237894 164000
rect 238758 163200 238814 164000
rect 239586 163200 239642 164000
rect 240414 163200 240470 164000
rect 241334 163200 241390 164000
rect 242162 163200 242218 164000
rect 243082 163200 243138 164000
rect 243910 163200 243966 164000
rect 244830 163200 244886 164000
rect 245658 163200 245714 164000
rect 246486 163200 246542 164000
rect 247406 163200 247462 164000
rect 248234 163200 248290 164000
rect 249154 163200 249210 164000
rect 249982 163200 250038 164000
rect 250902 163200 250958 164000
rect 251730 163200 251786 164000
rect 252558 163200 252614 164000
rect 253478 163200 253534 164000
rect 254124 163464 254176 163470
rect 254124 163406 254176 163412
rect 223960 159050 223988 163200
rect 223948 159044 224000 159050
rect 223948 158986 224000 158992
rect 224592 158704 224644 158710
rect 224592 158646 224644 158652
rect 223946 158536 224002 158545
rect 223946 158471 224002 158480
rect 223396 156528 223448 156534
rect 223396 156470 223448 156476
rect 223960 151980 223988 158471
rect 224604 151980 224632 158646
rect 224880 154494 224908 163200
rect 225708 161362 225736 163200
rect 225696 161356 225748 161362
rect 225696 161298 225748 161304
rect 225052 159996 225104 160002
rect 225052 159938 225104 159944
rect 224960 159588 225012 159594
rect 224960 159530 225012 159536
rect 224972 157826 225000 159530
rect 224960 157820 225012 157826
rect 224960 157762 225012 157768
rect 225064 154834 225092 159938
rect 226524 157956 226576 157962
rect 226524 157898 226576 157904
rect 225880 155168 225932 155174
rect 225880 155110 225932 155116
rect 225052 154828 225104 154834
rect 225052 154770 225104 154776
rect 224868 154488 224920 154494
rect 224868 154430 224920 154436
rect 225234 152960 225290 152969
rect 225234 152895 225290 152904
rect 225248 151980 225276 152895
rect 225892 151980 225920 155110
rect 226536 151980 226564 157898
rect 226628 155922 226656 163200
rect 227456 158794 227484 163200
rect 228376 159594 228404 163200
rect 228364 159588 228416 159594
rect 228364 159530 228416 159536
rect 227456 158766 227760 158794
rect 226616 155916 226668 155922
rect 226616 155858 226668 155864
rect 227168 154828 227220 154834
rect 227168 154770 227220 154776
rect 227180 151980 227208 154770
rect 227732 152522 227760 158766
rect 229100 158636 229152 158642
rect 229100 158578 229152 158584
rect 227810 152824 227866 152833
rect 227810 152759 227866 152768
rect 227720 152516 227772 152522
rect 227720 152458 227772 152464
rect 227824 151980 227852 152759
rect 228456 152380 228508 152386
rect 228456 152322 228508 152328
rect 228468 151980 228496 152322
rect 229112 151980 229140 158578
rect 229204 152930 229232 163200
rect 230032 158642 230060 163200
rect 230952 158778 230980 163200
rect 231780 161474 231808 163200
rect 231596 161446 231808 161474
rect 230940 158772 230992 158778
rect 230940 158714 230992 158720
rect 230020 158636 230072 158642
rect 230020 158578 230072 158584
rect 231032 156664 231084 156670
rect 231032 156606 231084 156612
rect 229742 156496 229798 156505
rect 229742 156431 229798 156440
rect 229192 152924 229244 152930
rect 229192 152866 229244 152872
rect 229756 151980 229784 156431
rect 230388 152312 230440 152318
rect 230388 152254 230440 152260
rect 230400 151980 230428 152254
rect 231044 151980 231072 156606
rect 231596 154562 231624 161446
rect 232700 160750 232728 163200
rect 233424 162036 233476 162042
rect 233424 161978 233476 161984
rect 232964 160812 233016 160818
rect 232964 160754 233016 160760
rect 232688 160744 232740 160750
rect 232688 160686 232740 160692
rect 232320 160064 232372 160070
rect 232320 160006 232372 160012
rect 231768 159044 231820 159050
rect 231768 158986 231820 158992
rect 231780 157146 231808 158986
rect 231676 157140 231728 157146
rect 231676 157082 231728 157088
rect 231768 157140 231820 157146
rect 231768 157082 231820 157088
rect 231584 154556 231636 154562
rect 231584 154498 231636 154504
rect 231688 151980 231716 157082
rect 232332 151980 232360 160006
rect 232976 151980 233004 160754
rect 233436 156618 233464 161978
rect 233528 156738 233556 163200
rect 234356 159118 234384 163200
rect 234896 162104 234948 162110
rect 234896 162046 234948 162052
rect 234344 159112 234396 159118
rect 234344 159054 234396 159060
rect 234252 158024 234304 158030
rect 234252 157966 234304 157972
rect 233516 156732 233568 156738
rect 233516 156674 233568 156680
rect 233436 156590 233648 156618
rect 233620 151980 233648 156590
rect 234264 151980 234292 157966
rect 234908 151980 234936 162046
rect 235276 159866 235304 163200
rect 235264 159860 235316 159866
rect 235264 159802 235316 159808
rect 236104 152998 236132 163200
rect 236828 158092 236880 158098
rect 236828 158034 236880 158040
rect 236184 156460 236236 156466
rect 236184 156402 236236 156408
rect 235540 152992 235592 152998
rect 235540 152934 235592 152940
rect 236092 152992 236144 152998
rect 236092 152934 236144 152940
rect 235552 151980 235580 152934
rect 236196 151980 236224 156402
rect 236840 151980 236868 158034
rect 237024 155174 237052 163200
rect 237852 158914 237880 163200
rect 238116 160540 238168 160546
rect 238116 160482 238168 160488
rect 237840 158908 237892 158914
rect 237840 158850 237892 158856
rect 237472 155236 237524 155242
rect 237472 155178 237524 155184
rect 237012 155168 237064 155174
rect 237012 155110 237064 155116
rect 237484 151980 237512 155178
rect 238128 151980 238156 160482
rect 238772 159798 238800 163200
rect 238852 161492 238904 161498
rect 238852 161434 238904 161440
rect 238760 159792 238812 159798
rect 238760 159734 238812 159740
rect 238668 159248 238720 159254
rect 238668 159190 238720 159196
rect 238680 154574 238708 159190
rect 238760 154624 238812 154630
rect 238680 154572 238760 154574
rect 238680 154566 238812 154572
rect 238680 154546 238800 154566
rect 238864 154442 238892 161434
rect 239600 160818 239628 163200
rect 240324 162240 240376 162246
rect 240324 162182 240376 162188
rect 239588 160812 239640 160818
rect 239588 160754 239640 160760
rect 240048 158908 240100 158914
rect 240048 158850 240100 158856
rect 239404 158160 239456 158166
rect 239404 158102 239456 158108
rect 238772 154414 238892 154442
rect 238772 151980 238800 154414
rect 239416 151980 239444 158102
rect 240060 158098 240088 158850
rect 240048 158092 240100 158098
rect 240048 158034 240100 158040
rect 240336 156618 240364 162182
rect 240428 156738 240456 163200
rect 241348 158794 241376 163200
rect 241348 158766 241560 158794
rect 240416 156732 240468 156738
rect 240416 156674 240468 156680
rect 240336 156590 240732 156618
rect 240048 154624 240100 154630
rect 240048 154566 240100 154572
rect 240060 151980 240088 154566
rect 240704 151980 240732 156590
rect 241336 155780 241388 155786
rect 241336 155722 241388 155728
rect 241348 151980 241376 155722
rect 241532 152386 241560 158766
rect 241980 155304 242032 155310
rect 241980 155246 242032 155252
rect 241520 152380 241572 152386
rect 241520 152322 241572 152328
rect 241992 151980 242020 155246
rect 242176 153814 242204 163200
rect 243096 161498 243124 163200
rect 243820 162172 243872 162178
rect 243820 162114 243872 162120
rect 243084 161492 243136 161498
rect 243084 161434 243136 161440
rect 243268 160880 243320 160886
rect 243268 160822 243320 160828
rect 242164 153808 242216 153814
rect 242164 153750 242216 153756
rect 242624 152448 242676 152454
rect 242624 152390 242676 152396
rect 242636 151980 242664 152390
rect 243280 151980 243308 160822
rect 243832 156618 243860 162114
rect 243924 158030 243952 163200
rect 244844 159322 244872 163200
rect 245672 160002 245700 163200
rect 246396 161560 246448 161566
rect 246396 161502 246448 161508
rect 245660 159996 245712 160002
rect 245660 159938 245712 159944
rect 245660 159452 245712 159458
rect 245660 159394 245712 159400
rect 245200 159384 245252 159390
rect 245200 159326 245252 159332
rect 244832 159316 244884 159322
rect 244832 159258 244884 159264
rect 243912 158024 243964 158030
rect 243912 157966 243964 157972
rect 244556 156800 244608 156806
rect 244556 156742 244608 156748
rect 243832 156590 243952 156618
rect 243924 151980 243952 156590
rect 244568 151980 244596 156742
rect 245212 151980 245240 159326
rect 245672 155786 245700 159394
rect 246408 156618 246436 161502
rect 246500 160886 246528 163200
rect 247316 161628 247368 161634
rect 247316 161570 247368 161576
rect 246488 160880 246540 160886
rect 246488 160822 246540 160828
rect 247132 157888 247184 157894
rect 247132 157830 247184 157836
rect 246408 156590 246528 156618
rect 245660 155780 245712 155786
rect 245660 155722 245712 155728
rect 245842 152416 245898 152425
rect 245842 152351 245898 152360
rect 245856 151980 245884 152351
rect 246500 151980 246528 156590
rect 247144 151980 247172 157830
rect 247328 156618 247356 161570
rect 247420 158778 247448 163200
rect 248248 159050 248276 163200
rect 249064 162376 249116 162382
rect 249064 162318 249116 162324
rect 248512 161696 248564 161702
rect 248512 161638 248564 161644
rect 248420 160948 248472 160954
rect 248420 160890 248472 160896
rect 248236 159044 248288 159050
rect 248236 158986 248288 158992
rect 247408 158772 247460 158778
rect 247408 158714 247460 158720
rect 247960 158772 248012 158778
rect 247960 158714 248012 158720
rect 247328 156590 247816 156618
rect 247788 151980 247816 156590
rect 247972 155242 248000 158714
rect 247960 155236 248012 155242
rect 247960 155178 248012 155184
rect 248432 151980 248460 160890
rect 248524 156806 248552 161638
rect 248512 156800 248564 156806
rect 248512 156742 248564 156748
rect 249076 151980 249104 162318
rect 249168 153746 249196 163200
rect 249996 160954 250024 163200
rect 249984 160948 250036 160954
rect 249984 160890 250036 160896
rect 250916 158166 250944 163200
rect 251640 162308 251692 162314
rect 251640 162250 251692 162256
rect 250996 161424 251048 161430
rect 250996 161366 251048 161372
rect 250904 158160 250956 158166
rect 250904 158102 250956 158108
rect 249708 156800 249760 156806
rect 249708 156742 249760 156748
rect 249156 153740 249208 153746
rect 249156 153682 249208 153688
rect 249720 151980 249748 156742
rect 250352 155780 250404 155786
rect 250352 155722 250404 155728
rect 250364 151980 250392 155722
rect 251008 151980 251036 161366
rect 251088 159044 251140 159050
rect 251088 158986 251140 158992
rect 251100 155417 251128 158986
rect 251086 155408 251142 155417
rect 251086 155343 251142 155352
rect 251652 151980 251680 162250
rect 251744 159186 251772 163200
rect 252572 159390 252600 163200
rect 252928 162580 252980 162586
rect 252928 162522 252980 162528
rect 252560 159384 252612 159390
rect 252560 159326 252612 159332
rect 251732 159180 251784 159186
rect 251732 159122 251784 159128
rect 252284 155372 252336 155378
rect 252284 155314 252336 155320
rect 252296 151980 252324 155314
rect 252940 151980 252968 162522
rect 253492 161430 253520 163200
rect 253480 161424 253532 161430
rect 253480 161366 253532 161372
rect 253480 161016 253532 161022
rect 253480 160958 253532 160964
rect 253204 159112 253256 159118
rect 253204 159054 253256 159060
rect 253216 156466 253244 159054
rect 253204 156460 253256 156466
rect 253204 156402 253256 156408
rect 253492 151980 253520 160958
rect 254032 158228 254084 158234
rect 254032 158170 254084 158176
rect 254044 157418 254072 158170
rect 254032 157412 254084 157418
rect 254032 157354 254084 157360
rect 254136 151980 254164 163406
rect 254306 163200 254362 164000
rect 255226 163200 255282 164000
rect 256054 163200 256110 164000
rect 256882 163200 256938 164000
rect 257802 163200 257858 164000
rect 258630 163200 258686 164000
rect 259550 163200 259606 164000
rect 260378 163200 260434 164000
rect 261298 163200 261354 164000
rect 262126 163200 262182 164000
rect 262954 163200 263010 164000
rect 263060 163254 263272 163282
rect 254320 158234 254348 163200
rect 255240 161022 255268 163200
rect 255228 161016 255280 161022
rect 255228 160958 255280 160964
rect 255964 160676 256016 160682
rect 255964 160618 256016 160624
rect 254308 158228 254360 158234
rect 254308 158170 254360 158176
rect 254768 157412 254820 157418
rect 254768 157354 254820 157360
rect 254780 151980 254808 157354
rect 255412 153876 255464 153882
rect 255412 153818 255464 153824
rect 255424 151980 255452 153818
rect 255976 153762 256004 160618
rect 256068 153882 256096 163200
rect 256896 160682 256924 163200
rect 256884 160676 256936 160682
rect 256884 160618 256936 160624
rect 257816 157962 257844 163200
rect 258080 162444 258132 162450
rect 258080 162386 258132 162392
rect 257804 157956 257856 157962
rect 257804 157898 257856 157904
rect 258092 156806 258120 162386
rect 258540 160608 258592 160614
rect 258540 160550 258592 160556
rect 258080 156800 258132 156806
rect 258080 156742 258132 156748
rect 257342 156632 257398 156641
rect 257342 156567 257398 156576
rect 256700 155440 256752 155446
rect 256700 155382 256752 155388
rect 256056 153876 256108 153882
rect 256056 153818 256108 153824
rect 255976 153734 256096 153762
rect 256068 151980 256096 153734
rect 256712 151980 256740 155382
rect 257356 151980 257384 156567
rect 258552 156210 258580 160550
rect 258644 159458 258672 163200
rect 259564 160070 259592 163200
rect 259552 160064 259604 160070
rect 259552 160006 259604 160012
rect 258632 159452 258684 159458
rect 258632 159394 258684 159400
rect 259920 158296 259972 158302
rect 259920 158238 259972 158244
rect 259276 156800 259328 156806
rect 259276 156742 259328 156748
rect 258552 156182 258672 156210
rect 257986 153912 258042 153921
rect 257986 153847 258042 153856
rect 258000 151980 258028 153847
rect 258644 151980 258672 156182
rect 259288 151980 259316 156742
rect 259932 151980 259960 158238
rect 260392 155378 260420 163200
rect 261208 161764 261260 161770
rect 261208 161706 261260 161712
rect 260564 159928 260616 159934
rect 260564 159870 260616 159876
rect 260576 157894 260604 159870
rect 260564 157888 260616 157894
rect 260564 157830 260616 157836
rect 261220 156618 261248 161706
rect 261312 158778 261340 163200
rect 262140 158794 262168 163200
rect 262968 163146 262996 163200
rect 263060 163146 263088 163254
rect 262968 163118 263088 163146
rect 261300 158772 261352 158778
rect 261300 158714 261352 158720
rect 261944 158772 261996 158778
rect 262140 158766 262260 158794
rect 261944 158714 261996 158720
rect 261220 156590 261892 156618
rect 260380 155372 260432 155378
rect 260380 155314 260432 155320
rect 260562 153776 260618 153785
rect 260562 153711 260618 153720
rect 260576 151980 260604 153711
rect 261208 153128 261260 153134
rect 261208 153070 261260 153076
rect 261220 151980 261248 153070
rect 261864 151980 261892 156590
rect 261956 155310 261984 158714
rect 261944 155304 261996 155310
rect 261944 155246 261996 155252
rect 262232 152454 262260 158766
rect 262496 158364 262548 158370
rect 262496 158306 262548 158312
rect 262220 152448 262272 152454
rect 262220 152390 262272 152396
rect 262508 151980 262536 158306
rect 263244 153950 263272 163254
rect 263874 163200 263930 164000
rect 264702 163200 264758 164000
rect 265622 163200 265678 164000
rect 266450 163200 266506 164000
rect 267370 163200 267426 164000
rect 268198 163200 268254 164000
rect 269026 163200 269082 164000
rect 269946 163200 270002 164000
rect 270774 163200 270830 164000
rect 271694 163200 271750 164000
rect 272522 163200 272578 164000
rect 273350 163200 273406 164000
rect 274270 163200 274326 164000
rect 274376 163254 274588 163282
rect 263784 161084 263836 161090
rect 263784 161026 263836 161032
rect 263140 153944 263192 153950
rect 263140 153886 263192 153892
rect 263232 153944 263284 153950
rect 263232 153886 263284 153892
rect 263152 151980 263180 153886
rect 263796 151980 263824 161026
rect 263888 160614 263916 163200
rect 263876 160608 263928 160614
rect 263876 160550 263928 160556
rect 264716 158001 264744 163200
rect 265072 161832 265124 161838
rect 265072 161774 265124 161780
rect 264980 159724 265032 159730
rect 264980 159666 265032 159672
rect 264702 157992 264758 158001
rect 264702 157927 264758 157936
rect 264428 155508 264480 155514
rect 264428 155450 264480 155456
rect 264440 151980 264468 155450
rect 264992 154834 265020 159666
rect 264980 154828 265032 154834
rect 264980 154770 265032 154776
rect 265084 151980 265112 161774
rect 265636 161090 265664 163200
rect 265624 161084 265676 161090
rect 265624 161026 265676 161032
rect 266464 159934 266492 163200
rect 267004 162648 267056 162654
rect 267004 162590 267056 162596
rect 266452 159928 266504 159934
rect 266452 159870 266504 159876
rect 265714 154048 265770 154057
rect 265714 153983 265770 153992
rect 265728 151980 265756 153983
rect 266360 153196 266412 153202
rect 266360 153138 266412 153144
rect 266372 151980 266400 153138
rect 267016 151980 267044 162590
rect 267384 155446 267412 163200
rect 268212 158302 268240 163200
rect 268934 160712 268990 160721
rect 268934 160647 268990 160656
rect 268200 158296 268252 158302
rect 268200 158238 268252 158244
rect 267372 155440 267424 155446
rect 267372 155382 267424 155388
rect 267648 154828 267700 154834
rect 267648 154770 267700 154776
rect 267660 151980 267688 154770
rect 268292 154012 268344 154018
rect 268292 153954 268344 153960
rect 268304 151980 268332 153954
rect 268948 151980 268976 160647
rect 269040 159254 269068 163200
rect 269028 159248 269080 159254
rect 269028 159190 269080 159196
rect 269580 156868 269632 156874
rect 269580 156810 269632 156816
rect 269592 151980 269620 156810
rect 269960 154018 269988 163200
rect 270406 159488 270462 159497
rect 270406 159423 270462 159432
rect 270224 158432 270276 158438
rect 270224 158374 270276 158380
rect 269948 154012 270000 154018
rect 269948 153954 270000 153960
rect 270236 151980 270264 158374
rect 270420 158370 270448 159423
rect 270408 158364 270460 158370
rect 270408 158306 270460 158312
rect 270788 155514 270816 163200
rect 271512 161152 271564 161158
rect 271512 161094 271564 161100
rect 270776 155508 270828 155514
rect 270776 155450 270828 155456
rect 270866 154184 270922 154193
rect 270866 154119 270922 154128
rect 270880 151980 270908 154119
rect 271524 151980 271552 161094
rect 271708 156641 271736 163200
rect 272432 159316 272484 159322
rect 272432 159258 272484 159264
rect 272064 159180 272116 159186
rect 272064 159122 272116 159128
rect 271694 156632 271750 156641
rect 271694 156567 271750 156576
rect 272076 156398 272104 159122
rect 272156 156936 272208 156942
rect 272156 156878 272208 156884
rect 272064 156392 272116 156398
rect 272064 156334 272116 156340
rect 272168 151980 272196 156878
rect 272444 156330 272472 159258
rect 272536 159118 272564 163200
rect 273364 159730 273392 163200
rect 274284 163146 274312 163200
rect 274376 163146 274404 163254
rect 274284 163118 274404 163146
rect 273352 159724 273404 159730
rect 273352 159666 273404 159672
rect 274086 159352 274142 159361
rect 274086 159287 274142 159296
rect 272524 159112 272576 159118
rect 272524 159054 272576 159060
rect 272800 157004 272852 157010
rect 272800 156946 272852 156952
rect 272432 156324 272484 156330
rect 272432 156266 272484 156272
rect 272812 151980 272840 156946
rect 273442 154320 273498 154329
rect 273442 154255 273498 154264
rect 273456 151980 273484 154255
rect 274100 151980 274128 159287
rect 274560 153202 274588 163254
rect 275098 163200 275154 164000
rect 276018 163200 276074 164000
rect 276846 163200 276902 164000
rect 277766 163200 277822 164000
rect 278594 163200 278650 164000
rect 279422 163200 279478 164000
rect 280342 163200 280398 164000
rect 281170 163200 281226 164000
rect 282090 163200 282146 164000
rect 282918 163200 282974 164000
rect 283838 163200 283894 164000
rect 284666 163200 284722 164000
rect 285494 163200 285550 164000
rect 286414 163200 286470 164000
rect 287242 163200 287298 164000
rect 288162 163200 288218 164000
rect 288990 163200 289046 164000
rect 289818 163200 289874 164000
rect 290738 163200 290794 164000
rect 291566 163200 291622 164000
rect 292486 163200 292542 164000
rect 293314 163200 293370 164000
rect 294234 163200 294290 164000
rect 295062 163200 295118 164000
rect 295890 163200 295946 164000
rect 296810 163200 296866 164000
rect 297638 163200 297694 164000
rect 298558 163200 298614 164000
rect 299386 163200 299442 164000
rect 300306 163200 300362 164000
rect 301134 163200 301190 164000
rect 301962 163200 302018 164000
rect 302882 163200 302938 164000
rect 303710 163200 303766 164000
rect 304630 163200 304686 164000
rect 304736 163254 304948 163282
rect 275112 155786 275140 163200
rect 276032 159322 276060 163200
rect 276112 159520 276164 159526
rect 276112 159462 276164 159468
rect 276020 159316 276072 159322
rect 276020 159258 276072 159264
rect 275376 157888 275428 157894
rect 275376 157830 275428 157836
rect 275100 155780 275152 155786
rect 275100 155722 275152 155728
rect 274732 155576 274784 155582
rect 274732 155518 274784 155524
rect 274548 153196 274600 153202
rect 274548 153138 274600 153144
rect 274744 151980 274772 155518
rect 275388 151980 275416 157830
rect 276124 156874 276152 159462
rect 276860 158438 276888 163200
rect 276848 158432 276900 158438
rect 276848 158374 276900 158380
rect 276112 156868 276164 156874
rect 276112 156810 276164 156816
rect 277308 156596 277360 156602
rect 277308 156538 277360 156544
rect 276018 154456 276074 154465
rect 276018 154391 276074 154400
rect 276032 151980 276060 154391
rect 276664 152584 276716 152590
rect 276664 152526 276716 152532
rect 276676 151980 276704 152526
rect 277320 151980 277348 156538
rect 277780 155582 277808 163200
rect 277952 161220 278004 161226
rect 277952 161162 278004 161168
rect 277768 155576 277820 155582
rect 277768 155518 277820 155524
rect 277964 151980 277992 161162
rect 278608 156806 278636 163200
rect 279240 158364 279292 158370
rect 279240 158306 279292 158312
rect 278596 156800 278648 156806
rect 278596 156742 278648 156748
rect 278596 154080 278648 154086
rect 278596 154022 278648 154028
rect 278608 151980 278636 154022
rect 279252 151980 279280 158306
rect 279436 152590 279464 163200
rect 280356 159361 280384 163200
rect 280988 159656 281040 159662
rect 280988 159598 281040 159604
rect 280342 159352 280398 159361
rect 280342 159287 280398 159296
rect 279884 157072 279936 157078
rect 279884 157014 279936 157020
rect 279424 152584 279476 152590
rect 279424 152526 279476 152532
rect 279896 151980 279924 157014
rect 280526 155272 280582 155281
rect 280526 155207 280582 155216
rect 280540 151980 280568 155207
rect 281000 153678 281028 159598
rect 281184 158370 281212 163200
rect 281448 158432 281500 158438
rect 281448 158374 281500 158380
rect 281172 158364 281224 158370
rect 281172 158306 281224 158312
rect 281460 154154 281488 158374
rect 282104 155650 282132 163200
rect 282184 159452 282236 159458
rect 282184 159394 282236 159400
rect 282196 156602 282224 159394
rect 282932 159050 282960 163200
rect 283012 159112 283064 159118
rect 283012 159054 283064 159060
rect 282920 159044 282972 159050
rect 282920 158986 282972 158992
rect 283024 157282 283052 159054
rect 283104 158500 283156 158506
rect 283104 158442 283156 158448
rect 282460 157276 282512 157282
rect 282460 157218 282512 157224
rect 283012 157276 283064 157282
rect 283012 157218 283064 157224
rect 282184 156596 282236 156602
rect 282184 156538 282236 156544
rect 281816 155644 281868 155650
rect 281816 155586 281868 155592
rect 282092 155644 282144 155650
rect 282092 155586 282144 155592
rect 281172 154148 281224 154154
rect 281172 154090 281224 154096
rect 281448 154148 281500 154154
rect 281448 154090 281500 154096
rect 280988 153672 281040 153678
rect 280988 153614 281040 153620
rect 281184 151980 281212 154090
rect 281828 151980 281856 155586
rect 282472 151980 282500 157218
rect 283116 151980 283144 158442
rect 283852 157758 283880 163200
rect 284680 158137 284708 163200
rect 284666 158128 284722 158137
rect 284666 158063 284722 158072
rect 283840 157752 283892 157758
rect 283840 157694 283892 157700
rect 284944 157208 284996 157214
rect 284944 157150 284996 157156
rect 283748 154216 283800 154222
rect 283748 154158 283800 154164
rect 283760 151980 283788 154158
rect 284300 152652 284352 152658
rect 284300 152594 284352 152600
rect 284312 151980 284340 152594
rect 284956 151980 284984 157150
rect 285508 156874 285536 163200
rect 286428 158438 286456 163200
rect 286876 161288 286928 161294
rect 286876 161230 286928 161236
rect 286416 158432 286468 158438
rect 286416 158374 286468 158380
rect 285680 157752 285732 157758
rect 285680 157694 285732 157700
rect 285588 156936 285640 156942
rect 285588 156878 285640 156884
rect 285496 156868 285548 156874
rect 285496 156810 285548 156816
rect 285600 151980 285628 156878
rect 285692 154086 285720 157694
rect 286232 154284 286284 154290
rect 286232 154226 286284 154232
rect 285680 154080 285732 154086
rect 285680 154022 285732 154028
rect 286244 151980 286272 154226
rect 286888 151980 286916 161230
rect 287256 158982 287284 163200
rect 288176 161474 288204 163200
rect 288176 161446 288296 161474
rect 287244 158976 287296 158982
rect 287244 158918 287296 158924
rect 288164 157820 288216 157826
rect 288164 157762 288216 157768
rect 287520 155100 287572 155106
rect 287520 155042 287572 155048
rect 287532 151980 287560 155042
rect 288176 151980 288204 157762
rect 288268 155106 288296 161446
rect 289004 156942 289032 163200
rect 289728 159588 289780 159594
rect 289728 159530 289780 159536
rect 288992 156936 289044 156942
rect 288992 156878 289044 156884
rect 288256 155100 288308 155106
rect 288256 155042 288308 155048
rect 288808 154352 288860 154358
rect 288808 154294 288860 154300
rect 288820 151980 288848 154294
rect 289740 154290 289768 159530
rect 289832 159186 289860 163200
rect 289820 159180 289872 159186
rect 289820 159122 289872 159128
rect 290752 158778 290780 163200
rect 291108 159248 291160 159254
rect 291108 159190 291160 159196
rect 290740 158772 290792 158778
rect 290740 158714 290792 158720
rect 290740 157344 290792 157350
rect 290740 157286 290792 157292
rect 290096 155712 290148 155718
rect 290096 155654 290148 155660
rect 289728 154284 289780 154290
rect 289728 154226 289780 154232
rect 289452 152720 289504 152726
rect 289452 152662 289504 152668
rect 289464 151980 289492 152662
rect 290108 151980 290136 155654
rect 290752 151980 290780 157286
rect 291120 155281 291148 159190
rect 291580 157894 291608 163200
rect 291844 159860 291896 159866
rect 291844 159802 291896 159808
rect 291568 157888 291620 157894
rect 291568 157830 291620 157836
rect 291106 155272 291162 155281
rect 291106 155207 291162 155216
rect 291856 154426 291884 159802
rect 292500 156777 292528 163200
rect 293328 159118 293356 163200
rect 294248 159526 294276 163200
rect 294236 159520 294288 159526
rect 294236 159462 294288 159468
rect 293960 159316 294012 159322
rect 293960 159258 294012 159264
rect 293316 159112 293368 159118
rect 293316 159054 293368 159060
rect 292764 158772 292816 158778
rect 292764 158714 292816 158720
rect 292672 158568 292724 158574
rect 292672 158510 292724 158516
rect 292486 156768 292542 156777
rect 292486 156703 292542 156712
rect 291384 154420 291436 154426
rect 291384 154362 291436 154368
rect 291844 154420 291896 154426
rect 291844 154362 291896 154368
rect 291396 151980 291424 154362
rect 292028 152788 292080 152794
rect 292028 152730 292080 152736
rect 292040 151980 292068 152730
rect 292684 151980 292712 158510
rect 292776 154222 292804 158714
rect 293316 155848 293368 155854
rect 293316 155790 293368 155796
rect 292764 154216 292816 154222
rect 292764 154158 292816 154164
rect 293328 151980 293356 155790
rect 293972 155038 294000 159258
rect 295076 158506 295104 163200
rect 295064 158500 295116 158506
rect 295064 158442 295116 158448
rect 295800 157140 295852 157146
rect 295800 157082 295852 157088
rect 295248 156528 295300 156534
rect 295248 156470 295300 156476
rect 293960 155032 294012 155038
rect 293960 154974 294012 154980
rect 293960 153672 294012 153678
rect 293960 153614 294012 153620
rect 293972 151980 294000 153614
rect 294604 152856 294656 152862
rect 294604 152798 294656 152804
rect 294616 151980 294644 152798
rect 295260 151980 295288 156470
rect 295812 154442 295840 157082
rect 295904 157010 295932 163200
rect 296628 159792 296680 159798
rect 296628 159734 296680 159740
rect 295892 157004 295944 157010
rect 295892 156946 295944 156952
rect 296640 154494 296668 159734
rect 296824 159322 296852 163200
rect 297180 161356 297232 161362
rect 297180 161298 297232 161304
rect 296812 159316 296864 159322
rect 296812 159258 296864 159264
rect 296536 154488 296588 154494
rect 295812 154414 295932 154442
rect 296536 154430 296588 154436
rect 296628 154488 296680 154494
rect 296628 154430 296680 154436
rect 295904 151980 295932 154414
rect 296548 151980 296576 154430
rect 297192 151980 297220 161298
rect 297652 155854 297680 163200
rect 297824 155916 297876 155922
rect 297824 155858 297876 155864
rect 297640 155848 297692 155854
rect 297640 155790 297692 155796
rect 297836 151980 297864 155858
rect 298100 155848 298152 155854
rect 298100 155790 298152 155796
rect 298112 154358 298140 155790
rect 298572 155718 298600 163200
rect 299400 157078 299428 163200
rect 299388 157072 299440 157078
rect 299388 157014 299440 157020
rect 298560 155712 298612 155718
rect 298560 155654 298612 155660
rect 298100 154352 298152 154358
rect 298100 154294 298152 154300
rect 300320 154290 300348 163200
rect 301148 159594 301176 163200
rect 301780 159996 301832 160002
rect 301780 159938 301832 159944
rect 301136 159588 301188 159594
rect 301136 159530 301188 159536
rect 301044 158704 301096 158710
rect 301044 158646 301096 158652
rect 300400 158636 300452 158642
rect 300400 158578 300452 158584
rect 299112 154284 299164 154290
rect 299112 154226 299164 154232
rect 300308 154284 300360 154290
rect 300308 154226 300360 154232
rect 298468 152516 298520 152522
rect 298468 152458 298520 152464
rect 298480 151980 298508 152458
rect 299124 151980 299152 154226
rect 299756 152924 299808 152930
rect 299756 152866 299808 152872
rect 299768 151980 299796 152866
rect 300412 151980 300440 158578
rect 301056 151980 301084 158646
rect 301792 154562 301820 159938
rect 301976 158574 302004 163200
rect 302332 160744 302384 160750
rect 302332 160686 302384 160692
rect 301964 158568 302016 158574
rect 301964 158510 302016 158516
rect 301688 154556 301740 154562
rect 301688 154498 301740 154504
rect 301780 154556 301832 154562
rect 301780 154498 301832 154504
rect 301700 151980 301728 154498
rect 302344 151980 302372 160686
rect 302896 155854 302924 163200
rect 303724 159254 303752 163200
rect 304644 163146 304672 163200
rect 304736 163146 304764 163254
rect 304644 163118 304764 163146
rect 303712 159248 303764 159254
rect 303712 159190 303764 159196
rect 302976 156664 303028 156670
rect 302976 156606 303028 156612
rect 302884 155848 302936 155854
rect 302884 155790 302936 155796
rect 302988 151980 303016 156606
rect 303620 156460 303672 156466
rect 303620 156402 303672 156408
rect 303632 151980 303660 156402
rect 304920 154426 304948 163254
rect 305458 163200 305514 164000
rect 306378 163200 306434 164000
rect 307206 163200 307262 164000
rect 308034 163200 308090 164000
rect 308954 163200 309010 164000
rect 309782 163200 309838 164000
rect 310702 163200 310758 164000
rect 311530 163200 311586 164000
rect 312358 163200 312414 164000
rect 313278 163200 313334 164000
rect 314106 163200 314162 164000
rect 315026 163200 315082 164000
rect 315854 163200 315910 164000
rect 316774 163200 316830 164000
rect 317602 163200 317658 164000
rect 318430 163200 318486 164000
rect 319350 163200 319406 164000
rect 320178 163200 320234 164000
rect 321098 163200 321154 164000
rect 321926 163200 321982 164000
rect 322846 163200 322902 164000
rect 323674 163200 323730 164000
rect 324502 163200 324558 164000
rect 325422 163200 325478 164000
rect 326250 163200 326306 164000
rect 327170 163200 327226 164000
rect 327998 163200 328054 164000
rect 328826 163200 328882 164000
rect 329746 163200 329802 164000
rect 330574 163200 330630 164000
rect 331494 163200 331550 164000
rect 332322 163200 332378 164000
rect 333242 163200 333298 164000
rect 334070 163200 334126 164000
rect 334898 163200 334954 164000
rect 335818 163200 335874 164000
rect 336646 163200 336702 164000
rect 337566 163200 337622 164000
rect 338394 163200 338450 164000
rect 339314 163200 339370 164000
rect 340142 163200 340198 164000
rect 340970 163200 341026 164000
rect 341890 163200 341946 164000
rect 342718 163200 342774 164000
rect 343638 163200 343694 164000
rect 344466 163200 344522 164000
rect 345386 163200 345442 164000
rect 346214 163200 346270 164000
rect 347042 163200 347098 164000
rect 347962 163200 348018 164000
rect 348790 163200 348846 164000
rect 349710 163200 349766 164000
rect 350538 163200 350594 164000
rect 351366 163200 351422 164000
rect 352286 163200 352342 164000
rect 353114 163200 353170 164000
rect 354034 163200 354090 164000
rect 354862 163200 354918 164000
rect 355782 163200 355838 164000
rect 356610 163200 356666 164000
rect 357438 163200 357494 164000
rect 358358 163200 358414 164000
rect 359186 163200 359242 164000
rect 360106 163200 360162 164000
rect 360934 163200 360990 164000
rect 361854 163200 361910 164000
rect 362682 163200 362738 164000
rect 363510 163200 363566 164000
rect 364430 163200 364486 164000
rect 365258 163200 365314 164000
rect 366178 163200 366234 164000
rect 367006 163200 367062 164000
rect 367834 163200 367890 164000
rect 368754 163200 368810 164000
rect 369582 163200 369638 164000
rect 370502 163200 370558 164000
rect 371330 163200 371386 164000
rect 372250 163200 372306 164000
rect 373078 163200 373134 164000
rect 373906 163200 373962 164000
rect 374826 163200 374882 164000
rect 375654 163200 375710 164000
rect 376574 163200 376630 164000
rect 377402 163200 377458 164000
rect 378322 163200 378378 164000
rect 379150 163200 379206 164000
rect 379978 163200 380034 164000
rect 380898 163200 380954 164000
rect 381726 163200 381782 164000
rect 382646 163200 382702 164000
rect 383474 163200 383530 164000
rect 384394 163200 384450 164000
rect 385222 163200 385278 164000
rect 386050 163200 386106 164000
rect 386970 163200 387026 164000
rect 387798 163200 387854 164000
rect 388718 163200 388774 164000
rect 389546 163200 389602 164000
rect 390374 163200 390430 164000
rect 391294 163200 391350 164000
rect 392122 163200 392178 164000
rect 393042 163200 393098 164000
rect 393870 163200 393926 164000
rect 394790 163200 394846 164000
rect 395618 163200 395674 164000
rect 396446 163200 396502 164000
rect 397366 163200 397422 164000
rect 398194 163200 398250 164000
rect 399114 163200 399170 164000
rect 399942 163200 399998 164000
rect 400862 163200 400918 164000
rect 401690 163200 401746 164000
rect 402518 163200 402574 164000
rect 403438 163200 403494 164000
rect 404266 163200 404322 164000
rect 405186 163200 405242 164000
rect 406014 163200 406070 164000
rect 406842 163200 406898 164000
rect 407762 163200 407818 164000
rect 408590 163200 408646 164000
rect 409510 163200 409566 164000
rect 410338 163200 410394 164000
rect 411258 163200 411314 164000
rect 412086 163200 412142 164000
rect 412914 163200 412970 164000
rect 413834 163200 413890 164000
rect 414662 163200 414718 164000
rect 415582 163200 415638 164000
rect 416410 163200 416466 164000
rect 417330 163200 417386 164000
rect 418158 163200 418214 164000
rect 418986 163200 419042 164000
rect 419092 163254 419304 163282
rect 305472 158642 305500 163200
rect 305460 158636 305512 158642
rect 305460 158578 305512 158584
rect 306196 158092 306248 158098
rect 306196 158034 306248 158040
rect 305552 155168 305604 155174
rect 305552 155110 305604 155116
rect 304264 154420 304316 154426
rect 304264 154362 304316 154368
rect 304908 154420 304960 154426
rect 304908 154362 304960 154368
rect 304276 151980 304304 154362
rect 304908 152992 304960 152998
rect 304908 152934 304960 152940
rect 304920 151980 304948 152934
rect 305564 151980 305592 155110
rect 306208 151980 306236 158034
rect 306392 157146 306420 163200
rect 307220 158778 307248 163200
rect 307484 160812 307536 160818
rect 307484 160754 307536 160760
rect 307208 158772 307260 158778
rect 307208 158714 307260 158720
rect 306380 157140 306432 157146
rect 306380 157082 306432 157088
rect 306840 153672 306892 153678
rect 306840 153614 306892 153620
rect 306852 151980 306880 153614
rect 307496 151980 307524 160754
rect 308048 159662 308076 163200
rect 308036 159656 308088 159662
rect 308036 159598 308088 159604
rect 308312 159180 308364 159186
rect 308312 159122 308364 159128
rect 308128 156732 308180 156738
rect 308128 156674 308180 156680
rect 308140 151980 308168 156674
rect 308324 156534 308352 159122
rect 308864 158772 308916 158778
rect 308864 158714 308916 158720
rect 308312 156528 308364 156534
rect 308312 156470 308364 156476
rect 308876 154494 308904 158714
rect 308968 158098 308996 163200
rect 309692 161492 309744 161498
rect 309692 161434 309744 161440
rect 308956 158092 309008 158098
rect 308956 158034 309008 158040
rect 309704 156618 309732 161434
rect 309796 156738 309824 163200
rect 310244 159384 310296 159390
rect 310244 159326 310296 159332
rect 309784 156732 309836 156738
rect 309784 156674 309836 156680
rect 309704 156590 310100 156618
rect 308864 154488 308916 154494
rect 308864 154430 308916 154436
rect 309416 153808 309468 153814
rect 309416 153750 309468 153756
rect 308772 152924 308824 152930
rect 308772 152866 308824 152872
rect 308784 151980 308812 152866
rect 309428 151980 309456 153750
rect 310072 151980 310100 156590
rect 310256 153270 310284 159326
rect 310716 159186 310744 163200
rect 310704 159180 310756 159186
rect 310704 159122 310756 159128
rect 311072 159044 311124 159050
rect 311072 158986 311124 158992
rect 310704 158024 310756 158030
rect 310704 157966 310756 157972
rect 310244 153264 310296 153270
rect 310244 153206 310296 153212
rect 310716 151980 310744 157966
rect 311084 155174 311112 158986
rect 311544 158778 311572 163200
rect 311900 160064 311952 160070
rect 311900 160006 311952 160012
rect 311532 158772 311584 158778
rect 311532 158714 311584 158720
rect 311348 156324 311400 156330
rect 311348 156266 311400 156272
rect 311072 155168 311124 155174
rect 311072 155110 311124 155116
rect 311360 151980 311388 156266
rect 311912 153678 311940 160006
rect 312372 158710 312400 163200
rect 312636 160880 312688 160886
rect 312636 160822 312688 160828
rect 312360 158704 312412 158710
rect 312360 158646 312412 158652
rect 311992 154556 312044 154562
rect 311992 154498 312044 154504
rect 311900 153672 311952 153678
rect 311900 153614 311952 153620
rect 312004 151980 312032 154498
rect 312648 151980 312676 160822
rect 313292 156738 313320 163200
rect 314120 158778 314148 163200
rect 315040 159390 315068 163200
rect 315120 160948 315172 160954
rect 315120 160890 315172 160896
rect 315028 159384 315080 159390
rect 315028 159326 315080 159332
rect 313740 158772 313792 158778
rect 313740 158714 313792 158720
rect 314108 158772 314160 158778
rect 314108 158714 314160 158720
rect 313280 156732 313332 156738
rect 313280 156674 313332 156680
rect 313280 155236 313332 155242
rect 313280 155178 313332 155184
rect 313292 151980 313320 155178
rect 313752 154562 313780 158714
rect 313922 155408 313978 155417
rect 313922 155343 313978 155352
rect 313740 154556 313792 154562
rect 313740 154498 313792 154504
rect 313936 151980 313964 155343
rect 314568 153740 314620 153746
rect 314568 153682 314620 153688
rect 314580 151980 314608 153682
rect 315132 151980 315160 160890
rect 315764 158160 315816 158166
rect 315764 158102 315816 158108
rect 315776 151980 315804 158102
rect 315868 158030 315896 163200
rect 316224 159928 316276 159934
rect 316224 159870 316276 159876
rect 315856 158024 315908 158030
rect 315856 157966 315908 157972
rect 316236 153814 316264 159870
rect 316788 157214 316816 163200
rect 317616 159050 317644 163200
rect 317696 161424 317748 161430
rect 317696 161366 317748 161372
rect 317604 159044 317656 159050
rect 317604 158986 317656 158992
rect 316776 157208 316828 157214
rect 316776 157150 316828 157156
rect 316408 156392 316460 156398
rect 316408 156334 316460 156340
rect 316224 153808 316276 153814
rect 316224 153750 316276 153756
rect 316420 151980 316448 156334
rect 317052 153264 317104 153270
rect 317052 153206 317104 153212
rect 317064 151980 317092 153206
rect 317708 151980 317736 161366
rect 318444 158846 318472 163200
rect 318984 161016 319036 161022
rect 318984 160958 319036 160964
rect 318432 158840 318484 158846
rect 318432 158782 318484 158788
rect 318708 158772 318760 158778
rect 318708 158714 318760 158720
rect 318340 158228 318392 158234
rect 318340 158170 318392 158176
rect 318352 151980 318380 158170
rect 318720 157826 318748 158714
rect 318708 157820 318760 157826
rect 318708 157762 318760 157768
rect 318996 151980 319024 160958
rect 319364 155242 319392 163200
rect 320192 158166 320220 163200
rect 320272 160676 320324 160682
rect 320272 160618 320324 160624
rect 320180 158160 320232 158166
rect 320180 158102 320232 158108
rect 319352 155236 319404 155242
rect 319352 155178 319404 155184
rect 319628 153876 319680 153882
rect 319628 153818 319680 153824
rect 319640 151980 319668 153818
rect 320284 151980 320312 160618
rect 321112 158778 321140 163200
rect 321940 159866 321968 163200
rect 321928 159860 321980 159866
rect 321928 159802 321980 159808
rect 321100 158772 321152 158778
rect 321100 158714 321152 158720
rect 321744 158772 321796 158778
rect 321744 158714 321796 158720
rect 320916 157956 320968 157962
rect 320916 157898 320968 157904
rect 320928 151980 320956 157898
rect 321560 156596 321612 156602
rect 321560 156538 321612 156544
rect 321572 151980 321600 156538
rect 321756 153882 321784 158714
rect 322860 158234 322888 163200
rect 322940 159112 322992 159118
rect 322940 159054 322992 159060
rect 322848 158228 322900 158234
rect 322848 158170 322900 158176
rect 322952 155417 322980 159054
rect 322938 155408 322994 155417
rect 322848 155372 322900 155378
rect 322938 155343 322994 155352
rect 322848 155314 322900 155320
rect 321744 153876 321796 153882
rect 321744 153818 321796 153824
rect 322204 153672 322256 153678
rect 322204 153614 322256 153620
rect 322216 151980 322244 153614
rect 322860 151980 322888 155314
rect 323688 155310 323716 163200
rect 324516 159798 324544 163200
rect 325332 160608 325384 160614
rect 325332 160550 325384 160556
rect 324504 159792 324556 159798
rect 324504 159734 324556 159740
rect 324320 158840 324372 158846
rect 324320 158782 324372 158788
rect 323492 155304 323544 155310
rect 323492 155246 323544 155252
rect 323676 155304 323728 155310
rect 323676 155246 323728 155252
rect 323504 151980 323532 155246
rect 324332 153746 324360 158782
rect 324780 153944 324832 153950
rect 324780 153886 324832 153892
rect 324320 153740 324372 153746
rect 324320 153682 324372 153688
rect 324136 153128 324188 153134
rect 324136 153070 324188 153076
rect 324148 151980 324176 153070
rect 324792 151980 324820 153886
rect 325344 153762 325372 160550
rect 325436 153950 325464 163200
rect 326066 157992 326122 158001
rect 326066 157927 326122 157936
rect 325424 153944 325476 153950
rect 325424 153886 325476 153892
rect 325344 153734 325464 153762
rect 325436 151980 325464 153734
rect 326080 151980 326108 157927
rect 326264 155922 326292 163200
rect 326712 161084 326764 161090
rect 326712 161026 326764 161032
rect 326252 155916 326304 155922
rect 326252 155858 326304 155864
rect 326724 151980 326752 161026
rect 327184 157350 327212 163200
rect 328012 158778 328040 163200
rect 328840 159730 328868 163200
rect 328368 159724 328420 159730
rect 328368 159666 328420 159672
rect 328828 159724 328880 159730
rect 328828 159666 328880 159672
rect 328000 158772 328052 158778
rect 328000 158714 328052 158720
rect 327172 157344 327224 157350
rect 327172 157286 327224 157292
rect 328000 155440 328052 155446
rect 328000 155382 328052 155388
rect 327356 153808 327408 153814
rect 327356 153750 327408 153756
rect 327368 151980 327396 153750
rect 328012 151980 328040 155382
rect 328380 153678 328408 159666
rect 328644 158296 328696 158302
rect 328644 158238 328696 158244
rect 328368 153672 328420 153678
rect 328368 153614 328420 153620
rect 328656 151980 328684 158238
rect 329760 155378 329788 163200
rect 330588 156602 330616 163200
rect 331508 160002 331536 163200
rect 331496 159996 331548 160002
rect 331496 159938 331548 159944
rect 330760 158772 330812 158778
rect 330760 158714 330812 158720
rect 330576 156596 330628 156602
rect 330576 156538 330628 156544
rect 330576 155508 330628 155514
rect 330576 155450 330628 155456
rect 329748 155372 329800 155378
rect 329748 155314 329800 155320
rect 329286 155272 329342 155281
rect 329286 155207 329342 155216
rect 329300 151980 329328 155207
rect 329932 154012 329984 154018
rect 329932 153954 329984 153960
rect 329944 151980 329972 153954
rect 330588 151980 330616 155450
rect 330772 153814 330800 158714
rect 331864 157276 331916 157282
rect 331864 157218 331916 157224
rect 331218 156632 331274 156641
rect 331218 156567 331274 156576
rect 330760 153808 330812 153814
rect 330760 153750 330812 153756
rect 331232 151980 331260 156567
rect 331876 151980 331904 157218
rect 332336 154018 332364 163200
rect 332600 159316 332652 159322
rect 332600 159258 332652 159264
rect 332612 154970 332640 159258
rect 333256 155446 333284 163200
rect 334084 158302 334112 163200
rect 334072 158296 334124 158302
rect 334072 158238 334124 158244
rect 334912 155786 334940 163200
rect 335832 157282 335860 163200
rect 335820 157276 335872 157282
rect 335820 157218 335872 157224
rect 336372 156800 336424 156806
rect 336372 156742 336424 156748
rect 333796 155780 333848 155786
rect 333796 155722 333848 155728
rect 334900 155780 334952 155786
rect 334900 155722 334952 155728
rect 333244 155440 333296 155446
rect 333244 155382 333296 155388
rect 332600 154964 332652 154970
rect 332600 154906 332652 154912
rect 332324 154012 332376 154018
rect 332324 153954 332376 153960
rect 332508 153672 332560 153678
rect 332508 153614 332560 153620
rect 332520 151980 332548 153614
rect 333152 153196 333204 153202
rect 333152 153138 333204 153144
rect 333164 151980 333192 153138
rect 333808 151980 333836 155722
rect 335728 155576 335780 155582
rect 335728 155518 335780 155524
rect 334440 155032 334492 155038
rect 334440 154974 334492 154980
rect 334452 151980 334480 154974
rect 335084 154148 335136 154154
rect 335084 154090 335136 154096
rect 335096 151980 335124 154090
rect 335740 151980 335768 155518
rect 336384 151980 336412 156742
rect 336660 155514 336688 163200
rect 337200 157276 337252 157282
rect 337200 157218 337252 157224
rect 336648 155508 336700 155514
rect 336648 155450 336700 155456
rect 337212 154154 337240 157218
rect 337580 156806 337608 163200
rect 338408 160070 338436 163200
rect 338396 160064 338448 160070
rect 338396 160006 338448 160012
rect 339328 159934 339356 163200
rect 339316 159928 339368 159934
rect 339316 159870 339368 159876
rect 337658 159352 337714 159361
rect 337658 159287 337714 159296
rect 337568 156800 337620 156806
rect 337568 156742 337620 156748
rect 337200 154148 337252 154154
rect 337200 154090 337252 154096
rect 337016 152584 337068 152590
rect 337016 152526 337068 152532
rect 337028 151980 337056 152526
rect 337672 151980 337700 159287
rect 339408 159248 339460 159254
rect 339408 159190 339460 159196
rect 338304 158364 338356 158370
rect 338304 158306 338356 158312
rect 338316 151980 338344 158306
rect 339420 157758 339448 159190
rect 339408 157752 339460 157758
rect 339408 157694 339460 157700
rect 338948 155644 339000 155650
rect 338948 155586 339000 155592
rect 338960 151980 338988 155586
rect 340156 155582 340184 163200
rect 340788 158432 340840 158438
rect 340788 158374 340840 158380
rect 340144 155576 340196 155582
rect 340144 155518 340196 155524
rect 339592 155168 339644 155174
rect 339592 155110 339644 155116
rect 339604 151980 339632 155110
rect 340800 154154 340828 158374
rect 340878 158128 340934 158137
rect 340878 158063 340934 158072
rect 340788 154148 340840 154154
rect 340788 154090 340840 154096
rect 340236 154080 340288 154086
rect 340236 154022 340288 154028
rect 340248 151980 340276 154022
rect 340892 151980 340920 158063
rect 340984 156874 341012 163200
rect 341904 157690 341932 163200
rect 342732 159458 342760 163200
rect 342720 159452 342772 159458
rect 342720 159394 342772 159400
rect 342260 159044 342312 159050
rect 342260 158986 342312 158992
rect 341892 157684 341944 157690
rect 341892 157626 341944 157632
rect 341524 156936 341576 156942
rect 341524 156878 341576 156884
rect 340972 156868 341024 156874
rect 340972 156810 341024 156816
rect 341536 151980 341564 156878
rect 342272 156398 342300 158986
rect 342812 158976 342864 158982
rect 342812 158918 342864 158924
rect 342260 156392 342312 156398
rect 342260 156334 342312 156340
rect 342168 154148 342220 154154
rect 342168 154090 342220 154096
rect 342180 151980 342208 154090
rect 342824 151980 342852 158918
rect 343548 157684 343600 157690
rect 343548 157626 343600 157632
rect 343456 155100 343508 155106
rect 343456 155042 343508 155048
rect 343468 151980 343496 155042
rect 343560 154086 343588 157626
rect 343652 155650 343680 163200
rect 344480 158370 344508 163200
rect 345400 159322 345428 163200
rect 345388 159316 345440 159322
rect 345388 159258 345440 159264
rect 346228 158778 346256 163200
rect 346308 159180 346360 159186
rect 346308 159122 346360 159128
rect 346216 158772 346268 158778
rect 346216 158714 346268 158720
rect 344468 158364 344520 158370
rect 344468 158306 344520 158312
rect 345940 157888 345992 157894
rect 345940 157830 345992 157836
rect 344744 156528 344796 156534
rect 344744 156470 344796 156476
rect 344100 156460 344152 156466
rect 344100 156402 344152 156408
rect 343640 155644 343692 155650
rect 343640 155586 343692 155592
rect 343548 154080 343600 154086
rect 343548 154022 343600 154028
rect 344112 151980 344140 156402
rect 344756 151980 344784 156470
rect 345388 154216 345440 154222
rect 345388 154158 345440 154164
rect 345400 151980 345428 154158
rect 345952 151980 345980 157830
rect 346320 155106 346348 159122
rect 347056 156942 347084 163200
rect 347688 159520 347740 159526
rect 347688 159462 347740 159468
rect 347044 156936 347096 156942
rect 347044 156878 347096 156884
rect 346582 156768 346638 156777
rect 346582 156703 346638 156712
rect 346308 155100 346360 155106
rect 346308 155042 346360 155048
rect 346596 151980 346624 156703
rect 347700 156074 347728 159462
rect 347976 157962 348004 163200
rect 348516 158500 348568 158506
rect 348516 158442 348568 158448
rect 347964 157956 348016 157962
rect 347964 157898 348016 157904
rect 347700 156046 347912 156074
rect 347226 155408 347282 155417
rect 347226 155343 347282 155352
rect 347240 151980 347268 155343
rect 347884 151980 347912 156046
rect 348528 151980 348556 158442
rect 348804 157282 348832 163200
rect 349724 159254 349752 163200
rect 350172 159588 350224 159594
rect 350172 159530 350224 159536
rect 349712 159248 349764 159254
rect 349712 159190 349764 159196
rect 348792 157276 348844 157282
rect 348792 157218 348844 157224
rect 349160 157004 349212 157010
rect 349160 156946 349212 156952
rect 349172 151980 349200 156946
rect 349804 154964 349856 154970
rect 349804 154906 349856 154912
rect 349816 151980 349844 154906
rect 350184 154222 350212 159530
rect 350552 158438 350580 163200
rect 350540 158432 350592 158438
rect 350540 158374 350592 158380
rect 351380 155718 351408 163200
rect 351736 157072 351788 157078
rect 351736 157014 351788 157020
rect 351092 155712 351144 155718
rect 351092 155654 351144 155660
rect 351368 155712 351420 155718
rect 351368 155654 351420 155660
rect 350448 154352 350500 154358
rect 350448 154294 350500 154300
rect 350172 154216 350224 154222
rect 350172 154158 350224 154164
rect 350460 151980 350488 154294
rect 351104 151980 351132 155654
rect 351748 151980 351776 157014
rect 351920 155780 351972 155786
rect 351920 155722 351972 155728
rect 351932 153678 351960 155722
rect 352300 155174 352328 163200
rect 353128 159594 353156 163200
rect 353116 159588 353168 159594
rect 353116 159530 353168 159536
rect 352472 158772 352524 158778
rect 352472 158714 352524 158720
rect 352288 155168 352340 155174
rect 352288 155110 352340 155116
rect 352484 154290 352512 158714
rect 353668 158568 353720 158574
rect 353668 158510 353720 158516
rect 352380 154284 352432 154290
rect 352380 154226 352432 154232
rect 352472 154284 352524 154290
rect 352472 154226 352524 154232
rect 351920 153672 351972 153678
rect 351920 153614 351972 153620
rect 352392 151980 352420 154226
rect 353024 154216 353076 154222
rect 353024 154158 353076 154164
rect 353036 151980 353064 154158
rect 353680 151980 353708 158510
rect 354048 158506 354076 163200
rect 354036 158500 354088 158506
rect 354036 158442 354088 158448
rect 354312 155848 354364 155854
rect 354312 155790 354364 155796
rect 354324 151980 354352 155790
rect 354876 155786 354904 163200
rect 354956 157752 355008 157758
rect 354956 157694 355008 157700
rect 354864 155780 354916 155786
rect 354864 155722 354916 155728
rect 354968 151980 354996 157694
rect 355796 157010 355824 163200
rect 356428 159656 356480 159662
rect 356428 159598 356480 159604
rect 356244 158636 356296 158642
rect 356244 158578 356296 158584
rect 355784 157004 355836 157010
rect 355784 156946 355836 156952
rect 355600 154420 355652 154426
rect 355600 154362 355652 154368
rect 355612 151980 355640 154362
rect 356256 151980 356284 158578
rect 356440 155990 356468 159598
rect 356624 157894 356652 163200
rect 356612 157888 356664 157894
rect 356612 157830 356664 157836
rect 356888 157140 356940 157146
rect 356888 157082 356940 157088
rect 356428 155984 356480 155990
rect 356428 155926 356480 155932
rect 356900 151980 356928 157082
rect 357452 157078 357480 163200
rect 358372 158574 358400 163200
rect 358360 158568 358412 158574
rect 358360 158510 358412 158516
rect 359200 158098 359228 163200
rect 360120 159526 360148 163200
rect 360108 159520 360160 159526
rect 360108 159462 360160 159468
rect 360200 159248 360252 159254
rect 360200 159190 360252 159196
rect 358820 158092 358872 158098
rect 358820 158034 358872 158040
rect 359188 158092 359240 158098
rect 359188 158034 359240 158040
rect 357624 157888 357676 157894
rect 357624 157830 357676 157836
rect 357440 157072 357492 157078
rect 357440 157014 357492 157020
rect 357532 154488 357584 154494
rect 357532 154430 357584 154436
rect 357544 151980 357572 154430
rect 357636 154222 357664 157830
rect 358176 155984 358228 155990
rect 358176 155926 358228 155932
rect 357624 154216 357676 154222
rect 357624 154158 357676 154164
rect 358188 151980 358216 155926
rect 358832 151980 358860 158034
rect 359464 156664 359516 156670
rect 359464 156606 359516 156612
rect 359476 151980 359504 156606
rect 360108 155100 360160 155106
rect 360108 155042 360160 155048
rect 360120 151980 360148 155042
rect 360212 154494 360240 159190
rect 360948 157146 360976 163200
rect 361396 158704 361448 158710
rect 361396 158646 361448 158652
rect 360936 157140 360988 157146
rect 360936 157082 360988 157088
rect 360752 154556 360804 154562
rect 360752 154498 360804 154504
rect 360200 154488 360252 154494
rect 360200 154430 360252 154436
rect 360764 151980 360792 154498
rect 361408 151980 361436 158646
rect 361868 156670 361896 163200
rect 362592 157820 362644 157826
rect 362592 157762 362644 157768
rect 362040 156732 362092 156738
rect 362040 156674 362092 156680
rect 361856 156664 361908 156670
rect 361856 156606 361908 156612
rect 362052 151980 362080 156674
rect 362604 154850 362632 157762
rect 362696 155854 362724 163200
rect 363328 159384 363380 159390
rect 363328 159326 363380 159332
rect 362684 155848 362736 155854
rect 362684 155790 362736 155796
rect 362604 154822 362724 154850
rect 362696 151980 362724 154822
rect 363340 151980 363368 159326
rect 363524 158778 363552 163200
rect 363512 158772 363564 158778
rect 363512 158714 363564 158720
rect 364444 158642 364472 163200
rect 364432 158636 364484 158642
rect 364432 158578 364484 158584
rect 365272 158030 365300 163200
rect 366192 159186 366220 163200
rect 366916 159860 366968 159866
rect 366916 159802 366968 159808
rect 366180 159180 366232 159186
rect 366180 159122 366232 159128
rect 366272 158772 366324 158778
rect 366272 158714 366324 158720
rect 363972 158024 364024 158030
rect 363972 157966 364024 157972
rect 365260 158024 365312 158030
rect 365260 157966 365312 157972
rect 363984 151980 364012 157966
rect 364616 157208 364668 157214
rect 364616 157150 364668 157156
rect 364628 151980 364656 157150
rect 365260 156460 365312 156466
rect 365260 156402 365312 156408
rect 365272 151980 365300 156402
rect 366284 154358 366312 158714
rect 366548 155236 366600 155242
rect 366548 155178 366600 155184
rect 366272 154352 366324 154358
rect 366272 154294 366324 154300
rect 365904 153740 365956 153746
rect 365904 153682 365956 153688
rect 365916 151980 365944 153682
rect 366560 151980 366588 155178
rect 366928 154426 366956 159802
rect 367020 159662 367048 163200
rect 367008 159656 367060 159662
rect 367008 159598 367060 159604
rect 367192 158160 367244 158166
rect 367192 158102 367244 158108
rect 366916 154420 366968 154426
rect 366916 154362 366968 154368
rect 367204 151980 367232 158102
rect 367848 157214 367876 163200
rect 368768 158166 368796 163200
rect 369124 158228 369176 158234
rect 369124 158170 369176 158176
rect 368756 158160 368808 158166
rect 368756 158102 368808 158108
rect 367836 157208 367888 157214
rect 367836 157150 367888 157156
rect 368480 154420 368532 154426
rect 368480 154362 368532 154368
rect 367836 153876 367888 153882
rect 367836 153818 367888 153824
rect 367848 151980 367876 153818
rect 368492 151980 368520 154362
rect 369136 151980 369164 158170
rect 369596 155242 369624 163200
rect 370412 159792 370464 159798
rect 370412 159734 370464 159740
rect 369768 155304 369820 155310
rect 369768 155246 369820 155252
rect 369584 155236 369636 155242
rect 369584 155178 369636 155184
rect 369780 151980 369808 155246
rect 370424 151980 370452 159734
rect 370516 153882 370544 163200
rect 371344 155310 371372 163200
rect 372264 156738 372292 163200
rect 372712 159996 372764 160002
rect 372712 159938 372764 159944
rect 372344 157344 372396 157350
rect 372344 157286 372396 157292
rect 372252 156732 372304 156738
rect 372252 156674 372304 156680
rect 371700 155916 371752 155922
rect 371700 155858 371752 155864
rect 371332 155304 371384 155310
rect 371332 155246 371384 155252
rect 371056 153944 371108 153950
rect 371056 153886 371108 153892
rect 370504 153876 370556 153882
rect 370504 153818 370556 153824
rect 371068 151980 371096 153886
rect 371712 151980 371740 155858
rect 372356 151980 372384 157286
rect 372620 155236 372672 155242
rect 372620 155178 372672 155184
rect 372632 154426 372660 155178
rect 372724 155106 372752 159938
rect 373092 159254 373120 163200
rect 373632 159724 373684 159730
rect 373632 159666 373684 159672
rect 373080 159248 373132 159254
rect 373080 159190 373132 159196
rect 372712 155100 372764 155106
rect 372712 155042 372764 155048
rect 372620 154420 372672 154426
rect 372620 154362 372672 154368
rect 372988 153808 373040 153814
rect 372988 153750 373040 153756
rect 373000 151980 373028 153750
rect 373644 151980 373672 159666
rect 373920 159390 373948 163200
rect 373908 159384 373960 159390
rect 373908 159326 373960 159332
rect 374276 155372 374328 155378
rect 374276 155314 374328 155320
rect 374288 151980 374316 155314
rect 374840 155242 374868 163200
rect 375668 158234 375696 163200
rect 376588 159866 376616 163200
rect 376668 160064 376720 160070
rect 376668 160006 376720 160012
rect 376576 159860 376628 159866
rect 376576 159802 376628 159808
rect 375656 158228 375708 158234
rect 375656 158170 375708 158176
rect 374920 156596 374972 156602
rect 374920 156538 374972 156544
rect 374828 155236 374880 155242
rect 374828 155178 374880 155184
rect 374932 151980 374960 156538
rect 375564 155100 375616 155106
rect 375564 155042 375616 155048
rect 375576 151980 375604 155042
rect 376680 154562 376708 160006
rect 377416 158846 377444 163200
rect 378048 159180 378100 159186
rect 378048 159122 378100 159128
rect 377404 158840 377456 158846
rect 377404 158782 377456 158788
rect 377404 158296 377456 158302
rect 377404 158238 377456 158244
rect 376760 155440 376812 155446
rect 376760 155382 376812 155388
rect 376668 154556 376720 154562
rect 376668 154498 376720 154504
rect 376208 154012 376260 154018
rect 376208 153954 376260 153960
rect 376220 151980 376248 153954
rect 376772 151980 376800 155382
rect 377416 151980 377444 158238
rect 378060 155922 378088 159122
rect 378336 158302 378364 163200
rect 378324 158296 378376 158302
rect 378324 158238 378376 158244
rect 379164 157350 379192 163200
rect 379992 159730 380020 163200
rect 380912 159798 380940 163200
rect 381268 159928 381320 159934
rect 381268 159870 381320 159876
rect 380900 159792 380952 159798
rect 380900 159734 380952 159740
rect 379980 159724 380032 159730
rect 379980 159666 380032 159672
rect 379520 159316 379572 159322
rect 379520 159258 379572 159264
rect 379428 158840 379480 158846
rect 379428 158782 379480 158788
rect 379152 157344 379204 157350
rect 379152 157286 379204 157292
rect 378048 155916 378100 155922
rect 378048 155858 378100 155864
rect 379336 155508 379388 155514
rect 379336 155450 379388 155456
rect 378692 154148 378744 154154
rect 378692 154090 378744 154096
rect 378048 153672 378100 153678
rect 378048 153614 378100 153620
rect 378060 151980 378088 153614
rect 378704 151980 378732 154090
rect 379348 151980 379376 155450
rect 379440 154018 379468 158782
rect 379428 154012 379480 154018
rect 379428 153954 379480 153960
rect 379532 153338 379560 159258
rect 379980 156800 380032 156806
rect 379980 156742 380032 156748
rect 379520 153332 379572 153338
rect 379520 153274 379572 153280
rect 379992 151980 380020 156742
rect 380624 154556 380676 154562
rect 380624 154498 380676 154504
rect 380636 151980 380664 154498
rect 381280 151980 381308 159870
rect 381740 155378 381768 163200
rect 382280 159452 382332 159458
rect 382280 159394 382332 159400
rect 381912 155576 381964 155582
rect 381912 155518 381964 155524
rect 381728 155372 381780 155378
rect 381728 155314 381780 155320
rect 381924 151980 381952 155518
rect 382292 153270 382320 159394
rect 382660 158778 382688 163200
rect 382648 158772 382700 158778
rect 382648 158714 382700 158720
rect 382556 156868 382608 156874
rect 382556 156810 382608 156816
rect 382280 153264 382332 153270
rect 382280 153206 382332 153212
rect 382568 151980 382596 156810
rect 383200 154080 383252 154086
rect 383200 154022 383252 154028
rect 383212 151980 383240 154022
rect 383488 153950 383516 163200
rect 384408 159050 384436 163200
rect 384396 159044 384448 159050
rect 384396 158986 384448 158992
rect 384212 158772 384264 158778
rect 384212 158714 384264 158720
rect 384224 155514 384252 158714
rect 384948 158364 385000 158370
rect 384948 158306 385000 158312
rect 384488 155644 384540 155650
rect 384488 155586 384540 155592
rect 384212 155508 384264 155514
rect 384212 155450 384264 155456
rect 383476 153944 383528 153950
rect 383476 153886 383528 153892
rect 383844 153264 383896 153270
rect 383844 153206 383896 153212
rect 383856 151980 383884 153206
rect 384500 151980 384528 155586
rect 384960 154574 384988 158306
rect 385236 155446 385264 163200
rect 385960 159588 386012 159594
rect 385960 159530 386012 159536
rect 385224 155440 385276 155446
rect 385224 155382 385276 155388
rect 384960 154546 385172 154574
rect 385972 154562 386000 159530
rect 386064 159066 386092 163200
rect 386984 159594 387012 163200
rect 386972 159588 387024 159594
rect 386972 159530 387024 159536
rect 387812 159458 387840 163200
rect 387800 159452 387852 159458
rect 387800 159394 387852 159400
rect 388444 159248 388496 159254
rect 388444 159190 388496 159196
rect 386064 159038 386460 159066
rect 386432 156806 386460 159038
rect 387708 157956 387760 157962
rect 387708 157898 387760 157904
rect 387064 156936 387116 156942
rect 387064 156878 387116 156884
rect 386420 156800 386472 156806
rect 386420 156742 386472 156748
rect 385144 151980 385172 154546
rect 385960 154556 386012 154562
rect 385960 154498 386012 154504
rect 386420 154284 386472 154290
rect 386420 154226 386472 154232
rect 385776 153332 385828 153338
rect 385776 153274 385828 153280
rect 385788 151980 385816 153274
rect 386432 151980 386460 154226
rect 387076 151980 387104 156878
rect 387720 151980 387748 157898
rect 388456 157282 388484 159190
rect 388352 157276 388404 157282
rect 388352 157218 388404 157224
rect 388444 157276 388496 157282
rect 388444 157218 388496 157224
rect 387800 155168 387852 155174
rect 387800 155110 387852 155116
rect 387812 153542 387840 155110
rect 387800 153536 387852 153542
rect 387800 153478 387852 153484
rect 388364 151980 388392 157218
rect 388732 155582 388760 163200
rect 389560 158370 389588 163200
rect 389640 158432 389692 158438
rect 389640 158374 389692 158380
rect 389548 158364 389600 158370
rect 389548 158306 389600 158312
rect 388720 155576 388772 155582
rect 388720 155518 388772 155524
rect 388996 154488 389048 154494
rect 388996 154430 389048 154436
rect 389008 151980 389036 154430
rect 389652 151980 389680 158374
rect 390284 155712 390336 155718
rect 390284 155654 390336 155660
rect 390296 151980 390324 155654
rect 390388 154086 390416 163200
rect 390560 159044 390612 159050
rect 390560 158986 390612 158992
rect 390572 154494 390600 158986
rect 390560 154488 390612 154494
rect 390560 154430 390612 154436
rect 391308 154154 391336 163200
rect 391940 159860 391992 159866
rect 391940 159802 391992 159808
rect 391952 154562 391980 159802
rect 392136 156874 392164 163200
rect 393056 159474 393084 163200
rect 393884 159866 393912 163200
rect 394804 159934 394832 163200
rect 394792 159928 394844 159934
rect 394792 159870 394844 159876
rect 393872 159860 393924 159866
rect 393872 159802 393924 159808
rect 393056 159446 393360 159474
rect 392216 158500 392268 158506
rect 392216 158442 392268 158448
rect 392124 156868 392176 156874
rect 392124 156810 392176 156816
rect 391572 154556 391624 154562
rect 391572 154498 391624 154504
rect 391940 154556 391992 154562
rect 391940 154498 391992 154504
rect 391296 154148 391348 154154
rect 391296 154090 391348 154096
rect 390376 154080 390428 154086
rect 390376 154022 390428 154028
rect 390928 153536 390980 153542
rect 390928 153478 390980 153484
rect 390940 151980 390968 153478
rect 391584 151980 391612 154498
rect 392228 151980 392256 158442
rect 392860 155780 392912 155786
rect 392860 155722 392912 155728
rect 392872 151980 392900 155722
rect 393332 155650 393360 159446
rect 395436 158568 395488 158574
rect 395436 158510 395488 158516
rect 394608 158092 394660 158098
rect 394608 158034 394660 158040
rect 393504 157004 393556 157010
rect 393504 156946 393556 156952
rect 393320 155644 393372 155650
rect 393320 155586 393372 155592
rect 393516 151980 393544 156946
rect 394620 154290 394648 158034
rect 394792 157072 394844 157078
rect 394792 157014 394844 157020
rect 394608 154284 394660 154290
rect 394608 154226 394660 154232
rect 394148 154216 394200 154222
rect 394148 154158 394200 154164
rect 394160 151980 394188 154158
rect 394804 151980 394832 157014
rect 395448 151980 395476 158510
rect 395632 158098 395660 163200
rect 396460 158778 396488 163200
rect 397276 159656 397328 159662
rect 397276 159598 397328 159604
rect 396724 159520 396776 159526
rect 396724 159462 396776 159468
rect 396448 158772 396500 158778
rect 396448 158714 396500 158720
rect 395620 158092 395672 158098
rect 395620 158034 395672 158040
rect 396080 154284 396132 154290
rect 396080 154226 396132 154232
rect 396092 151980 396120 154226
rect 396736 151980 396764 159462
rect 397288 155990 397316 159598
rect 397380 158794 397408 163200
rect 398208 158846 398236 163200
rect 398196 158840 398248 158846
rect 397380 158766 397500 158794
rect 398196 158782 398248 158788
rect 397368 157140 397420 157146
rect 397368 157082 397420 157088
rect 397276 155984 397328 155990
rect 397276 155926 397328 155932
rect 397380 151980 397408 157082
rect 397472 154222 397500 158766
rect 399128 156670 399156 163200
rect 399956 159746 399984 163200
rect 399956 159718 400260 159746
rect 399392 158840 399444 158846
rect 399392 158782 399444 158788
rect 398012 156664 398064 156670
rect 398012 156606 398064 156612
rect 399116 156664 399168 156670
rect 399116 156606 399168 156612
rect 397460 154216 397512 154222
rect 397460 154158 397512 154164
rect 398024 151980 398052 156606
rect 398656 155848 398708 155854
rect 398656 155790 398708 155796
rect 398668 151980 398696 155790
rect 399404 154358 399432 158782
rect 399944 158636 399996 158642
rect 399944 158578 399996 158584
rect 399300 154352 399352 154358
rect 399300 154294 399352 154300
rect 399392 154352 399444 154358
rect 399392 154294 399444 154300
rect 399312 151980 399340 154294
rect 399956 151980 399984 158578
rect 400232 158030 400260 159718
rect 400876 159526 400904 163200
rect 401704 159662 401732 163200
rect 401692 159656 401744 159662
rect 401692 159598 401744 159604
rect 400864 159520 400916 159526
rect 400864 159462 400916 159468
rect 400220 158024 400272 158030
rect 400220 157966 400272 157972
rect 400588 157956 400640 157962
rect 400588 157898 400640 157904
rect 400600 151980 400628 157898
rect 402428 157208 402480 157214
rect 402428 157150 402480 157156
rect 401876 155984 401928 155990
rect 401876 155926 401928 155932
rect 401232 155916 401284 155922
rect 401232 155858 401284 155864
rect 401244 151980 401272 155858
rect 401888 151980 401916 155926
rect 402440 154578 402468 157150
rect 402532 156942 402560 163200
rect 403452 158846 403480 163200
rect 403440 158840 403492 158846
rect 403440 158782 403492 158788
rect 403164 158160 403216 158166
rect 403164 158102 403216 158108
rect 402520 156936 402572 156942
rect 402520 156878 402572 156884
rect 402440 154550 402560 154578
rect 402532 151980 402560 154550
rect 403176 151980 403204 158102
rect 403808 154420 403860 154426
rect 403808 154362 403860 154368
rect 403820 151980 403848 154362
rect 404280 154290 404308 163200
rect 405096 155304 405148 155310
rect 405096 155246 405148 155252
rect 404268 154284 404320 154290
rect 404268 154226 404320 154232
rect 404452 153876 404504 153882
rect 404452 153818 404504 153824
rect 404464 151980 404492 153818
rect 405108 151980 405136 155246
rect 405200 153814 405228 163200
rect 405648 158840 405700 158846
rect 405648 158782 405700 158788
rect 405660 155718 405688 158782
rect 406028 158166 406056 163200
rect 406752 159384 406804 159390
rect 406752 159326 406804 159332
rect 406016 158160 406068 158166
rect 406016 158102 406068 158108
rect 406384 157276 406436 157282
rect 406384 157218 406436 157224
rect 405740 156732 405792 156738
rect 405740 156674 405792 156680
rect 405648 155712 405700 155718
rect 405648 155654 405700 155660
rect 405188 153808 405240 153814
rect 405188 153750 405240 153756
rect 405752 151980 405780 156674
rect 406396 151980 406424 157218
rect 406764 155666 406792 159326
rect 406856 158794 406884 163200
rect 407776 159390 407804 163200
rect 408604 160002 408632 163200
rect 408592 159996 408644 160002
rect 408592 159938 408644 159944
rect 407764 159384 407816 159390
rect 407764 159326 407816 159332
rect 406856 158766 407160 158794
rect 406764 155638 407068 155666
rect 407040 151980 407068 155638
rect 407132 155310 407160 158766
rect 408224 158228 408276 158234
rect 408224 158170 408276 158176
rect 407120 155304 407172 155310
rect 407120 155246 407172 155252
rect 407580 155236 407632 155242
rect 407580 155178 407632 155184
rect 407592 151980 407620 155178
rect 408236 151980 408264 158170
rect 408500 157344 408552 157350
rect 408500 157286 408552 157292
rect 408512 153882 408540 157286
rect 409524 155242 409552 163200
rect 410156 158296 410208 158302
rect 410156 158238 410208 158244
rect 409512 155236 409564 155242
rect 409512 155178 409564 155184
rect 408868 154556 408920 154562
rect 408868 154498 408920 154504
rect 408500 153876 408552 153882
rect 408500 153818 408552 153824
rect 408880 151980 408908 154498
rect 409512 154012 409564 154018
rect 409512 153954 409564 153960
rect 409524 151980 409552 153954
rect 410168 151980 410196 158238
rect 410352 157010 410380 163200
rect 411168 159724 411220 159730
rect 411168 159666 411220 159672
rect 410340 157004 410392 157010
rect 410340 156946 410392 156952
rect 411180 153898 411208 159666
rect 411272 154018 411300 163200
rect 411996 159792 412048 159798
rect 411996 159734 412048 159740
rect 412008 155802 412036 159734
rect 412100 159730 412128 163200
rect 412088 159724 412140 159730
rect 412088 159666 412140 159672
rect 412008 155774 412128 155802
rect 411260 154012 411312 154018
rect 411260 153954 411312 153960
rect 410800 153876 410852 153882
rect 411180 153870 411484 153898
rect 410800 153818 410852 153824
rect 410812 151980 410840 153818
rect 411456 151980 411484 153870
rect 412100 151980 412128 155774
rect 412928 155378 412956 163200
rect 413848 155786 413876 163200
rect 414676 161474 414704 163200
rect 414676 161446 414796 161474
rect 413836 155780 413888 155786
rect 413836 155722 413888 155728
rect 413376 155508 413428 155514
rect 413376 155450 413428 155456
rect 412732 155372 412784 155378
rect 412732 155314 412784 155320
rect 412916 155372 412968 155378
rect 412916 155314 412968 155320
rect 412744 151980 412772 155314
rect 413388 151980 413416 155450
rect 414664 154488 414716 154494
rect 414664 154430 414716 154436
rect 414020 153944 414072 153950
rect 414020 153886 414072 153892
rect 414032 151980 414060 153886
rect 414676 151980 414704 154430
rect 414768 153950 414796 161446
rect 415216 159588 415268 159594
rect 415216 159530 415268 159536
rect 414756 153944 414808 153950
rect 414756 153886 414808 153892
rect 415228 153746 415256 159530
rect 415308 155440 415360 155446
rect 415308 155382 415360 155388
rect 415216 153740 415268 153746
rect 415216 153682 415268 153688
rect 415320 151980 415348 155382
rect 415596 154426 415624 163200
rect 415952 156800 416004 156806
rect 415952 156742 416004 156748
rect 415584 154420 415636 154426
rect 415584 154362 415636 154368
rect 415964 151980 415992 156742
rect 416424 155446 416452 163200
rect 417240 159452 417292 159458
rect 417240 159394 417292 159400
rect 416412 155440 416464 155446
rect 416412 155382 416464 155388
rect 416596 153740 416648 153746
rect 416596 153682 416648 153688
rect 416608 151980 416636 153682
rect 417252 151980 417280 159394
rect 417344 156738 417372 163200
rect 418172 160070 418200 163200
rect 419000 163146 419028 163200
rect 419092 163146 419120 163254
rect 419000 163118 419120 163146
rect 418160 160064 418212 160070
rect 418160 160006 418212 160012
rect 418528 158364 418580 158370
rect 418528 158306 418580 158312
rect 417332 156732 417384 156738
rect 417332 156674 417384 156680
rect 417884 155576 417936 155582
rect 417884 155518 417936 155524
rect 417896 151980 417924 155518
rect 418540 151980 418568 158306
rect 419276 154086 419304 163254
rect 419906 163200 419962 164000
rect 420734 163200 420790 164000
rect 421654 163200 421710 164000
rect 422482 163200 422538 164000
rect 423402 163200 423458 164000
rect 424230 163200 424286 164000
rect 425058 163200 425114 164000
rect 425978 163200 426034 164000
rect 426806 163200 426862 164000
rect 427726 163200 427782 164000
rect 428554 163200 428610 164000
rect 429382 163200 429438 164000
rect 430302 163200 430358 164000
rect 431130 163200 431186 164000
rect 432050 163200 432106 164000
rect 432878 163200 432934 164000
rect 432984 163254 433288 163282
rect 419920 155582 419948 163200
rect 420460 156868 420512 156874
rect 420460 156810 420512 156816
rect 419908 155576 419960 155582
rect 419908 155518 419960 155524
rect 419816 154148 419868 154154
rect 419816 154090 419868 154096
rect 419172 154080 419224 154086
rect 419172 154022 419224 154028
rect 419264 154080 419316 154086
rect 419264 154022 419316 154028
rect 419184 151980 419212 154022
rect 419828 151980 419856 154090
rect 420472 151980 420500 156810
rect 420748 156806 420776 163200
rect 420920 159928 420972 159934
rect 420920 159870 420972 159876
rect 420736 156800 420788 156806
rect 420736 156742 420788 156748
rect 420932 153270 420960 159870
rect 421668 159594 421696 163200
rect 421748 159860 421800 159866
rect 421748 159802 421800 159808
rect 421656 159588 421708 159594
rect 421656 159530 421708 159536
rect 421104 155644 421156 155650
rect 421104 155586 421156 155592
rect 420920 153264 420972 153270
rect 420920 153206 420972 153212
rect 421116 151980 421144 155586
rect 421760 151980 421788 159802
rect 422496 154154 422524 163200
rect 423416 158098 423444 163200
rect 423680 158432 423732 158438
rect 423680 158374 423732 158380
rect 423036 158092 423088 158098
rect 423036 158034 423088 158040
rect 423404 158092 423456 158098
rect 423404 158034 423456 158040
rect 422484 154148 422536 154154
rect 422484 154090 422536 154096
rect 422392 153264 422444 153270
rect 422392 153206 422444 153212
rect 422404 151980 422432 153206
rect 423048 151980 423076 158034
rect 423692 151980 423720 158374
rect 424244 155650 424272 163200
rect 424232 155644 424284 155650
rect 424232 155586 424284 155592
rect 424968 154352 425020 154358
rect 424968 154294 425020 154300
rect 424324 154216 424376 154222
rect 424324 154158 424376 154164
rect 424336 151980 424364 154158
rect 424980 151980 425008 154294
rect 425072 154222 425100 163200
rect 425992 159798 426020 163200
rect 425980 159792 426032 159798
rect 425980 159734 426032 159740
rect 426820 158846 426848 163200
rect 427544 159656 427596 159662
rect 427544 159598 427596 159604
rect 426900 159520 426952 159526
rect 426900 159462 426952 159468
rect 426808 158840 426860 158846
rect 426808 158782 426860 158788
rect 426256 158024 426308 158030
rect 426256 157966 426308 157972
rect 425612 156664 425664 156670
rect 425612 156606 425664 156612
rect 425060 154216 425112 154222
rect 425060 154158 425112 154164
rect 425624 151980 425652 156606
rect 426268 151980 426296 157966
rect 426912 151980 426940 159462
rect 427556 151980 427584 159598
rect 427740 158778 427768 163200
rect 427728 158772 427780 158778
rect 427728 158714 427780 158720
rect 428188 156936 428240 156942
rect 428188 156878 428240 156884
rect 428200 151980 428228 156878
rect 428568 154358 428596 163200
rect 429396 159526 429424 163200
rect 429384 159520 429436 159526
rect 429384 159462 429436 159468
rect 429384 158840 429436 158846
rect 429384 158782 429436 158788
rect 429200 157004 429252 157010
rect 429200 156946 429252 156952
rect 428832 155712 428884 155718
rect 428832 155654 428884 155660
rect 428556 154352 428608 154358
rect 428556 154294 428608 154300
rect 428844 151980 428872 155654
rect 429212 153270 429240 156946
rect 429396 155786 429424 158782
rect 429384 155780 429436 155786
rect 429384 155722 429436 155728
rect 430316 155718 430344 163200
rect 431144 159662 431172 163200
rect 432064 159866 432092 163200
rect 432892 163146 432920 163200
rect 432984 163146 433012 163254
rect 432892 163118 433012 163146
rect 432696 159996 432748 160002
rect 432696 159938 432748 159944
rect 432052 159860 432104 159866
rect 432052 159802 432104 159808
rect 431132 159656 431184 159662
rect 431132 159598 431184 159604
rect 432052 159384 432104 159390
rect 432052 159326 432104 159332
rect 430580 158772 430632 158778
rect 430580 158714 430632 158720
rect 430592 155922 430620 158714
rect 430764 158160 430816 158166
rect 430764 158102 430816 158108
rect 430580 155916 430632 155922
rect 430580 155858 430632 155864
rect 430304 155712 430356 155718
rect 430304 155654 430356 155660
rect 429476 154284 429528 154290
rect 429476 154226 429528 154232
rect 429200 153264 429252 153270
rect 429200 153206 429252 153212
rect 429488 151980 429516 154226
rect 430120 153876 430172 153882
rect 430120 153818 430172 153824
rect 430132 151980 430160 153818
rect 430776 151980 430804 158102
rect 431408 155304 431460 155310
rect 431408 155246 431460 155252
rect 431420 151980 431448 155246
rect 432064 151980 432092 159326
rect 432708 151980 432736 159938
rect 433260 153882 433288 163254
rect 433798 163200 433854 164000
rect 434626 163200 434682 164000
rect 435454 163200 435510 164000
rect 436374 163200 436430 164000
rect 437202 163200 437258 164000
rect 438122 163200 438178 164000
rect 438950 163200 439006 164000
rect 439870 163200 439926 164000
rect 440698 163200 440754 164000
rect 441526 163200 441582 164000
rect 442446 163200 442502 164000
rect 443274 163200 443330 164000
rect 444194 163200 444250 164000
rect 445022 163200 445078 164000
rect 445850 163200 445906 164000
rect 446770 163200 446826 164000
rect 447598 163200 447654 164000
rect 448518 163200 448574 164000
rect 449346 163200 449402 164000
rect 450266 163200 450322 164000
rect 451094 163200 451150 164000
rect 451922 163200 451978 164000
rect 452842 163200 452898 164000
rect 453670 163200 453726 164000
rect 454590 163200 454646 164000
rect 455418 163200 455474 164000
rect 456338 163200 456394 164000
rect 457166 163200 457222 164000
rect 457994 163200 458050 164000
rect 458914 163200 458970 164000
rect 459742 163200 459798 164000
rect 460662 163200 460718 164000
rect 461490 163200 461546 164000
rect 462410 163200 462466 164000
rect 463238 163200 463294 164000
rect 464066 163200 464122 164000
rect 464986 163200 465042 164000
rect 465814 163200 465870 164000
rect 466734 163200 466790 164000
rect 467562 163200 467618 164000
rect 468390 163200 468446 164000
rect 469310 163200 469366 164000
rect 470138 163200 470194 164000
rect 471058 163200 471114 164000
rect 471886 163200 471942 164000
rect 472806 163200 472862 164000
rect 473634 163200 473690 164000
rect 474462 163200 474518 164000
rect 475382 163200 475438 164000
rect 476210 163200 476266 164000
rect 477130 163200 477186 164000
rect 477958 163200 478014 164000
rect 478878 163200 478934 164000
rect 479706 163200 479762 164000
rect 480534 163200 480590 164000
rect 481454 163200 481510 164000
rect 482282 163200 482338 164000
rect 483202 163200 483258 164000
rect 484030 163200 484086 164000
rect 484858 163200 484914 164000
rect 485778 163200 485834 164000
rect 486606 163200 486662 164000
rect 487526 163200 487582 164000
rect 488354 163200 488410 164000
rect 489274 163200 489330 164000
rect 490102 163200 490158 164000
rect 490930 163200 490986 164000
rect 491036 163254 491248 163282
rect 433812 155242 433840 163200
rect 434640 156670 434668 163200
rect 435272 159724 435324 159730
rect 435272 159666 435324 159672
rect 434628 156664 434680 156670
rect 434628 156606 434680 156612
rect 433340 155236 433392 155242
rect 433340 155178 433392 155184
rect 433800 155236 433852 155242
rect 433800 155178 433852 155184
rect 433248 153876 433300 153882
rect 433248 153818 433300 153824
rect 433352 151980 433380 155178
rect 434628 154012 434680 154018
rect 434628 153954 434680 153960
rect 433984 153264 434036 153270
rect 433984 153206 434036 153212
rect 433996 151980 434024 153206
rect 434640 151980 434668 153954
rect 435284 151980 435312 159666
rect 435468 158982 435496 163200
rect 436008 159860 436060 159866
rect 436008 159802 436060 159808
rect 435456 158976 435508 158982
rect 435456 158918 435508 158924
rect 435916 155508 435968 155514
rect 435916 155450 435968 155456
rect 435928 151980 435956 155450
rect 436020 154290 436048 159802
rect 436008 154284 436060 154290
rect 436008 154226 436060 154232
rect 436388 154018 436416 163200
rect 436560 155372 436612 155378
rect 436560 155314 436612 155320
rect 436376 154012 436428 154018
rect 436376 153954 436428 153960
rect 436572 151980 436600 155314
rect 437216 155310 437244 163200
rect 437480 159656 437532 159662
rect 437480 159598 437532 159604
rect 437492 155854 437520 159598
rect 437480 155848 437532 155854
rect 437480 155790 437532 155796
rect 438136 155378 438164 163200
rect 438964 156874 438992 163200
rect 439688 160064 439740 160070
rect 439688 160006 439740 160012
rect 438952 156868 439004 156874
rect 438952 156810 439004 156816
rect 439044 156732 439096 156738
rect 439044 156674 439096 156680
rect 438400 155440 438452 155446
rect 438400 155382 438452 155388
rect 438124 155372 438176 155378
rect 438124 155314 438176 155320
rect 437204 155304 437256 155310
rect 437204 155246 437256 155252
rect 437848 154420 437900 154426
rect 437848 154362 437900 154368
rect 437204 153944 437256 153950
rect 437204 153886 437256 153892
rect 437216 151980 437244 153886
rect 437860 151980 437888 154362
rect 438412 151980 438440 155382
rect 439056 151980 439084 156674
rect 439700 151980 439728 160006
rect 439884 159458 439912 163200
rect 439872 159452 439924 159458
rect 439872 159394 439924 159400
rect 440240 156800 440292 156806
rect 440240 156742 440292 156748
rect 440252 153270 440280 156742
rect 440712 155446 440740 163200
rect 441540 156738 441568 163200
rect 442460 159662 442488 163200
rect 442448 159656 442500 159662
rect 442448 159598 442500 159604
rect 442264 159588 442316 159594
rect 442264 159530 442316 159536
rect 441528 156732 441580 156738
rect 441528 156674 441580 156680
rect 440976 155576 441028 155582
rect 440976 155518 441028 155524
rect 440700 155440 440752 155446
rect 440700 155382 440752 155388
rect 440332 154080 440384 154086
rect 440332 154022 440384 154028
rect 440240 153264 440292 153270
rect 440240 153206 440292 153212
rect 440344 151980 440372 154022
rect 440988 151980 441016 155518
rect 441620 153264 441672 153270
rect 441620 153206 441672 153212
rect 441632 151980 441660 153206
rect 442276 151980 442304 159530
rect 442816 158976 442868 158982
rect 442816 158918 442868 158924
rect 442828 154086 442856 158918
rect 443288 158030 443316 163200
rect 444208 159118 444236 163200
rect 444196 159112 444248 159118
rect 444196 159054 444248 159060
rect 445036 158778 445064 163200
rect 445864 160002 445892 163200
rect 445852 159996 445904 160002
rect 445852 159938 445904 159944
rect 445484 159792 445536 159798
rect 445484 159734 445536 159740
rect 445024 158772 445076 158778
rect 445024 158714 445076 158720
rect 443552 158092 443604 158098
rect 443552 158034 443604 158040
rect 443276 158024 443328 158030
rect 443276 157966 443328 157972
rect 442908 154148 442960 154154
rect 442908 154090 442960 154096
rect 442816 154080 442868 154086
rect 442816 154022 442868 154028
rect 442920 151980 442948 154090
rect 443564 151980 443592 158034
rect 444196 155644 444248 155650
rect 444196 155586 444248 155592
rect 444208 151980 444236 155586
rect 444840 154216 444892 154222
rect 444840 154158 444892 154164
rect 444852 151980 444880 154158
rect 445496 151980 445524 159734
rect 445668 159656 445720 159662
rect 445668 159598 445720 159604
rect 445680 155514 445708 159598
rect 446404 159452 446456 159458
rect 446404 159394 446456 159400
rect 446416 155786 446444 159394
rect 446784 158846 446812 163200
rect 447612 159662 447640 163200
rect 448532 159730 448560 163200
rect 448520 159724 448572 159730
rect 448520 159666 448572 159672
rect 447600 159656 447652 159662
rect 447600 159598 447652 159604
rect 449360 159594 449388 163200
rect 450280 159866 450308 163200
rect 451108 159934 451136 163200
rect 451096 159928 451148 159934
rect 451096 159870 451148 159876
rect 450268 159860 450320 159866
rect 450268 159802 450320 159808
rect 451936 159798 451964 163200
rect 452856 160070 452884 163200
rect 452844 160064 452896 160070
rect 452844 160006 452896 160012
rect 451924 159792 451976 159798
rect 451924 159734 451976 159740
rect 449348 159588 449400 159594
rect 449348 159530 449400 159536
rect 446864 159520 446916 159526
rect 446864 159462 446916 159468
rect 446772 158840 446824 158846
rect 446772 158782 446824 158788
rect 446876 155922 446904 159462
rect 453684 159390 453712 163200
rect 454604 159458 454632 163200
rect 454592 159452 454644 159458
rect 454592 159394 454644 159400
rect 453672 159384 453724 159390
rect 453672 159326 453724 159332
rect 455432 159254 455460 163200
rect 456352 159322 456380 163200
rect 456892 159996 456944 160002
rect 456892 159938 456944 159944
rect 456340 159316 456392 159322
rect 456340 159258 456392 159264
rect 455420 159248 455472 159254
rect 455420 159190 455472 159196
rect 447232 159112 447284 159118
rect 447232 159054 447284 159060
rect 447140 158772 447192 158778
rect 447140 158714 447192 158720
rect 446772 155916 446824 155922
rect 446772 155858 446824 155864
rect 446864 155916 446916 155922
rect 446864 155858 446916 155864
rect 446128 155780 446180 155786
rect 446128 155722 446180 155728
rect 446404 155780 446456 155786
rect 446404 155722 446456 155728
rect 445668 155508 445720 155514
rect 445668 155450 445720 155456
rect 446140 151980 446168 155722
rect 446784 151980 446812 155858
rect 447152 155582 447180 158714
rect 447244 155650 447272 159054
rect 451740 158840 451792 158846
rect 451740 158782 451792 158788
rect 449900 156664 449952 156670
rect 449900 156606 449952 156612
rect 448060 155916 448112 155922
rect 448060 155858 448112 155864
rect 447232 155644 447284 155650
rect 447232 155586 447284 155592
rect 447140 155576 447192 155582
rect 447140 155518 447192 155524
rect 447416 154352 447468 154358
rect 447416 154294 447468 154300
rect 447428 151980 447456 154294
rect 448072 151980 448100 155858
rect 449348 155848 449400 155854
rect 449348 155790 449400 155796
rect 448704 155712 448756 155718
rect 448704 155654 448756 155660
rect 448716 151980 448744 155654
rect 449360 151980 449388 155790
rect 449912 153270 449940 156606
rect 451280 155236 451332 155242
rect 451280 155178 451332 155184
rect 449992 154012 450044 154018
rect 449992 153954 450044 153960
rect 449900 153264 449952 153270
rect 449900 153206 449952 153212
rect 450004 151980 450032 153954
rect 450636 153876 450688 153882
rect 450636 153818 450688 153824
rect 450648 151980 450676 153818
rect 451292 151980 451320 155178
rect 451752 153882 451780 158782
rect 455144 156868 455196 156874
rect 455144 156810 455196 156816
rect 454500 155372 454552 155378
rect 454500 155314 454552 155320
rect 453856 155304 453908 155310
rect 453856 155246 453908 155252
rect 452568 154080 452620 154086
rect 452568 154022 452620 154028
rect 451740 153876 451792 153882
rect 451740 153818 451792 153824
rect 451924 153264 451976 153270
rect 451924 153206 451976 153212
rect 451936 151980 451964 153206
rect 452580 151980 452608 154022
rect 453212 153944 453264 153950
rect 453212 153886 453264 153892
rect 453224 151980 453252 153886
rect 453868 151980 453896 155246
rect 454512 151980 454540 155314
rect 455156 151980 455184 156810
rect 455788 155780 455840 155786
rect 455788 155722 455840 155728
rect 455800 151980 455828 155722
rect 456432 155440 456484 155446
rect 456432 155382 456484 155388
rect 456444 151980 456472 155382
rect 456904 154562 456932 159938
rect 457180 159186 457208 163200
rect 458008 159594 458036 163200
rect 458928 160002 458956 163200
rect 458916 159996 458968 160002
rect 458916 159938 458968 159944
rect 458180 159656 458232 159662
rect 458180 159598 458232 159604
rect 457996 159588 458048 159594
rect 457996 159530 458048 159536
rect 457168 159180 457220 159186
rect 457168 159122 457220 159128
rect 457076 156732 457128 156738
rect 457076 156674 457128 156680
rect 456892 154556 456944 154562
rect 456892 154498 456944 154504
rect 457088 151980 457116 156674
rect 457720 155508 457772 155514
rect 457720 155450 457772 155456
rect 457732 151980 457760 155450
rect 458192 153270 458220 159598
rect 459560 159520 459612 159526
rect 459560 159462 459612 159468
rect 458364 158024 458416 158030
rect 458364 157966 458416 157972
rect 458180 153264 458232 153270
rect 458180 153206 458232 153212
rect 458376 151980 458404 157966
rect 459008 155644 459060 155650
rect 459008 155586 459060 155592
rect 459020 151980 459048 155586
rect 459572 153406 459600 159462
rect 459756 159050 459784 163200
rect 459836 159724 459888 159730
rect 459836 159666 459888 159672
rect 459744 159044 459796 159050
rect 459744 158986 459796 158992
rect 459652 155576 459704 155582
rect 459652 155518 459704 155524
rect 459560 153400 459612 153406
rect 459560 153342 459612 153348
rect 459664 151980 459692 155518
rect 459848 153338 459876 159666
rect 460676 159662 460704 163200
rect 460664 159656 460716 159662
rect 460664 159598 460716 159604
rect 461504 158846 461532 163200
rect 462136 159928 462188 159934
rect 462136 159870 462188 159876
rect 461492 158840 461544 158846
rect 461492 158782 461544 158788
rect 460296 154556 460348 154562
rect 460296 154498 460348 154504
rect 459836 153332 459888 153338
rect 459836 153274 459888 153280
rect 460308 151980 460336 154498
rect 462148 154154 462176 159870
rect 462228 159860 462280 159866
rect 462228 159802 462280 159808
rect 462240 154562 462268 159802
rect 462424 159526 462452 163200
rect 462872 159792 462924 159798
rect 462872 159734 462924 159740
rect 462412 159520 462464 159526
rect 462412 159462 462464 159468
rect 462228 154556 462280 154562
rect 462228 154498 462280 154504
rect 462136 154148 462188 154154
rect 462136 154090 462188 154096
rect 460940 153876 460992 153882
rect 460940 153818 460992 153824
rect 460952 151980 460980 153818
rect 462884 153610 462912 159734
rect 463252 158914 463280 163200
rect 463792 160064 463844 160070
rect 463792 160006 463844 160012
rect 463700 159384 463752 159390
rect 463700 159326 463752 159332
rect 463240 158908 463292 158914
rect 463240 158850 463292 158856
rect 463516 154556 463568 154562
rect 463516 154498 463568 154504
rect 462872 153604 462924 153610
rect 462872 153546 462924 153552
rect 462872 153400 462924 153406
rect 462872 153342 462924 153348
rect 462228 153332 462280 153338
rect 462228 153274 462280 153280
rect 461584 153264 461636 153270
rect 461584 153206 461636 153212
rect 461596 151980 461624 153206
rect 462240 151980 462268 153274
rect 462884 151980 462912 153342
rect 463528 151980 463556 154498
rect 463712 153882 463740 159326
rect 463700 153876 463752 153882
rect 463700 153818 463752 153824
rect 463804 153474 463832 160006
rect 464080 159118 464108 163200
rect 464068 159112 464120 159118
rect 464068 159054 464120 159060
rect 465000 158778 465028 163200
rect 465828 159798 465856 163200
rect 465816 159792 465868 159798
rect 465816 159734 465868 159740
rect 466368 159452 466420 159458
rect 466368 159394 466420 159400
rect 465632 159044 465684 159050
rect 465632 158986 465684 158992
rect 464988 158772 465040 158778
rect 464988 158714 465040 158720
rect 465644 154290 465672 158986
rect 466380 154574 466408 159394
rect 466748 158982 466776 163200
rect 467380 159248 467432 159254
rect 467380 159190 467432 159196
rect 466736 158976 466788 158982
rect 466736 158918 466788 158924
rect 466828 158840 466880 158846
rect 466828 158782 466880 158788
rect 466380 154546 466776 154574
rect 465632 154284 465684 154290
rect 465632 154226 465684 154232
rect 464160 154148 464212 154154
rect 464160 154090 464212 154096
rect 463792 153468 463844 153474
rect 463792 153410 463844 153416
rect 464172 151980 464200 154090
rect 466092 153876 466144 153882
rect 466092 153818 466144 153824
rect 464804 153604 464856 153610
rect 464804 153546 464856 153552
rect 464816 151980 464844 153546
rect 465448 153468 465500 153474
rect 465448 153410 465500 153416
rect 465460 151980 465488 153410
rect 466104 151980 466132 153818
rect 466748 151980 466776 154546
rect 466840 153474 466868 158782
rect 466828 153468 466880 153474
rect 466828 153410 466880 153416
rect 467392 151980 467420 159190
rect 467576 158846 467604 163200
rect 468404 159934 468432 163200
rect 468392 159928 468444 159934
rect 468392 159870 468444 159876
rect 469324 159594 469352 163200
rect 469864 159996 469916 160002
rect 469864 159938 469916 159944
rect 469128 159588 469180 159594
rect 469128 159530 469180 159536
rect 469312 159588 469364 159594
rect 469312 159530 469364 159536
rect 468208 159520 468260 159526
rect 468208 159462 468260 159468
rect 467748 159316 467800 159322
rect 467748 159258 467800 159264
rect 467564 158840 467616 158846
rect 467564 158782 467616 158788
rect 467760 154574 467788 159258
rect 468116 158908 468168 158914
rect 468116 158850 468168 158856
rect 467760 154546 468064 154574
rect 468036 151980 468064 154546
rect 468128 153406 468156 158850
rect 468116 153400 468168 153406
rect 468116 153342 468168 153348
rect 468220 153338 468248 159462
rect 468668 159180 468720 159186
rect 468668 159122 468720 159128
rect 468208 153332 468260 153338
rect 468208 153274 468260 153280
rect 468680 151980 468708 159122
rect 469140 153762 469168 159530
rect 469312 159112 469364 159118
rect 469312 159054 469364 159060
rect 469220 158772 469272 158778
rect 469220 158714 469272 158720
rect 469232 153882 469260 158714
rect 469324 154086 469352 159054
rect 469312 154080 469364 154086
rect 469312 154022 469364 154028
rect 469220 153876 469272 153882
rect 469220 153818 469272 153824
rect 469140 153734 469260 153762
rect 469232 151980 469260 153734
rect 469876 151980 469904 159938
rect 470152 159866 470180 163200
rect 470140 159860 470192 159866
rect 470140 159802 470192 159808
rect 471072 159050 471100 163200
rect 471900 159934 471928 163200
rect 471888 159928 471940 159934
rect 471888 159870 471940 159876
rect 471888 159792 471940 159798
rect 471888 159734 471940 159740
rect 471152 159656 471204 159662
rect 471152 159598 471204 159604
rect 471060 159044 471112 159050
rect 471060 158986 471112 158992
rect 470508 154284 470560 154290
rect 470508 154226 470560 154232
rect 470520 151980 470548 154226
rect 471164 151980 471192 159598
rect 471900 154426 471928 159734
rect 472820 158914 472848 163200
rect 473648 159390 473676 163200
rect 473728 159860 473780 159866
rect 473728 159802 473780 159808
rect 473636 159384 473688 159390
rect 473636 159326 473688 159332
rect 473268 158976 473320 158982
rect 473268 158918 473320 158924
rect 472808 158908 472860 158914
rect 472808 158850 472860 158856
rect 473176 158840 473228 158846
rect 473176 158782 473228 158788
rect 471888 154420 471940 154426
rect 471888 154362 471940 154368
rect 473188 154154 473216 158782
rect 473280 154562 473308 158918
rect 473268 154556 473320 154562
rect 473268 154498 473320 154504
rect 473740 154290 473768 159802
rect 474476 159118 474504 163200
rect 475396 160002 475424 163200
rect 475384 159996 475436 160002
rect 475384 159938 475436 159944
rect 476120 159928 476172 159934
rect 476120 159870 476172 159876
rect 475752 159724 475804 159730
rect 475752 159666 475804 159672
rect 474740 159588 474792 159594
rect 474740 159530 474792 159536
rect 474464 159112 474516 159118
rect 474464 159054 474516 159060
rect 473728 154284 473780 154290
rect 473728 154226 473780 154232
rect 473176 154148 473228 154154
rect 473176 154090 473228 154096
rect 473728 154080 473780 154086
rect 473728 154022 473780 154028
rect 471796 153468 471848 153474
rect 471796 153410 471848 153416
rect 471808 151980 471836 153410
rect 473084 153400 473136 153406
rect 473084 153342 473136 153348
rect 472440 153332 472492 153338
rect 472440 153274 472492 153280
rect 472452 151980 472480 153274
rect 473096 151980 473124 153342
rect 473740 151980 473768 154022
rect 474752 154018 474780 159530
rect 475764 154562 475792 159666
rect 475660 154556 475712 154562
rect 475660 154498 475712 154504
rect 475752 154556 475804 154562
rect 475752 154498 475804 154504
rect 475016 154420 475068 154426
rect 475016 154362 475068 154368
rect 474740 154012 474792 154018
rect 474740 153954 474792 153960
rect 474372 153876 474424 153882
rect 474372 153818 474424 153824
rect 474384 151980 474412 153818
rect 475028 151980 475056 154362
rect 475672 151980 475700 154498
rect 476132 154426 476160 159870
rect 476224 158778 476252 163200
rect 476396 159044 476448 159050
rect 476396 158986 476448 158992
rect 476212 158772 476264 158778
rect 476212 158714 476264 158720
rect 476120 154420 476172 154426
rect 476120 154362 476172 154368
rect 476304 154148 476356 154154
rect 476304 154090 476356 154096
rect 476316 151980 476344 154090
rect 476408 153270 476436 158986
rect 477144 158846 477172 163200
rect 477972 159934 478000 163200
rect 477960 159928 478012 159934
rect 477960 159870 478012 159876
rect 478892 159798 478920 163200
rect 478880 159792 478932 159798
rect 478880 159734 478932 159740
rect 479720 159526 479748 163200
rect 479708 159520 479760 159526
rect 479708 159462 479760 159468
rect 478972 159384 479024 159390
rect 478972 159326 479024 159332
rect 478880 159112 478932 159118
rect 478880 159054 478932 159060
rect 477500 158908 477552 158914
rect 477500 158850 477552 158856
rect 477132 158840 477184 158846
rect 477132 158782 477184 158788
rect 477512 154290 477540 158850
rect 478236 154556 478288 154562
rect 478236 154498 478288 154504
rect 476948 154284 477000 154290
rect 476948 154226 477000 154232
rect 477500 154284 477552 154290
rect 477500 154226 477552 154232
rect 476396 153264 476448 153270
rect 476396 153206 476448 153212
rect 476960 151980 476988 154226
rect 477592 154012 477644 154018
rect 477592 153954 477644 153960
rect 477604 151980 477632 153954
rect 478248 151980 478276 154498
rect 478892 153338 478920 159054
rect 478880 153332 478932 153338
rect 478880 153274 478932 153280
rect 478984 153270 479012 159326
rect 480548 159050 480576 163200
rect 481088 159996 481140 160002
rect 481088 159938 481140 159944
rect 480536 159044 480588 159050
rect 480536 158986 480588 158992
rect 479524 154420 479576 154426
rect 479524 154362 479576 154368
rect 478972 153264 479024 153270
rect 478972 153206 479024 153212
rect 478880 153196 478932 153202
rect 478880 153138 478932 153144
rect 478892 151980 478920 153138
rect 479536 151980 479564 154362
rect 480168 154284 480220 154290
rect 480168 154226 480220 154232
rect 480180 151980 480208 154226
rect 481100 153610 481128 159938
rect 481468 158982 481496 163200
rect 481456 158976 481508 158982
rect 481456 158918 481508 158924
rect 482296 158914 482324 163200
rect 482284 158908 482336 158914
rect 482284 158850 482336 158856
rect 482008 158840 482060 158846
rect 482008 158782 482060 158788
rect 482020 154018 482048 158782
rect 483216 158778 483244 163200
rect 484044 160070 484072 163200
rect 484032 160064 484084 160070
rect 484032 160006 484084 160012
rect 484032 159928 484084 159934
rect 484032 159870 484084 159876
rect 482744 158772 482796 158778
rect 482744 158714 482796 158720
rect 483204 158772 483256 158778
rect 483204 158714 483256 158720
rect 482008 154012 482060 154018
rect 482008 153954 482060 153960
rect 481088 153604 481140 153610
rect 481088 153546 481140 153552
rect 482100 153604 482152 153610
rect 482100 153546 482152 153552
rect 481456 153332 481508 153338
rect 481456 153274 481508 153280
rect 480812 153264 480864 153270
rect 480812 153206 480864 153212
rect 480824 151980 480852 153206
rect 481468 151980 481496 153274
rect 482112 151980 482140 153546
rect 482756 151980 482784 158714
rect 483388 154012 483440 154018
rect 483388 153954 483440 153960
rect 483400 151980 483428 153954
rect 484044 151980 484072 159870
rect 484676 159792 484728 159798
rect 484676 159734 484728 159740
rect 484688 151980 484716 159734
rect 484872 158846 484900 163200
rect 485320 159520 485372 159526
rect 485320 159462 485372 159468
rect 484860 158840 484912 158846
rect 484860 158782 484912 158788
rect 485332 151980 485360 159462
rect 485792 158778 485820 163200
rect 486620 160070 486648 163200
rect 486608 160064 486660 160070
rect 486608 160006 486660 160012
rect 485964 159044 486016 159050
rect 485964 158986 486016 158992
rect 485504 158772 485556 158778
rect 485504 158714 485556 158720
rect 485780 158772 485832 158778
rect 485780 158714 485832 158720
rect 485516 154154 485544 158714
rect 485504 154148 485556 154154
rect 485504 154090 485556 154096
rect 485976 151980 486004 158986
rect 487540 158982 487568 163200
rect 488264 160064 488316 160070
rect 488264 160006 488316 160012
rect 486608 158976 486660 158982
rect 486608 158918 486660 158924
rect 487528 158976 487580 158982
rect 487528 158918 487580 158924
rect 486620 151980 486648 158918
rect 487252 158908 487304 158914
rect 487252 158850 487304 158856
rect 486976 158840 487028 158846
rect 486976 158782 487028 158788
rect 486988 154494 487016 158782
rect 486976 154488 487028 154494
rect 486976 154430 487028 154436
rect 487264 151980 487292 158850
rect 487804 158772 487856 158778
rect 487804 158714 487856 158720
rect 487816 154562 487844 158714
rect 487804 154556 487856 154562
rect 487804 154498 487856 154504
rect 487896 154148 487948 154154
rect 487896 154090 487948 154096
rect 487908 151980 487936 154090
rect 488276 153474 488304 160006
rect 488368 158794 488396 163200
rect 488724 159996 488776 160002
rect 488724 159938 488776 159944
rect 488632 158976 488684 158982
rect 488632 158918 488684 158924
rect 488368 158766 488580 158794
rect 488264 153468 488316 153474
rect 488264 153410 488316 153416
rect 488552 153406 488580 158766
rect 488540 153400 488592 153406
rect 488540 153342 488592 153348
rect 488644 153270 488672 158918
rect 488632 153264 488684 153270
rect 488632 153206 488684 153212
rect 488736 153082 488764 159938
rect 489288 158914 489316 163200
rect 489276 158908 489328 158914
rect 489276 158850 489328 158856
rect 490116 158778 490144 163200
rect 490944 163146 490972 163200
rect 491036 163146 491064 163254
rect 490944 163118 491064 163146
rect 491220 159066 491248 163254
rect 491850 163200 491906 164000
rect 492678 163200 492734 164000
rect 493598 163200 493654 164000
rect 494426 163200 494482 164000
rect 495346 163200 495402 164000
rect 496174 163200 496230 164000
rect 497002 163200 497058 164000
rect 497922 163200 497978 164000
rect 498750 163200 498806 164000
rect 499670 163200 499726 164000
rect 499776 163254 500080 163282
rect 491220 159038 491340 159066
rect 491208 158908 491260 158914
rect 491208 158850 491260 158856
rect 490104 158772 490156 158778
rect 490104 158714 490156 158720
rect 489828 154556 489880 154562
rect 489828 154498 489880 154504
rect 489184 154488 489236 154494
rect 489184 154430 489236 154436
rect 488552 153054 488764 153082
rect 488552 151980 488580 153054
rect 489196 151980 489224 154430
rect 489840 151980 489868 154498
rect 491220 154154 491248 158850
rect 491312 154290 491340 159038
rect 491864 158846 491892 163200
rect 492692 158914 492720 163200
rect 492680 158908 492732 158914
rect 492680 158850 492732 158856
rect 491852 158840 491904 158846
rect 491852 158782 491904 158788
rect 493612 158778 493640 163200
rect 494440 158846 494468 163200
rect 494980 158908 495032 158914
rect 494980 158850 495032 158856
rect 493968 158840 494020 158846
rect 493968 158782 494020 158788
rect 494428 158840 494480 158846
rect 494428 158782 494480 158788
rect 491576 158772 491628 158778
rect 491576 158714 491628 158720
rect 493600 158772 493652 158778
rect 493600 158714 493652 158720
rect 491588 154562 491616 158714
rect 491576 154556 491628 154562
rect 491576 154498 491628 154504
rect 493048 154556 493100 154562
rect 493980 154544 494008 158782
rect 493980 154516 494376 154544
rect 493048 154498 493100 154504
rect 491300 154284 491352 154290
rect 491300 154226 491352 154232
rect 491208 154148 491260 154154
rect 491208 154090 491260 154096
rect 492404 154148 492456 154154
rect 492404 154090 492456 154096
rect 490472 153468 490524 153474
rect 490472 153410 490524 153416
rect 490484 151980 490512 153410
rect 491760 153400 491812 153406
rect 491760 153342 491812 153348
rect 491116 153264 491168 153270
rect 491116 153206 491168 153212
rect 491128 151980 491156 153206
rect 491772 151980 491800 153342
rect 492416 151980 492444 154090
rect 493060 151980 493088 154498
rect 493692 154284 493744 154290
rect 493692 154226 493744 154232
rect 493704 151980 493732 154226
rect 494348 151980 494376 154516
rect 494992 151980 495020 158850
rect 495360 158794 495388 163200
rect 495256 158772 495308 158778
rect 495360 158766 495480 158794
rect 496188 158778 496216 163200
rect 497016 158846 497044 163200
rect 496268 158840 496320 158846
rect 496268 158782 496320 158788
rect 497004 158840 497056 158846
rect 497004 158782 497056 158788
rect 495256 158714 495308 158720
rect 495268 154442 495296 158714
rect 495452 154562 495480 158766
rect 496176 158772 496228 158778
rect 496176 158714 496228 158720
rect 495440 154556 495492 154562
rect 495440 154498 495492 154504
rect 495268 154414 495664 154442
rect 495636 151980 495664 154414
rect 496280 151980 496308 158782
rect 497936 158778 497964 163200
rect 498200 158840 498252 158846
rect 498200 158782 498252 158788
rect 497556 158772 497608 158778
rect 497556 158714 497608 158720
rect 497924 158772 497976 158778
rect 497924 158714 497976 158720
rect 496912 154556 496964 154562
rect 496912 154498 496964 154504
rect 496924 151980 496952 154498
rect 497568 151980 497596 158714
rect 498212 151980 498240 158782
rect 498764 154562 498792 163200
rect 499684 163146 499712 163200
rect 499776 163146 499804 163254
rect 499684 163118 499804 163146
rect 498844 158772 498896 158778
rect 498844 158714 498896 158720
rect 498752 154556 498804 154562
rect 498752 154498 498804 154504
rect 498856 151980 498884 158714
rect 499488 154556 499540 154562
rect 499488 154498 499540 154504
rect 499500 151980 499528 154498
rect 500052 151980 500080 163254
rect 500498 163200 500554 164000
rect 501418 163200 501474 164000
rect 501984 163254 502196 163282
rect 500512 161474 500540 163200
rect 501432 161474 501460 163200
rect 500512 161446 500724 161474
rect 500696 151980 500724 161446
rect 501340 161446 501460 161474
rect 501340 151980 501368 161446
rect 501984 151980 502012 163254
rect 502168 163146 502196 163254
rect 502246 163200 502302 164000
rect 502628 163254 503024 163282
rect 502260 163146 502288 163200
rect 502168 163118 502288 163146
rect 502628 151980 502656 163254
rect 502996 163146 503024 163254
rect 503074 163200 503130 164000
rect 503732 163254 503944 163282
rect 503088 163146 503116 163200
rect 502996 163118 503116 163146
rect 503732 158778 503760 163254
rect 503916 163146 503944 163254
rect 503994 163200 504050 164000
rect 504822 163200 504878 164000
rect 505742 163200 505798 164000
rect 506570 163200 506626 164000
rect 507398 163200 507454 164000
rect 508318 163200 508374 164000
rect 509146 163200 509202 164000
rect 510066 163200 510122 164000
rect 510894 163200 510950 164000
rect 511814 163200 511870 164000
rect 512642 163200 512698 164000
rect 513470 163200 513526 164000
rect 514390 163200 514446 164000
rect 514772 163254 515168 163282
rect 504008 163146 504036 163200
rect 503916 163118 504036 163146
rect 504548 158840 504600 158846
rect 504548 158782 504600 158788
rect 503260 158772 503312 158778
rect 503260 158714 503312 158720
rect 503720 158772 503772 158778
rect 503720 158714 503772 158720
rect 503904 158772 503956 158778
rect 503904 158714 503956 158720
rect 503272 151980 503300 158714
rect 503916 151980 503944 158714
rect 504560 151980 504588 158782
rect 504836 158778 504864 163200
rect 505756 158846 505784 163200
rect 506480 158908 506532 158914
rect 506480 158850 506532 158856
rect 505744 158840 505796 158846
rect 505744 158782 505796 158788
rect 505836 158840 505888 158846
rect 505836 158782 505888 158788
rect 504824 158772 504876 158778
rect 504824 158714 504876 158720
rect 505192 158772 505244 158778
rect 505192 158714 505244 158720
rect 505204 151980 505232 158714
rect 505848 151980 505876 158782
rect 506492 151980 506520 158850
rect 506584 158778 506612 163200
rect 507124 158976 507176 158982
rect 507124 158918 507176 158924
rect 506572 158772 506624 158778
rect 506572 158714 506624 158720
rect 507136 151980 507164 158918
rect 507412 158846 507440 163200
rect 508332 158914 508360 163200
rect 509160 158982 509188 163200
rect 509148 158976 509200 158982
rect 509148 158918 509200 158924
rect 509700 158976 509752 158982
rect 509700 158918 509752 158924
rect 508320 158908 508372 158914
rect 508320 158850 508372 158856
rect 508412 158908 508464 158914
rect 508412 158850 508464 158856
rect 507400 158840 507452 158846
rect 507400 158782 507452 158788
rect 507768 158840 507820 158846
rect 507768 158782 507820 158788
rect 507780 151980 507808 158782
rect 508424 151980 508452 158850
rect 509056 158772 509108 158778
rect 509056 158714 509108 158720
rect 509068 151980 509096 158714
rect 509712 151980 509740 158918
rect 510080 158846 510108 163200
rect 510908 158914 510936 163200
rect 510896 158908 510948 158914
rect 510896 158850 510948 158856
rect 510068 158840 510120 158846
rect 510068 158782 510120 158788
rect 510988 158840 511040 158846
rect 510988 158782 511040 158788
rect 510344 154488 510396 154494
rect 510344 154430 510396 154436
rect 510356 151980 510384 154430
rect 511000 151980 511028 158782
rect 511828 158778 511856 163200
rect 512656 158982 512684 163200
rect 512644 158976 512696 158982
rect 512644 158918 512696 158924
rect 511816 158772 511868 158778
rect 511816 158714 511868 158720
rect 512276 154556 512328 154562
rect 512276 154498 512328 154504
rect 511632 154284 511684 154290
rect 511632 154226 511684 154232
rect 511644 151980 511672 154226
rect 512288 151980 512316 154498
rect 513484 154494 513512 163200
rect 514404 158846 514432 163200
rect 514392 158840 514444 158846
rect 514392 158782 514444 158788
rect 513472 154488 513524 154494
rect 513472 154430 513524 154436
rect 513564 154488 513616 154494
rect 513564 154430 513616 154436
rect 512920 154420 512972 154426
rect 512920 154362 512972 154368
rect 512932 151980 512960 154362
rect 513576 151980 513604 154430
rect 514208 154352 514260 154358
rect 514208 154294 514260 154300
rect 514220 151980 514248 154294
rect 514772 154290 514800 163254
rect 515140 163146 515168 163254
rect 515218 163200 515274 164000
rect 516138 163200 516194 164000
rect 516966 163200 517022 164000
rect 517624 163254 517836 163282
rect 515232 163146 515260 163200
rect 515140 163118 515260 163146
rect 516152 154562 516180 163200
rect 516140 154556 516192 154562
rect 516140 154498 516192 154504
rect 516980 154426 517008 163200
rect 517624 154494 517652 163254
rect 517808 163146 517836 163254
rect 517886 163200 517942 164000
rect 518714 163200 518770 164000
rect 518912 163254 519492 163282
rect 517900 163146 517928 163200
rect 517808 163118 517928 163146
rect 517612 154488 517664 154494
rect 517612 154430 517664 154436
rect 518728 154426 518756 163200
rect 516968 154420 517020 154426
rect 516968 154362 517020 154368
rect 518716 154420 518768 154426
rect 518716 154362 518768 154368
rect 518072 154352 518124 154358
rect 518072 154294 518124 154300
rect 514760 154284 514812 154290
rect 514760 154226 514812 154232
rect 517428 154148 517480 154154
rect 517428 154090 517480 154096
rect 515496 153604 515548 153610
rect 515496 153546 515548 153552
rect 514852 153468 514904 153474
rect 514852 153410 514904 153416
rect 514864 151980 514892 153410
rect 515508 151980 515536 153546
rect 516140 153400 516192 153406
rect 516140 153342 516192 153348
rect 516152 151980 516180 153342
rect 516784 153264 516836 153270
rect 516784 153206 516836 153212
rect 516796 151980 516824 153206
rect 517440 151980 517468 154090
rect 518084 151980 518112 154294
rect 518716 154216 518768 154222
rect 518716 154158 518768 154164
rect 518728 151980 518756 154158
rect 518912 153474 518940 163254
rect 519464 163146 519492 163254
rect 519542 163200 519598 164000
rect 520462 163200 520518 164000
rect 520752 163254 521240 163282
rect 519556 163146 519584 163200
rect 519464 163118 519584 163146
rect 520476 161474 520504 163200
rect 520292 161446 520504 161474
rect 520292 158794 520320 161446
rect 520200 158766 520320 158794
rect 520556 158840 520608 158846
rect 520556 158782 520608 158788
rect 520004 154556 520056 154562
rect 520004 154498 520056 154504
rect 519360 154420 519412 154426
rect 519360 154362 519412 154368
rect 518900 153468 518952 153474
rect 518900 153410 518952 153416
rect 519372 151980 519400 154362
rect 520016 151980 520044 154498
rect 520200 153610 520228 158766
rect 520188 153604 520240 153610
rect 520188 153546 520240 153552
rect 520568 153270 520596 158782
rect 520648 153604 520700 153610
rect 520648 153546 520700 153552
rect 520556 153264 520608 153270
rect 520556 153206 520608 153212
rect 520660 151980 520688 153546
rect 520752 153406 520780 163254
rect 521212 163146 521240 163254
rect 521290 163200 521346 164000
rect 522210 163200 522266 164000
rect 523038 163200 523094 164000
rect 523866 163200 523922 164000
rect 524786 163200 524842 164000
rect 525614 163200 525670 164000
rect 525812 163254 526484 163282
rect 521304 163146 521332 163200
rect 521212 163118 521332 163146
rect 522224 158846 522252 163200
rect 522212 158840 522264 158846
rect 522212 158782 522264 158788
rect 521660 158772 521712 158778
rect 521660 158714 521712 158720
rect 521292 154488 521344 154494
rect 521292 154430 521344 154436
rect 520740 153400 520792 153406
rect 520740 153342 520792 153348
rect 521304 151980 521332 154430
rect 521672 154358 521700 158714
rect 521660 154352 521712 154358
rect 521660 154294 521712 154300
rect 523052 154154 523080 163200
rect 523132 158840 523184 158846
rect 523132 158782 523184 158788
rect 523144 154426 523172 158782
rect 523880 158778 523908 163200
rect 523868 158772 523920 158778
rect 523868 158714 523920 158720
rect 523132 154420 523184 154426
rect 523132 154362 523184 154368
rect 524512 154420 524564 154426
rect 524512 154362 524564 154368
rect 523040 154148 523092 154154
rect 523040 154090 523092 154096
rect 523868 154148 523920 154154
rect 523868 154090 523920 154096
rect 523224 154080 523276 154086
rect 523224 154022 523276 154028
rect 522580 153400 522632 153406
rect 522580 153342 522632 153348
rect 521936 153332 521988 153338
rect 521936 153274 521988 153280
rect 521948 151980 521976 153274
rect 522592 151980 522620 153342
rect 523236 151980 523264 154022
rect 523880 151980 523908 154090
rect 524524 151980 524552 154362
rect 524800 154222 524828 163200
rect 525628 158846 525656 163200
rect 525616 158840 525668 158846
rect 525616 158782 525668 158788
rect 525812 154562 525840 163254
rect 526456 163146 526484 163254
rect 526534 163200 526590 164000
rect 527362 163200 527418 164000
rect 528282 163200 528338 164000
rect 528572 163254 529060 163282
rect 526548 163146 526576 163200
rect 526456 163118 526576 163146
rect 527180 158772 527232 158778
rect 527180 158714 527232 158720
rect 525800 154556 525852 154562
rect 525800 154498 525852 154504
rect 525800 154352 525852 154358
rect 525800 154294 525852 154300
rect 525156 154284 525208 154290
rect 525156 154226 525208 154232
rect 524788 154216 524840 154222
rect 524788 154158 524840 154164
rect 525168 151980 525196 154226
rect 525812 151980 525840 154294
rect 526444 154216 526496 154222
rect 526444 154158 526496 154164
rect 526456 151980 526484 154158
rect 527192 154086 527220 158714
rect 527180 154080 527232 154086
rect 527180 154022 527232 154028
rect 527088 153876 527140 153882
rect 527088 153818 527140 153824
rect 527100 151980 527128 153818
rect 527376 153610 527404 163200
rect 527732 154556 527784 154562
rect 527732 154498 527784 154504
rect 527364 153604 527416 153610
rect 527364 153546 527416 153552
rect 527744 151980 527772 154498
rect 528296 154494 528324 163200
rect 528284 154488 528336 154494
rect 528284 154430 528336 154436
rect 528376 154488 528428 154494
rect 528376 154430 528428 154436
rect 528388 151980 528416 154430
rect 528572 153338 528600 163254
rect 529032 163146 529060 163254
rect 529110 163200 529166 164000
rect 529938 163200 529994 164000
rect 530858 163200 530914 164000
rect 531332 163254 531636 163282
rect 529124 163146 529152 163200
rect 529032 163118 529152 163146
rect 529664 154012 529716 154018
rect 529664 153954 529716 153960
rect 529020 153944 529072 153950
rect 529020 153886 529072 153892
rect 528560 153332 528612 153338
rect 528560 153274 528612 153280
rect 529032 151980 529060 153886
rect 529676 151980 529704 153954
rect 529952 153406 529980 163200
rect 530872 158778 530900 163200
rect 530860 158772 530912 158778
rect 530860 158714 530912 158720
rect 531332 154154 531360 163254
rect 531608 163146 531636 163254
rect 531686 163200 531742 164000
rect 531792 163254 532556 163282
rect 531700 163146 531728 163200
rect 531608 163118 531728 163146
rect 531412 158772 531464 158778
rect 531412 158714 531464 158720
rect 531424 154290 531452 158714
rect 531792 154426 531820 163254
rect 532528 163146 532556 163254
rect 532606 163200 532662 164000
rect 533434 163200 533490 164000
rect 534092 163254 534304 163282
rect 532620 163146 532648 163200
rect 532528 163118 532648 163146
rect 533160 158976 533212 158982
rect 533160 158918 533212 158924
rect 532700 158908 532752 158914
rect 532700 158850 532752 158856
rect 531964 157412 532016 157418
rect 531964 157354 532016 157360
rect 531780 154420 531832 154426
rect 531780 154362 531832 154368
rect 531412 154284 531464 154290
rect 531412 154226 531464 154232
rect 531320 154148 531372 154154
rect 531320 154090 531372 154096
rect 529940 153400 529992 153406
rect 529940 153342 529992 153348
rect 531596 151564 531648 151570
rect 531596 151506 531648 151512
rect 531608 151201 531636 151506
rect 531594 151192 531650 151201
rect 127624 151156 127676 151162
rect 531594 151127 531650 151136
rect 127624 151098 127676 151104
rect 126978 150920 127034 150929
rect 126978 150855 127034 150864
rect 126992 150686 127020 150855
rect 126980 150680 127032 150686
rect 126980 150622 127032 150628
rect 126704 150476 126756 150482
rect 126704 150418 126756 150424
rect 126980 149048 127032 149054
rect 126978 149016 126980 149025
rect 127032 149016 127034 149025
rect 126978 148951 127034 148960
rect 126980 147620 127032 147626
rect 126980 147562 127032 147568
rect 126992 147121 127020 147562
rect 126978 147112 127034 147121
rect 126978 147047 127034 147056
rect 126980 146260 127032 146266
rect 126980 146202 127032 146208
rect 126992 145217 127020 146202
rect 126978 145208 127034 145217
rect 126978 145143 127034 145152
rect 126980 143540 127032 143546
rect 126980 143482 127032 143488
rect 126992 143313 127020 143482
rect 126978 143304 127034 143313
rect 126978 143239 127034 143248
rect 126980 140752 127032 140758
rect 126980 140694 127032 140700
rect 126992 139505 127020 140694
rect 126978 139496 127034 139505
rect 126978 139431 127034 139440
rect 126980 137964 127032 137970
rect 126980 137906 127032 137912
rect 126992 137465 127020 137906
rect 126978 137456 127034 137465
rect 126978 137391 127034 137400
rect 126980 136604 127032 136610
rect 126980 136546 127032 136552
rect 126992 135561 127020 136546
rect 126978 135552 127034 135561
rect 126978 135487 127034 135496
rect 126980 133884 127032 133890
rect 126980 133826 127032 133832
rect 126992 133657 127020 133826
rect 126978 133648 127034 133657
rect 126978 133583 127034 133592
rect 126980 132456 127032 132462
rect 126980 132398 127032 132404
rect 126992 131753 127020 132398
rect 126978 131744 127034 131753
rect 126978 131679 127034 131688
rect 126980 131096 127032 131102
rect 126980 131038 127032 131044
rect 126992 129849 127020 131038
rect 126978 129840 127034 129849
rect 126978 129775 127034 129784
rect 126980 128308 127032 128314
rect 126980 128250 127032 128256
rect 126992 127945 127020 128250
rect 126978 127936 127034 127945
rect 126978 127871 127034 127880
rect 126980 126948 127032 126954
rect 126980 126890 127032 126896
rect 126992 126041 127020 126890
rect 126978 126032 127034 126041
rect 126978 125967 127034 125976
rect 126334 124128 126390 124137
rect 126334 124063 126390 124072
rect 126980 122460 127032 122466
rect 126980 122402 127032 122408
rect 126992 122097 127020 122402
rect 126978 122088 127034 122097
rect 126978 122023 127034 122032
rect 126980 121440 127032 121446
rect 126980 121382 127032 121388
rect 126992 120193 127020 121382
rect 126978 120184 127034 120193
rect 126978 120119 127034 120128
rect 126980 118652 127032 118658
rect 126980 118594 127032 118600
rect 126992 118289 127020 118594
rect 126978 118280 127034 118289
rect 126978 118215 127034 118224
rect 126980 117292 127032 117298
rect 126980 117234 127032 117240
rect 126992 116385 127020 117234
rect 126978 116376 127034 116385
rect 126978 116311 127034 116320
rect 126980 113144 127032 113150
rect 126980 113086 127032 113092
rect 126992 112577 127020 113086
rect 126978 112568 127034 112577
rect 126978 112503 127034 112512
rect 126980 111784 127032 111790
rect 126980 111726 127032 111732
rect 126992 110673 127020 111726
rect 126978 110664 127034 110673
rect 126978 110599 127034 110608
rect 126980 108996 127032 109002
rect 126980 108938 127032 108944
rect 126992 108769 127020 108938
rect 126978 108760 127034 108769
rect 126978 108695 127034 108704
rect 126980 107636 127032 107642
rect 126980 107578 127032 107584
rect 126992 106729 127020 107578
rect 126978 106720 127034 106729
rect 126978 106655 127034 106664
rect 126980 104848 127032 104854
rect 126978 104816 126980 104825
rect 127032 104816 127034 104825
rect 126978 104751 127034 104760
rect 126980 103488 127032 103494
rect 126980 103430 127032 103436
rect 126992 102921 127020 103430
rect 126978 102912 127034 102921
rect 126978 102847 127034 102856
rect 126980 102128 127032 102134
rect 126980 102070 127032 102076
rect 126992 101017 127020 102070
rect 126978 101008 127034 101017
rect 126978 100943 127034 100952
rect 126980 99340 127032 99346
rect 126980 99282 127032 99288
rect 126992 99113 127020 99282
rect 126978 99104 127034 99113
rect 126978 99039 127034 99048
rect 126980 97980 127032 97986
rect 126980 97922 127032 97928
rect 126992 97209 127020 97922
rect 126978 97200 127034 97209
rect 126978 97135 127034 97144
rect 126980 96620 127032 96626
rect 126980 96562 127032 96568
rect 126992 95305 127020 96562
rect 126978 95296 127034 95305
rect 126978 95231 127034 95240
rect 126242 93256 126298 93265
rect 126242 93191 126298 93200
rect 127636 91361 127664 151098
rect 127900 150476 127952 150482
rect 127900 150418 127952 150424
rect 127716 149728 127768 149734
rect 127716 149670 127768 149676
rect 127728 114481 127756 149670
rect 127912 141409 127940 150418
rect 531976 147121 532004 157354
rect 532712 154222 532740 158850
rect 532792 158840 532844 158846
rect 532792 158782 532844 158788
rect 532804 154562 532832 158782
rect 532792 154556 532844 154562
rect 532792 154498 532844 154504
rect 533172 154494 533200 158918
rect 533448 158778 533476 163200
rect 534092 158794 534120 163254
rect 534276 163146 534304 163254
rect 534354 163200 534410 164000
rect 535182 163200 535238 164000
rect 535564 163254 535960 163282
rect 534368 163146 534396 163200
rect 534276 163118 534396 163146
rect 534722 163160 534778 163169
rect 534722 163095 534778 163104
rect 533436 158772 533488 158778
rect 533436 158714 533488 158720
rect 534000 158766 534120 158794
rect 533160 154488 533212 154494
rect 533160 154430 533212 154436
rect 534000 154358 534028 158766
rect 533988 154352 534040 154358
rect 533988 154294 534040 154300
rect 532700 154216 532752 154222
rect 532700 154158 532752 154164
rect 534736 151570 534764 163095
rect 535196 158914 535224 163200
rect 535184 158908 535236 158914
rect 535184 158850 535236 158856
rect 535458 158672 535514 158681
rect 535458 158607 535514 158616
rect 535472 157418 535500 158607
rect 535460 157412 535512 157418
rect 535460 157354 535512 157360
rect 535366 157176 535422 157185
rect 535366 157111 535422 157120
rect 535274 154048 535330 154057
rect 535274 153983 535330 153992
rect 534906 152552 534962 152561
rect 534906 152487 534962 152496
rect 534724 151564 534776 151570
rect 534724 151506 534776 151512
rect 532608 149932 532660 149938
rect 532608 149874 532660 149880
rect 532620 149841 532648 149874
rect 532606 149832 532662 149841
rect 532606 149767 532662 149776
rect 534722 149560 534778 149569
rect 534722 149495 534778 149504
rect 532332 149048 532384 149054
rect 532332 148990 532384 148996
rect 532344 148481 532372 148990
rect 532330 148472 532386 148481
rect 532330 148407 532386 148416
rect 531962 147112 532018 147121
rect 531962 147047 532018 147056
rect 532148 146124 532200 146130
rect 532148 146066 532200 146072
rect 532160 145761 532188 146066
rect 532146 145752 532202 145761
rect 532146 145687 532202 145696
rect 531780 144900 531832 144906
rect 531780 144842 531832 144848
rect 531792 144401 531820 144842
rect 531778 144392 531834 144401
rect 531778 144327 531834 144336
rect 531688 143268 531740 143274
rect 531688 143210 531740 143216
rect 531700 143041 531728 143210
rect 531686 143032 531742 143041
rect 531686 142967 531742 142976
rect 531964 141908 532016 141914
rect 531964 141850 532016 141856
rect 531976 141681 532004 141850
rect 531962 141672 532018 141681
rect 531962 141607 532018 141616
rect 127898 141400 127954 141409
rect 127898 141335 127954 141344
rect 531964 140752 532016 140758
rect 531964 140694 532016 140700
rect 531976 140321 532004 140694
rect 531962 140312 532018 140321
rect 531962 140247 532018 140256
rect 534736 139398 534764 149495
rect 534814 148064 534870 148073
rect 534814 147999 534870 148008
rect 531596 139392 531648 139398
rect 531596 139334 531648 139340
rect 534724 139392 534776 139398
rect 534724 139334 534776 139340
rect 531608 138961 531636 139334
rect 531594 138952 531650 138961
rect 531594 138887 531650 138896
rect 534828 137970 534856 147999
rect 534920 141914 534948 152487
rect 535182 151056 535238 151065
rect 535182 150991 535238 151000
rect 535090 146568 535146 146577
rect 535090 146503 535146 146512
rect 534998 144936 535054 144945
rect 534998 144871 535054 144880
rect 534908 141908 534960 141914
rect 534908 141850 534960 141856
rect 531412 137964 531464 137970
rect 531412 137906 531464 137912
rect 534816 137964 534868 137970
rect 534816 137906 534868 137912
rect 531424 137601 531452 137906
rect 531410 137592 531466 137601
rect 531410 137527 531466 137536
rect 532148 136400 532200 136406
rect 532148 136342 532200 136348
rect 532160 136241 532188 136342
rect 532146 136232 532202 136241
rect 532146 136167 532202 136176
rect 535012 134910 535040 144871
rect 535104 136406 535132 146503
rect 535196 140758 535224 150991
rect 535288 143274 535316 153983
rect 535380 146130 535408 157111
rect 535564 153882 535592 163254
rect 535932 163146 535960 163254
rect 536010 163200 536066 164000
rect 536930 163200 536986 164000
rect 537758 163200 537814 164000
rect 538678 163200 538734 164000
rect 539506 163200 539562 164000
rect 536024 163146 536052 163200
rect 535932 163118 536052 163146
rect 536102 161664 536158 161673
rect 536102 161599 536158 161608
rect 535552 153876 535604 153882
rect 535552 153818 535604 153824
rect 536116 149938 536144 161599
rect 536194 160168 536250 160177
rect 536194 160103 536250 160112
rect 536104 149932 536156 149938
rect 536104 149874 536156 149880
rect 536208 149054 536236 160103
rect 536944 158846 536972 163200
rect 537772 158982 537800 163200
rect 537760 158976 537812 158982
rect 537760 158918 537812 158924
rect 536932 158840 536984 158846
rect 536932 158782 536984 158788
rect 538692 158778 538720 163200
rect 539520 158778 539548 163200
rect 538680 158772 538732 158778
rect 538680 158714 538732 158720
rect 539508 158772 539560 158778
rect 539508 158714 539560 158720
rect 536286 155680 536342 155689
rect 536286 155615 536342 155624
rect 536196 149048 536248 149054
rect 536196 148990 536248 148996
rect 535368 146124 535420 146130
rect 535368 146066 535420 146072
rect 536300 144906 536328 155615
rect 536288 144900 536340 144906
rect 536288 144842 536340 144848
rect 536194 143440 536250 143449
rect 536194 143375 536250 143384
rect 535276 143268 535328 143274
rect 535276 143210 535328 143216
rect 536010 141944 536066 141953
rect 536010 141879 536066 141888
rect 535184 140752 535236 140758
rect 535184 140694 535236 140700
rect 535092 136400 535144 136406
rect 535092 136342 535144 136348
rect 531780 134904 531832 134910
rect 531778 134872 531780 134881
rect 535000 134904 535052 134910
rect 531832 134872 531834 134881
rect 535000 134846 535052 134852
rect 531778 134807 531834 134816
rect 531780 133544 531832 133550
rect 531780 133486 531832 133492
rect 531792 133385 531820 133486
rect 531778 133376 531834 133385
rect 531778 133311 531834 133320
rect 536024 132054 536052 141879
rect 536208 133550 536236 143375
rect 536746 140448 536802 140457
rect 536746 140383 536802 140392
rect 536654 138952 536710 138961
rect 536654 138887 536710 138896
rect 536562 137456 536618 137465
rect 536562 137391 536618 137400
rect 536470 135824 536526 135833
rect 536470 135759 536526 135768
rect 536378 134328 536434 134337
rect 536378 134263 536434 134272
rect 536196 133544 536248 133550
rect 536196 133486 536248 133492
rect 536102 132832 536158 132841
rect 536102 132767 536158 132776
rect 531412 132048 531464 132054
rect 531410 132016 531412 132025
rect 536012 132048 536064 132054
rect 531464 132016 531466 132025
rect 536012 131990 536064 131996
rect 531410 131951 531466 131960
rect 532608 130688 532660 130694
rect 532606 130656 532608 130665
rect 532660 130656 532662 130665
rect 532606 130591 532662 130600
rect 531596 129464 531648 129470
rect 531596 129406 531648 129412
rect 531608 129305 531636 129406
rect 531594 129296 531650 129305
rect 531594 129231 531650 129240
rect 531964 128104 532016 128110
rect 531964 128046 532016 128052
rect 531976 127945 532004 128046
rect 531962 127936 532018 127945
rect 531962 127871 532018 127880
rect 531872 126608 531924 126614
rect 531870 126576 531872 126585
rect 531924 126576 531926 126585
rect 531870 126511 531926 126520
rect 532608 125248 532660 125254
rect 532606 125216 532608 125225
rect 532660 125216 532662 125225
rect 532606 125151 532662 125160
rect 535458 125216 535514 125225
rect 535458 125151 535514 125160
rect 531780 123888 531832 123894
rect 531778 123856 531780 123865
rect 531832 123856 531834 123865
rect 531778 123791 531834 123800
rect 532608 122528 532660 122534
rect 532606 122496 532608 122505
rect 532660 122496 532662 122505
rect 532606 122431 532662 122440
rect 532148 121168 532200 121174
rect 532146 121136 532148 121145
rect 532200 121136 532202 121145
rect 532146 121071 532202 121080
rect 532516 119944 532568 119950
rect 532516 119886 532568 119892
rect 532528 119785 532556 119886
rect 532514 119776 532570 119785
rect 532514 119711 532570 119720
rect 532608 118448 532660 118454
rect 532606 118416 532608 118425
rect 532660 118416 532662 118425
rect 532606 118351 532662 118360
rect 535472 117094 535500 125151
rect 536116 123894 536144 132767
rect 536286 131336 536342 131345
rect 536286 131271 536342 131280
rect 536194 129840 536250 129849
rect 536194 129775 536250 129784
rect 536104 123888 536156 123894
rect 536104 123830 536156 123836
rect 535642 122224 535698 122233
rect 535642 122159 535698 122168
rect 532332 117088 532384 117094
rect 532330 117056 532332 117065
rect 535460 117088 535512 117094
rect 532384 117056 532386 117065
rect 535460 117030 535512 117036
rect 532330 116991 532386 117000
rect 532608 115728 532660 115734
rect 532606 115696 532608 115705
rect 532660 115696 532662 115705
rect 532606 115631 532662 115640
rect 535550 114608 535606 114617
rect 535550 114543 535606 114552
rect 127714 114472 127770 114481
rect 127714 114407 127770 114416
rect 531688 114368 531740 114374
rect 531688 114310 531740 114316
rect 531700 114209 531728 114310
rect 531686 114200 531742 114209
rect 531686 114135 531742 114144
rect 535458 113112 535514 113121
rect 535458 113047 535514 113056
rect 531780 112940 531832 112946
rect 531780 112882 531832 112888
rect 531792 112849 531820 112882
rect 531778 112840 531834 112849
rect 531778 112775 531834 112784
rect 535472 111858 535500 113047
rect 532516 111852 532568 111858
rect 532516 111794 532568 111800
rect 535460 111852 535512 111858
rect 535460 111794 535512 111800
rect 531964 110152 532016 110158
rect 531962 110120 531964 110129
rect 532016 110120 532018 110129
rect 531962 110055 532018 110064
rect 532424 109064 532476 109070
rect 532424 109006 532476 109012
rect 531780 108928 531832 108934
rect 531780 108870 531832 108876
rect 531792 108769 531820 108870
rect 531778 108760 531834 108769
rect 531778 108695 531834 108704
rect 532240 107704 532292 107710
rect 532240 107646 532292 107652
rect 531780 107432 531832 107438
rect 531778 107400 531780 107409
rect 531832 107400 531834 107409
rect 531778 107335 531834 107344
rect 532148 106344 532200 106350
rect 532148 106286 532200 106292
rect 532056 102196 532108 102202
rect 532056 102138 532108 102144
rect 532068 96393 532096 102138
rect 532160 100609 532188 106286
rect 532252 101969 532280 107646
rect 532436 103329 532464 109006
rect 532528 106049 532556 111794
rect 535458 111616 535514 111625
rect 535458 111551 535514 111560
rect 532608 111512 532660 111518
rect 532606 111480 532608 111489
rect 532660 111480 532662 111489
rect 532606 111415 532662 111424
rect 535472 110498 535500 111551
rect 532608 110492 532660 110498
rect 532608 110434 532660 110440
rect 535460 110492 535512 110498
rect 535460 110434 535512 110440
rect 532514 106040 532570 106049
rect 532514 105975 532570 105984
rect 532516 104916 532568 104922
rect 532516 104858 532568 104864
rect 532422 103320 532478 103329
rect 532422 103255 532478 103264
rect 532238 101960 532294 101969
rect 532238 101895 532294 101904
rect 532528 100994 532556 104858
rect 532620 104689 532648 110434
rect 535458 110120 535514 110129
rect 535458 110055 535514 110064
rect 535472 109070 535500 110055
rect 535460 109064 535512 109070
rect 535460 109006 535512 109012
rect 535458 108488 535514 108497
rect 535458 108423 535514 108432
rect 535472 107710 535500 108423
rect 535460 107704 535512 107710
rect 535460 107646 535512 107652
rect 535564 107438 535592 114543
rect 535656 114374 535684 122159
rect 536208 121174 536236 129775
rect 536300 122534 536328 131271
rect 536392 125254 536420 134263
rect 536484 126614 536512 135759
rect 536576 128110 536604 137391
rect 536668 129470 536696 138887
rect 536760 130694 536788 140383
rect 536748 130688 536800 130694
rect 536748 130630 536800 130636
rect 536656 129464 536708 129470
rect 536656 129406 536708 129412
rect 536654 128344 536710 128353
rect 536654 128279 536710 128288
rect 536564 128104 536616 128110
rect 536564 128046 536616 128052
rect 536472 126608 536524 126614
rect 536472 126550 536524 126556
rect 536380 125248 536432 125254
rect 536380 125190 536432 125196
rect 536378 123720 536434 123729
rect 536378 123655 536434 123664
rect 536288 122528 536340 122534
rect 536288 122470 536340 122476
rect 536196 121168 536248 121174
rect 536196 121110 536248 121116
rect 536286 120728 536342 120737
rect 536286 120663 536342 120672
rect 536194 117600 536250 117609
rect 536194 117535 536250 117544
rect 535644 114368 535696 114374
rect 535644 114310 535696 114316
rect 536208 110158 536236 117535
rect 536300 112946 536328 120663
rect 536392 115734 536420 123655
rect 536668 119950 536696 128279
rect 536746 126712 536802 126721
rect 536746 126647 536802 126656
rect 536656 119944 536708 119950
rect 536656 119886 536708 119892
rect 536470 119232 536526 119241
rect 536470 119167 536526 119176
rect 536380 115728 536432 115734
rect 536380 115670 536432 115676
rect 536288 112940 536340 112946
rect 536288 112882 536340 112888
rect 536484 111518 536512 119167
rect 536760 118454 536788 126647
rect 536748 118448 536800 118454
rect 536748 118390 536800 118396
rect 536654 116104 536710 116113
rect 536654 116039 536710 116048
rect 536472 111512 536524 111518
rect 536472 111454 536524 111460
rect 536196 110152 536248 110158
rect 536196 110094 536248 110100
rect 536668 108934 536696 116039
rect 536656 108928 536708 108934
rect 536656 108870 536708 108876
rect 535552 107432 535604 107438
rect 535552 107374 535604 107380
rect 535458 106992 535514 107001
rect 535458 106927 535514 106936
rect 535472 106350 535500 106927
rect 535460 106344 535512 106350
rect 535460 106286 535512 106292
rect 535458 105496 535514 105505
rect 535458 105431 535514 105440
rect 535472 104922 535500 105431
rect 535460 104916 535512 104922
rect 535460 104858 535512 104864
rect 532606 104680 532662 104689
rect 532606 104615 532662 104624
rect 535458 104000 535514 104009
rect 535458 103935 535514 103944
rect 535472 103766 535500 103935
rect 532608 103760 532660 103766
rect 532608 103702 532660 103708
rect 535460 103760 535512 103766
rect 535460 103702 535512 103708
rect 532252 100966 532556 100994
rect 532146 100600 532202 100609
rect 532146 100535 532202 100544
rect 532252 99249 532280 100966
rect 532620 100858 532648 103702
rect 535458 102504 535514 102513
rect 535458 102439 535514 102448
rect 535472 102202 535500 102439
rect 535460 102196 535512 102202
rect 535460 102138 535512 102144
rect 535458 101008 535514 101017
rect 535458 100943 535514 100952
rect 532436 100830 532648 100858
rect 532238 99240 532294 99249
rect 532238 99175 532294 99184
rect 532240 98048 532292 98054
rect 532240 97990 532292 97996
rect 532148 96688 532200 96694
rect 532148 96630 532200 96636
rect 532054 96384 532110 96393
rect 532054 96319 532110 96328
rect 532056 95260 532108 95266
rect 532056 95202 532108 95208
rect 127622 91352 127678 91361
rect 127622 91287 127678 91296
rect 531964 91112 532016 91118
rect 531964 91054 532016 91060
rect 126980 89684 127032 89690
rect 126980 89626 127032 89632
rect 126992 89457 127020 89626
rect 126978 89448 127034 89457
rect 126978 89383 127034 89392
rect 126980 88324 127032 88330
rect 126980 88266 127032 88272
rect 126992 87553 127020 88266
rect 126978 87544 127034 87553
rect 126978 87479 127034 87488
rect 126980 86964 127032 86970
rect 126980 86906 127032 86912
rect 126992 85649 127020 86906
rect 531976 86873 532004 91054
rect 532068 90953 532096 95202
rect 532160 92313 532188 96630
rect 532252 93673 532280 97990
rect 532436 97889 532464 100830
rect 535472 100774 535500 100943
rect 532608 100768 532660 100774
rect 532608 100710 532660 100716
rect 535460 100768 535512 100774
rect 535460 100710 535512 100716
rect 532422 97880 532478 97889
rect 532422 97815 532478 97824
rect 532620 95033 532648 100710
rect 535458 99376 535514 99385
rect 535458 99311 535514 99320
rect 535472 98054 535500 99311
rect 535460 98048 535512 98054
rect 535460 97990 535512 97996
rect 535458 97880 535514 97889
rect 535458 97815 535514 97824
rect 535472 96694 535500 97815
rect 535460 96688 535512 96694
rect 535460 96630 535512 96636
rect 535458 96384 535514 96393
rect 535458 96319 535514 96328
rect 535472 95266 535500 96319
rect 535460 95260 535512 95266
rect 535460 95202 535512 95208
rect 532606 95024 532662 95033
rect 532606 94959 532662 94968
rect 535458 94888 535514 94897
rect 535458 94823 535514 94832
rect 535472 94246 535500 94823
rect 532516 94240 532568 94246
rect 532516 94182 532568 94188
rect 535460 94240 535512 94246
rect 535460 94182 535512 94188
rect 532238 93664 532294 93673
rect 532238 93599 532294 93608
rect 532424 92540 532476 92546
rect 532424 92482 532476 92488
rect 532146 92304 532202 92313
rect 532146 92239 532202 92248
rect 532054 90944 532110 90953
rect 532054 90879 532110 90888
rect 532056 88392 532108 88398
rect 532056 88334 532108 88340
rect 531962 86864 532018 86873
rect 531962 86799 532018 86808
rect 126978 85640 127034 85649
rect 126978 85575 127034 85584
rect 126980 84176 127032 84182
rect 532068 84153 532096 88334
rect 532436 88233 532464 92482
rect 532528 89593 532556 94182
rect 535458 93392 535514 93401
rect 535458 93327 535514 93336
rect 535472 92546 535500 93327
rect 535460 92540 535512 92546
rect 535460 92482 535512 92488
rect 535458 91896 535514 91905
rect 535458 91831 535514 91840
rect 535472 91118 535500 91831
rect 535460 91112 535512 91118
rect 535460 91054 535512 91060
rect 535458 90264 535514 90273
rect 535458 90199 535514 90208
rect 535472 89758 535500 90199
rect 532608 89752 532660 89758
rect 532608 89694 532660 89700
rect 535460 89752 535512 89758
rect 535460 89694 535512 89700
rect 532514 89584 532570 89593
rect 532514 89519 532570 89528
rect 532422 88224 532478 88233
rect 532422 88159 532478 88168
rect 532332 87032 532384 87038
rect 532332 86974 532384 86980
rect 126980 84118 127032 84124
rect 532054 84144 532110 84153
rect 126992 83745 127020 84118
rect 532054 84079 532110 84088
rect 126978 83736 127034 83745
rect 126978 83671 127034 83680
rect 122104 82816 122156 82822
rect 122104 82758 122156 82764
rect 126980 82816 127032 82822
rect 532344 82793 532372 86974
rect 532516 85604 532568 85610
rect 532516 85546 532568 85552
rect 126980 82758 127032 82764
rect 532330 82784 532386 82793
rect 126992 81841 127020 82758
rect 532330 82719 532386 82728
rect 126978 81832 127034 81841
rect 126978 81767 127034 81776
rect 532528 81433 532556 85546
rect 532620 85513 532648 89694
rect 535458 88768 535514 88777
rect 535458 88703 535514 88712
rect 535472 88398 535500 88703
rect 535460 88392 535512 88398
rect 535460 88334 535512 88340
rect 535458 87272 535514 87281
rect 535458 87207 535514 87216
rect 535472 87038 535500 87207
rect 535460 87032 535512 87038
rect 535460 86974 535512 86980
rect 535458 85776 535514 85785
rect 535458 85711 535514 85720
rect 535472 85610 535500 85711
rect 535460 85604 535512 85610
rect 535460 85546 535512 85552
rect 532606 85504 532662 85513
rect 532606 85439 532662 85448
rect 535458 84280 535514 84289
rect 532608 84244 532660 84250
rect 535458 84215 535460 84224
rect 532608 84186 532660 84192
rect 535512 84215 535514 84224
rect 535460 84186 535512 84192
rect 532514 81424 532570 81433
rect 532514 81359 532570 81368
rect 532620 80073 532648 84186
rect 535642 82784 535698 82793
rect 535642 82719 535698 82728
rect 535550 81152 535606 81161
rect 535550 81087 535606 81096
rect 532606 80064 532662 80073
rect 117964 80028 118016 80034
rect 117964 79970 118016 79976
rect 126980 80028 127032 80034
rect 532606 79999 532662 80008
rect 126980 79970 127032 79976
rect 126992 79937 127020 79970
rect 126978 79928 127034 79937
rect 126978 79863 127034 79872
rect 535458 79656 535514 79665
rect 535458 79591 535514 79600
rect 532148 78736 532200 78742
rect 532146 78704 532148 78713
rect 532200 78704 532202 78713
rect 532146 78639 532202 78648
rect 116124 77988 116176 77994
rect 116124 77930 116176 77936
rect 126980 77988 127032 77994
rect 126980 77930 127032 77936
rect 116136 77897 116164 77930
rect 126992 77897 127020 77930
rect 116122 77888 116178 77897
rect 116122 77823 116178 77832
rect 126978 77888 127034 77897
rect 126978 77823 127034 77832
rect 532608 77240 532660 77246
rect 532606 77208 532608 77217
rect 532660 77208 532662 77217
rect 532606 77143 532662 77152
rect 126978 75984 127034 75993
rect 116584 75948 116636 75954
rect 126978 75919 126980 75928
rect 116584 75890 116636 75896
rect 127032 75919 127034 75928
rect 126980 75890 127032 75896
rect 116596 66473 116624 75890
rect 535472 75886 535500 79591
rect 535564 77246 535592 81087
rect 535656 78742 535684 82719
rect 535644 78736 535696 78742
rect 535644 78678 535696 78684
rect 536286 78160 536342 78169
rect 536286 78095 536342 78104
rect 535552 77240 535604 77246
rect 535552 77182 535604 77188
rect 535550 76664 535606 76673
rect 535550 76599 535606 76608
rect 532608 75880 532660 75886
rect 532606 75848 532608 75857
rect 535460 75880 535512 75886
rect 532660 75848 532662 75857
rect 535460 75822 535512 75828
rect 532606 75783 532662 75792
rect 532608 74520 532660 74526
rect 532606 74488 532608 74497
rect 532660 74488 532662 74497
rect 532606 74423 532662 74432
rect 126978 74080 127034 74089
rect 126978 74015 127034 74024
rect 126992 73234 127020 74015
rect 116768 73228 116820 73234
rect 116768 73170 116820 73176
rect 126980 73228 127032 73234
rect 126980 73170 127032 73176
rect 116676 71800 116728 71806
rect 116676 71742 116728 71748
rect 116582 66464 116638 66473
rect 116582 66399 116638 66408
rect 115204 62144 115256 62150
rect 115204 62086 115256 62092
rect 9016 4690 9352 4706
rect 49036 4690 49372 4706
rect 55660 4690 55996 4706
rect 62376 4690 62712 4706
rect 65688 4690 66024 4706
rect 75716 4690 75868 4706
rect 79028 4690 79364 4706
rect 82340 4690 82676 4706
rect 95680 4690 96016 4706
rect 9016 4684 9364 4690
rect 9016 4678 9312 4684
rect 49036 4684 49384 4690
rect 49036 4678 49332 4684
rect 9312 4626 9364 4632
rect 55660 4684 56008 4690
rect 55660 4678 55956 4684
rect 49332 4626 49384 4632
rect 62376 4684 62724 4690
rect 62376 4678 62672 4684
rect 55956 4626 56008 4632
rect 65688 4684 66036 4690
rect 65688 4678 65984 4684
rect 62672 4626 62724 4632
rect 75716 4684 75880 4690
rect 75716 4678 75828 4684
rect 65984 4626 66036 4632
rect 79028 4684 79376 4690
rect 79028 4678 79324 4684
rect 75828 4626 75880 4632
rect 82340 4684 82688 4690
rect 82340 4678 82636 4684
rect 79324 4626 79376 4632
rect 95680 4684 96028 4690
rect 95680 4678 95976 4684
rect 82636 4626 82688 4632
rect 95976 4626 96028 4632
rect 5704 4134 6040 4162
rect 6012 3602 6040 4134
rect 12314 3890 12342 4148
rect 15640 4134 15976 4162
rect 18952 4134 19288 4162
rect 22356 4134 22692 4162
rect 25668 4134 26004 4162
rect 12314 3862 12388 3890
rect 6000 3596 6052 3602
rect 6000 3538 6052 3544
rect 12360 2786 12388 3862
rect 15948 2854 15976 4134
rect 15936 2848 15988 2854
rect 15936 2790 15988 2796
rect 12348 2780 12400 2786
rect 12348 2722 12400 2728
rect 19260 2174 19288 4134
rect 19248 2168 19300 2174
rect 19248 2110 19300 2116
rect 22664 2038 22692 4134
rect 25976 2106 26004 4134
rect 28966 3890 28994 4148
rect 32292 4134 32628 4162
rect 35696 4134 35848 4162
rect 39008 4134 39344 4162
rect 42320 4134 42656 4162
rect 45632 4134 45968 4162
rect 28920 3862 28994 3890
rect 28920 2582 28948 3862
rect 28908 2576 28960 2582
rect 28908 2518 28960 2524
rect 32600 2514 32628 4134
rect 33692 3392 33744 3398
rect 33692 3334 33744 3340
rect 32588 2508 32640 2514
rect 32588 2450 32640 2456
rect 25964 2100 26016 2106
rect 25964 2042 26016 2048
rect 22652 2032 22704 2038
rect 22652 1974 22704 1980
rect 33704 800 33732 3334
rect 35820 2446 35848 4134
rect 39316 2990 39344 4134
rect 42628 3058 42656 4134
rect 45940 3126 45968 4134
rect 52334 3890 52362 4148
rect 58972 4134 59308 4162
rect 52334 3862 52408 3890
rect 52380 3194 52408 3862
rect 52368 3188 52420 3194
rect 52368 3130 52420 3136
rect 45928 3120 45980 3126
rect 45928 3062 45980 3068
rect 42616 3052 42668 3058
rect 42616 2994 42668 3000
rect 39304 2984 39356 2990
rect 39304 2926 39356 2932
rect 35808 2440 35860 2446
rect 35808 2382 35860 2388
rect 59280 1358 59308 4134
rect 68986 3890 69014 4148
rect 72312 4134 72648 4162
rect 85652 4134 85988 4162
rect 89056 4134 89392 4162
rect 68940 3862 69014 3890
rect 68940 3262 68968 3862
rect 68928 3256 68980 3262
rect 68928 3198 68980 3204
rect 72620 2310 72648 4134
rect 72608 2304 72660 2310
rect 72608 2246 72660 2252
rect 85960 2242 85988 4134
rect 89364 3330 89392 4134
rect 92354 3890 92382 4148
rect 98992 4134 99328 4162
rect 102396 4134 102732 4162
rect 105708 4134 106044 4162
rect 92354 3862 92428 3890
rect 91100 3460 91152 3466
rect 91100 3402 91152 3408
rect 89352 3324 89404 3330
rect 89352 3266 89404 3272
rect 91112 2786 91140 3402
rect 91100 2780 91152 2786
rect 91100 2722 91152 2728
rect 92400 2378 92428 3862
rect 99300 2786 99328 4134
rect 101128 2916 101180 2922
rect 101128 2858 101180 2864
rect 99288 2780 99340 2786
rect 99288 2722 99340 2728
rect 92388 2372 92440 2378
rect 92388 2314 92440 2320
rect 85948 2236 86000 2242
rect 85948 2178 86000 2184
rect 59268 1352 59320 1358
rect 59268 1294 59320 1300
rect 101140 800 101168 2858
rect 102704 2718 102732 4134
rect 105636 3528 105688 3534
rect 105636 3470 105688 3476
rect 105648 2786 105676 3470
rect 105636 2780 105688 2786
rect 105636 2722 105688 2728
rect 102692 2712 102744 2718
rect 102692 2654 102744 2660
rect 106016 1970 106044 4134
rect 109006 3890 109034 4148
rect 112332 4134 112668 4162
rect 108960 3862 109034 3890
rect 108960 2718 108988 3862
rect 108948 2712 109000 2718
rect 108948 2654 109000 2660
rect 112640 2650 112668 4134
rect 115216 2718 115244 62086
rect 115296 57248 115348 57254
rect 115296 57190 115348 57196
rect 115204 2712 115256 2718
rect 115204 2654 115256 2660
rect 112628 2644 112680 2650
rect 112628 2586 112680 2592
rect 115308 1970 115336 57190
rect 116584 53848 116636 53854
rect 116584 53790 116636 53796
rect 115940 21140 115992 21146
rect 115940 21082 115992 21088
rect 115952 20913 115980 21082
rect 115938 20904 115994 20913
rect 115938 20839 115994 20848
rect 115388 12504 115440 12510
rect 115388 12446 115440 12452
rect 115400 2174 115428 12446
rect 116596 5370 116624 53790
rect 116688 43761 116716 71742
rect 116780 55049 116808 73170
rect 535564 73166 535592 76599
rect 535642 75168 535698 75177
rect 535642 75103 535698 75112
rect 532424 73160 532476 73166
rect 532422 73128 532424 73137
rect 535552 73160 535604 73166
rect 532476 73128 532478 73137
rect 535552 73102 535604 73108
rect 532422 73063 532478 73072
rect 126978 72176 127034 72185
rect 126978 72111 127034 72120
rect 126992 71806 127020 72111
rect 535550 72040 535606 72049
rect 535550 71975 535606 71984
rect 126980 71800 127032 71806
rect 126980 71742 127032 71748
rect 532422 71768 532478 71777
rect 532422 71703 532424 71712
rect 532476 71703 532478 71712
rect 532424 71674 532476 71680
rect 531780 70576 531832 70582
rect 531780 70518 531832 70524
rect 535458 70544 535514 70553
rect 531792 70417 531820 70518
rect 535458 70479 535514 70488
rect 531778 70408 531834 70417
rect 531778 70343 531834 70352
rect 126978 70272 127034 70281
rect 126978 70207 127034 70216
rect 126992 69086 127020 70207
rect 531964 69828 532016 69834
rect 531964 69770 532016 69776
rect 120816 69080 120868 69086
rect 120816 69022 120868 69028
rect 126980 69080 127032 69086
rect 531976 69057 532004 69770
rect 126980 69022 127032 69028
rect 531962 69048 532018 69057
rect 118056 67652 118108 67658
rect 118056 67594 118108 67600
rect 116766 55040 116822 55049
rect 116766 54975 116822 54984
rect 117964 53100 118016 53106
rect 117964 53042 118016 53048
rect 116674 43752 116730 43761
rect 116674 43687 116730 43696
rect 116676 37324 116728 37330
rect 116676 37266 116728 37272
rect 116584 5364 116636 5370
rect 116584 5306 116636 5312
rect 116688 5098 116716 37266
rect 116860 33380 116912 33386
rect 116860 33322 116912 33328
rect 116872 32337 116900 33322
rect 116858 32328 116914 32337
rect 116858 32263 116914 32272
rect 116768 24880 116820 24886
rect 116768 24822 116820 24828
rect 116676 5092 116728 5098
rect 116676 5034 116728 5040
rect 116780 3058 116808 24822
rect 117226 9616 117282 9625
rect 117226 9551 117282 9560
rect 117240 9110 117268 9551
rect 117228 9104 117280 9110
rect 117228 9046 117280 9052
rect 117228 4208 117280 4214
rect 117228 4150 117280 4156
rect 117240 3602 117268 4150
rect 117228 3596 117280 3602
rect 117228 3538 117280 3544
rect 116768 3052 116820 3058
rect 116768 2994 116820 3000
rect 117976 2786 118004 53042
rect 118068 21146 118096 67594
rect 119344 63572 119396 63578
rect 119344 63514 119396 63520
rect 118148 38684 118200 38690
rect 118148 38626 118200 38632
rect 118056 21140 118108 21146
rect 118056 21082 118108 21088
rect 118056 13864 118108 13870
rect 118056 13806 118108 13812
rect 117964 2780 118016 2786
rect 117964 2722 118016 2728
rect 115388 2168 115440 2174
rect 115388 2110 115440 2116
rect 118068 2038 118096 13806
rect 118160 3262 118188 38626
rect 118148 3256 118200 3262
rect 118148 3198 118200 3204
rect 119356 2650 119384 63514
rect 120724 51128 120776 51134
rect 120724 51070 120776 51076
rect 119436 42832 119488 42838
rect 119436 42774 119488 42780
rect 119448 5166 119476 42774
rect 119528 27668 119580 27674
rect 119528 27610 119580 27616
rect 119436 5160 119488 5166
rect 119436 5102 119488 5108
rect 119540 3126 119568 27610
rect 120736 3330 120764 51070
rect 120828 33386 120856 69022
rect 531962 68983 532018 68992
rect 126978 68368 127034 68377
rect 126978 68303 127034 68312
rect 126992 67658 127020 68303
rect 535472 68202 535500 70479
rect 535564 69834 535592 71975
rect 535656 71738 535684 75103
rect 536300 74526 536328 78095
rect 536288 74520 536340 74526
rect 536288 74462 536340 74468
rect 535734 73672 535790 73681
rect 535734 73607 535790 73616
rect 535644 71732 535696 71738
rect 535644 71674 535696 71680
rect 535748 70582 535776 73607
rect 535736 70576 535788 70582
rect 535736 70518 535788 70524
rect 535552 69828 535604 69834
rect 535552 69770 535604 69776
rect 535550 69048 535606 69057
rect 535550 68983 535606 68992
rect 531964 68196 532016 68202
rect 531964 68138 532016 68144
rect 535460 68196 535512 68202
rect 535460 68138 535512 68144
rect 531976 67697 532004 68138
rect 531962 67688 532018 67697
rect 126980 67652 127032 67658
rect 531962 67623 532018 67632
rect 126980 67594 127032 67600
rect 535564 67590 535592 68983
rect 531964 67584 532016 67590
rect 535552 67584 535604 67590
rect 531964 67526 532016 67532
rect 535458 67552 535514 67561
rect 127438 66464 127494 66473
rect 127438 66399 127494 66408
rect 127452 66298 127480 66399
rect 531976 66337 532004 67526
rect 535552 67526 535604 67532
rect 535458 67487 535514 67496
rect 531962 66328 532018 66337
rect 124864 66292 124916 66298
rect 124864 66234 124916 66240
rect 127440 66292 127492 66298
rect 535472 66298 535500 67487
rect 531962 66263 532018 66272
rect 535460 66292 535512 66298
rect 127440 66234 127492 66240
rect 535460 66234 535512 66240
rect 123484 46980 123536 46986
rect 123484 46922 123536 46928
rect 122104 44192 122156 44198
rect 122104 44134 122156 44140
rect 120816 33380 120868 33386
rect 120816 33322 120868 33328
rect 120816 29028 120868 29034
rect 120816 28970 120868 28976
rect 120828 4894 120856 28970
rect 120908 18012 120960 18018
rect 120908 17954 120960 17960
rect 120816 4888 120868 4894
rect 120816 4830 120868 4836
rect 120724 3324 120776 3330
rect 120724 3266 120776 3272
rect 119528 3120 119580 3126
rect 119528 3062 119580 3068
rect 119344 2644 119396 2650
rect 119344 2586 119396 2592
rect 120920 2582 120948 17954
rect 122116 5234 122144 44134
rect 122196 31816 122248 31822
rect 122196 31758 122248 31764
rect 122104 5228 122156 5234
rect 122104 5170 122156 5176
rect 122208 3194 122236 31758
rect 122288 19372 122340 19378
rect 122288 19314 122340 19320
rect 122196 3188 122248 3194
rect 122196 3130 122248 3136
rect 120908 2576 120960 2582
rect 120908 2518 120960 2524
rect 122300 2514 122328 19314
rect 123496 5302 123524 46922
rect 123576 33176 123628 33182
rect 123576 33118 123628 33124
rect 123484 5296 123536 5302
rect 123484 5238 123536 5244
rect 123588 4962 123616 33118
rect 123668 22160 123720 22166
rect 123668 22102 123720 22108
rect 123576 4956 123628 4962
rect 123576 4898 123628 4904
rect 122288 2508 122340 2514
rect 122288 2450 122340 2456
rect 123680 2446 123708 22102
rect 124876 9110 124904 66234
rect 532148 66224 532200 66230
rect 532148 66166 532200 66172
rect 532160 64977 532188 66166
rect 535458 66056 535514 66065
rect 535458 65991 535514 66000
rect 532146 64968 532202 64977
rect 535472 64938 535500 65991
rect 532146 64903 532202 64912
rect 535460 64932 535512 64938
rect 535460 64874 535512 64880
rect 531320 64864 531372 64870
rect 531320 64806 531372 64812
rect 126978 64560 127034 64569
rect 126978 64495 127034 64504
rect 126992 63578 127020 64495
rect 531332 63617 531360 64806
rect 535458 64560 535514 64569
rect 535458 64495 535514 64504
rect 531318 63608 531374 63617
rect 126980 63572 127032 63578
rect 535472 63578 535500 64495
rect 531318 63543 531374 63552
rect 535460 63572 535512 63578
rect 126980 63514 127032 63520
rect 535460 63514 535512 63520
rect 532148 63504 532200 63510
rect 532148 63446 532200 63452
rect 126978 62520 127034 62529
rect 126978 62455 127034 62464
rect 126992 62150 127020 62455
rect 532160 62257 532188 63446
rect 535458 62928 535514 62937
rect 535458 62863 535514 62872
rect 532146 62248 532202 62257
rect 532146 62183 532202 62192
rect 535472 62150 535500 62863
rect 126980 62144 127032 62150
rect 126980 62086 127032 62092
rect 535460 62144 535512 62150
rect 535460 62086 535512 62092
rect 532332 62076 532384 62082
rect 532332 62018 532384 62024
rect 532344 60897 532372 62018
rect 535458 61432 535514 61441
rect 535458 61367 535514 61376
rect 532330 60888 532386 60897
rect 532330 60823 532386 60832
rect 535472 60790 535500 61367
rect 535460 60784 535512 60790
rect 535460 60726 535512 60732
rect 532516 60716 532568 60722
rect 532516 60658 532568 60664
rect 126978 60616 127034 60625
rect 126978 60551 127034 60560
rect 126992 57254 127020 60551
rect 532528 59401 532556 60658
rect 535458 59936 535514 59945
rect 535458 59871 535514 59880
rect 535472 59430 535500 59871
rect 535460 59424 535512 59430
rect 532514 59392 532570 59401
rect 535460 59366 535512 59372
rect 532514 59327 532570 59336
rect 532608 59356 532660 59362
rect 532608 59298 532660 59304
rect 127806 58712 127862 58721
rect 127806 58647 127862 58656
rect 126980 57248 127032 57254
rect 126980 57190 127032 57196
rect 127622 56808 127678 56817
rect 127622 56743 127678 56752
rect 126978 54904 127034 54913
rect 126978 54839 127034 54848
rect 126992 53854 127020 54839
rect 126980 53848 127032 53854
rect 126980 53790 127032 53796
rect 126980 51128 127032 51134
rect 126978 51096 126980 51105
rect 127032 51096 127034 51105
rect 126978 51031 127034 51040
rect 126242 49056 126298 49065
rect 126242 48991 126298 49000
rect 124956 41472 125008 41478
rect 124956 41414 125008 41420
rect 124864 9104 124916 9110
rect 124864 9046 124916 9052
rect 124312 9036 124364 9042
rect 124312 8978 124364 8984
rect 123668 2440 123720 2446
rect 123668 2382 123720 2388
rect 124324 2106 124352 8978
rect 124864 5568 124916 5574
rect 124864 5510 124916 5516
rect 124876 4826 124904 5510
rect 124864 4820 124916 4826
rect 124864 4762 124916 4768
rect 124968 2310 124996 41414
rect 125048 10940 125100 10946
rect 125048 10882 125100 10888
rect 125060 2378 125088 10882
rect 125048 2372 125100 2378
rect 125048 2314 125100 2320
rect 124956 2304 125008 2310
rect 124956 2246 125008 2252
rect 126256 2242 126284 48991
rect 126978 47152 127034 47161
rect 126978 47087 127034 47096
rect 126992 46986 127020 47087
rect 126980 46980 127032 46986
rect 126980 46922 127032 46928
rect 126978 45248 127034 45257
rect 126978 45183 127034 45192
rect 126992 44198 127020 45183
rect 126980 44192 127032 44198
rect 126980 44134 127032 44140
rect 126978 43344 127034 43353
rect 126978 43279 127034 43288
rect 126992 42838 127020 43279
rect 126980 42832 127032 42838
rect 126980 42774 127032 42780
rect 126980 41472 127032 41478
rect 126978 41440 126980 41449
rect 127032 41440 127034 41449
rect 126978 41375 127034 41384
rect 126978 39536 127034 39545
rect 126978 39471 127034 39480
rect 126992 38690 127020 39471
rect 126980 38684 127032 38690
rect 126980 38626 127032 38632
rect 126978 37632 127034 37641
rect 126978 37567 127034 37576
rect 126992 37330 127020 37567
rect 126980 37324 127032 37330
rect 126980 37266 127032 37272
rect 126334 35728 126390 35737
rect 126334 35663 126390 35672
rect 126348 5030 126376 35663
rect 126978 33688 127034 33697
rect 126978 33623 127034 33632
rect 126992 33182 127020 33623
rect 126980 33176 127032 33182
rect 126980 33118 127032 33124
rect 126980 31816 127032 31822
rect 126978 31784 126980 31793
rect 127032 31784 127034 31793
rect 126978 31719 127034 31728
rect 126978 29880 127034 29889
rect 126978 29815 127034 29824
rect 126992 29034 127020 29815
rect 126980 29028 127032 29034
rect 126980 28970 127032 28976
rect 126978 27976 127034 27985
rect 126978 27911 127034 27920
rect 126992 27674 127020 27911
rect 126980 27668 127032 27674
rect 126980 27610 127032 27616
rect 126978 26072 127034 26081
rect 126978 26007 127034 26016
rect 126992 24886 127020 26007
rect 126980 24880 127032 24886
rect 126980 24822 127032 24828
rect 126426 24168 126482 24177
rect 126426 24103 126482 24112
rect 126336 5024 126388 5030
rect 126336 4966 126388 4972
rect 126440 2990 126468 24103
rect 126978 22264 127034 22273
rect 126978 22199 127034 22208
rect 126992 22166 127020 22199
rect 126980 22160 127032 22166
rect 126980 22102 127032 22108
rect 126978 20360 127034 20369
rect 126978 20295 127034 20304
rect 126992 19378 127020 20295
rect 126980 19372 127032 19378
rect 126980 19314 127032 19320
rect 126978 18320 127034 18329
rect 126978 18255 127034 18264
rect 126992 18018 127020 18255
rect 126980 18012 127032 18018
rect 126980 17954 127032 17960
rect 127254 16416 127310 16425
rect 127254 16351 127310 16360
rect 126978 14512 127034 14521
rect 126978 14447 127034 14456
rect 126992 13870 127020 14447
rect 126980 13864 127032 13870
rect 126980 13806 127032 13812
rect 126978 12608 127034 12617
rect 126978 12543 127034 12552
rect 126992 12510 127020 12543
rect 126980 12504 127032 12510
rect 126980 12446 127032 12452
rect 127268 9042 127296 16351
rect 127256 9036 127308 9042
rect 127256 8978 127308 8984
rect 126978 6896 127034 6905
rect 126978 6831 127034 6840
rect 126992 5574 127020 6831
rect 126980 5568 127032 5574
rect 126980 5510 127032 5516
rect 126978 4992 127034 5001
rect 126978 4927 127034 4936
rect 126992 4214 127020 4927
rect 126980 4208 127032 4214
rect 126980 4150 127032 4156
rect 127636 3534 127664 56743
rect 127820 53106 127848 58647
rect 532620 58041 532648 59298
rect 535458 58440 535514 58449
rect 535458 58375 535514 58384
rect 532606 58032 532662 58041
rect 535472 58002 535500 58375
rect 532606 57967 532662 57976
rect 535460 57996 535512 58002
rect 535460 57938 535512 57944
rect 532424 57928 532476 57934
rect 532424 57870 532476 57876
rect 532436 56681 532464 57870
rect 535458 56944 535514 56953
rect 535458 56879 535514 56888
rect 532422 56672 532478 56681
rect 535472 56642 535500 56879
rect 532422 56607 532478 56616
rect 535460 56636 535512 56642
rect 535460 56578 535512 56584
rect 532608 56568 532660 56574
rect 532608 56510 532660 56516
rect 532620 55321 532648 56510
rect 535458 55448 535514 55457
rect 535458 55383 535514 55392
rect 532606 55312 532662 55321
rect 535472 55282 535500 55383
rect 532606 55247 532662 55256
rect 535460 55276 535512 55282
rect 535460 55218 535512 55224
rect 531320 55208 531372 55214
rect 531320 55150 531372 55156
rect 531332 53961 531360 55150
rect 531318 53952 531374 53961
rect 531318 53887 531374 53896
rect 535458 53816 535514 53825
rect 535458 53751 535514 53760
rect 127808 53100 127860 53106
rect 127808 53042 127860 53048
rect 535472 53038 535500 53751
rect 532148 53032 532200 53038
rect 127714 53000 127770 53009
rect 532148 52974 532200 52980
rect 535460 53032 535512 53038
rect 535460 52974 535512 52980
rect 127714 52935 127770 52944
rect 127728 10946 127756 52935
rect 532160 52601 532188 52974
rect 532146 52592 532202 52601
rect 532146 52527 532202 52536
rect 535458 52320 535514 52329
rect 535458 52255 535514 52264
rect 535472 51338 535500 52255
rect 532608 51332 532660 51338
rect 532608 51274 532660 51280
rect 535460 51332 535512 51338
rect 535460 51274 535512 51280
rect 532620 51241 532648 51274
rect 532606 51232 532662 51241
rect 532606 51167 532662 51176
rect 535458 50824 535514 50833
rect 535458 50759 535514 50768
rect 535472 50046 535500 50759
rect 532516 50040 532568 50046
rect 532516 49982 532568 49988
rect 535460 50040 535512 50046
rect 535460 49982 535512 49988
rect 532528 49881 532556 49982
rect 532514 49872 532570 49881
rect 532514 49807 532570 49816
rect 535458 49328 535514 49337
rect 535458 49263 535514 49272
rect 535472 48686 535500 49263
rect 531964 48680 532016 48686
rect 531964 48622 532016 48628
rect 535460 48680 535512 48686
rect 535460 48622 535512 48628
rect 531976 48521 532004 48622
rect 531962 48512 532018 48521
rect 531962 48447 532018 48456
rect 535458 47832 535514 47841
rect 535458 47767 535514 47776
rect 535472 47462 535500 47767
rect 532608 47456 532660 47462
rect 532608 47398 532660 47404
rect 535460 47456 535512 47462
rect 535460 47398 535512 47404
rect 532620 47161 532648 47398
rect 532606 47152 532662 47161
rect 532606 47087 532662 47096
rect 535458 46336 535514 46345
rect 535458 46271 535514 46280
rect 535472 45830 535500 46271
rect 532608 45824 532660 45830
rect 532606 45792 532608 45801
rect 535460 45824 535512 45830
rect 532660 45792 532662 45801
rect 535460 45766 535512 45772
rect 532606 45727 532662 45736
rect 535458 44704 535514 44713
rect 535458 44639 535514 44648
rect 535472 44606 535500 44639
rect 532516 44600 532568 44606
rect 532516 44542 532568 44548
rect 535460 44600 535512 44606
rect 535460 44542 535512 44548
rect 532528 44441 532556 44542
rect 532514 44432 532570 44441
rect 532514 44367 532570 44376
rect 535458 43208 535514 43217
rect 535458 43143 535514 43152
rect 535472 43110 535500 43143
rect 532608 43104 532660 43110
rect 532606 43072 532608 43081
rect 535460 43104 535512 43110
rect 532660 43072 532662 43081
rect 535460 43046 535512 43052
rect 532606 43007 532662 43016
rect 532608 41744 532660 41750
rect 532606 41712 532608 41721
rect 535460 41744 535512 41750
rect 532660 41712 532662 41721
rect 532606 41647 532662 41656
rect 535458 41712 535460 41721
rect 535512 41712 535514 41721
rect 535458 41647 535514 41656
rect 532606 40216 532662 40225
rect 532606 40151 532608 40160
rect 532660 40151 532662 40160
rect 535458 40216 535514 40225
rect 535458 40151 535460 40160
rect 532608 40122 532660 40128
rect 535512 40151 535514 40160
rect 535460 40122 535512 40128
rect 532606 38856 532662 38865
rect 532606 38791 532608 38800
rect 532660 38791 532662 38800
rect 535460 38820 535512 38826
rect 532608 38762 532660 38768
rect 535460 38762 535512 38768
rect 535472 38729 535500 38762
rect 535458 38720 535514 38729
rect 535458 38655 535514 38664
rect 532606 37496 532662 37505
rect 532606 37431 532608 37440
rect 532660 37431 532662 37440
rect 535368 37460 535420 37466
rect 532608 37402 532660 37408
rect 535368 37402 535420 37408
rect 535380 37233 535408 37402
rect 535366 37224 535422 37233
rect 535366 37159 535422 37168
rect 532330 36136 532386 36145
rect 532330 36071 532332 36080
rect 532384 36071 532386 36080
rect 535368 36100 535420 36106
rect 532332 36042 532384 36048
rect 535368 36042 535420 36048
rect 535380 35601 535408 36042
rect 535366 35592 535422 35601
rect 535366 35527 535422 35536
rect 532606 34776 532662 34785
rect 532606 34711 532608 34720
rect 532660 34711 532662 34720
rect 535368 34740 535420 34746
rect 532608 34682 532660 34688
rect 535368 34682 535420 34688
rect 535380 34105 535408 34682
rect 535366 34096 535422 34105
rect 535366 34031 535422 34040
rect 531962 33416 532018 33425
rect 531962 33351 531964 33360
rect 532016 33351 532018 33360
rect 535368 33380 535420 33386
rect 531964 33322 532016 33328
rect 535368 33322 535420 33328
rect 535380 32609 535408 33322
rect 535366 32600 535422 32609
rect 535366 32535 535422 32544
rect 532606 32056 532662 32065
rect 532606 31991 532608 32000
rect 532660 31991 532662 32000
rect 535368 32020 535420 32026
rect 532608 31962 532660 31968
rect 535368 31962 535420 31968
rect 535380 31113 535408 31962
rect 535366 31104 535422 31113
rect 535366 31039 535422 31048
rect 532606 30696 532662 30705
rect 532606 30631 532608 30640
rect 532660 30631 532662 30640
rect 535368 30660 535420 30666
rect 532608 30602 532660 30608
rect 535368 30602 535420 30608
rect 535380 29617 535408 30602
rect 535366 29608 535422 29617
rect 535366 29543 535422 29552
rect 532606 29336 532662 29345
rect 532606 29271 532608 29280
rect 532660 29271 532662 29280
rect 535368 29300 535420 29306
rect 532608 29242 532660 29248
rect 535368 29242 535420 29248
rect 535380 28121 535408 29242
rect 535366 28112 535422 28121
rect 535366 28047 535422 28056
rect 532606 27976 532662 27985
rect 532606 27911 532662 27920
rect 532620 27674 532648 27911
rect 532608 27668 532660 27674
rect 532608 27610 532660 27616
rect 535460 27600 535512 27606
rect 535460 27542 535512 27548
rect 532330 26616 532386 26625
rect 532330 26551 532332 26560
rect 532384 26551 532386 26560
rect 535368 26580 535420 26586
rect 532332 26522 532384 26528
rect 535368 26522 535420 26528
rect 532606 25256 532662 25265
rect 532606 25191 532662 25200
rect 532620 24886 532648 25191
rect 535380 24993 535408 26522
rect 535472 26489 535500 27542
rect 535458 26480 535514 26489
rect 535458 26415 535514 26424
rect 535366 24984 535422 24993
rect 535366 24919 535422 24928
rect 532608 24880 532660 24886
rect 532608 24822 532660 24828
rect 535368 24880 535420 24886
rect 535368 24822 535420 24828
rect 532054 23896 532110 23905
rect 532054 23831 532110 23840
rect 532068 23730 532096 23831
rect 532056 23724 532108 23730
rect 532056 23666 532108 23672
rect 535276 23724 535328 23730
rect 535276 23666 535328 23672
rect 531962 22400 532018 22409
rect 531962 22335 531964 22344
rect 532016 22335 532018 22344
rect 531964 22306 532016 22312
rect 535288 22001 535316 23666
rect 535380 23497 535408 24822
rect 535366 23488 535422 23497
rect 535366 23423 535422 23432
rect 535368 22364 535420 22370
rect 535368 22306 535420 22312
rect 535274 21992 535330 22001
rect 535274 21927 535330 21936
rect 531962 21040 532018 21049
rect 531962 20975 531964 20984
rect 532016 20975 532018 20984
rect 535276 21004 535328 21010
rect 531964 20946 532016 20952
rect 535276 20946 535328 20952
rect 531962 19680 532018 19689
rect 531962 19615 531964 19624
rect 532016 19615 532018 19624
rect 535184 19644 535236 19650
rect 531964 19586 532016 19592
rect 535184 19586 535236 19592
rect 532330 18320 532386 18329
rect 532330 18255 532386 18264
rect 532344 18018 532372 18255
rect 532332 18012 532384 18018
rect 532332 17954 532384 17960
rect 535196 17377 535224 19586
rect 535288 19009 535316 20946
rect 535380 20505 535408 22306
rect 535366 20496 535422 20505
rect 535366 20431 535422 20440
rect 535274 19000 535330 19009
rect 535274 18935 535330 18944
rect 535368 18012 535420 18018
rect 535368 17954 535420 17960
rect 535182 17368 535238 17377
rect 535182 17303 535238 17312
rect 532238 16960 532294 16969
rect 532238 16895 532240 16904
rect 532292 16895 532294 16904
rect 535276 16924 535328 16930
rect 532240 16866 532292 16872
rect 535276 16866 535328 16872
rect 532606 15600 532662 15609
rect 532606 15535 532608 15544
rect 532660 15535 532662 15544
rect 532608 15506 532660 15512
rect 535288 14385 535316 16866
rect 535380 15881 535408 17954
rect 535366 15872 535422 15881
rect 535366 15807 535422 15816
rect 535368 15564 535420 15570
rect 535368 15506 535420 15512
rect 535274 14376 535330 14385
rect 535274 14311 535330 14320
rect 532146 14240 532202 14249
rect 532146 14175 532148 14184
rect 532200 14175 532202 14184
rect 535276 14204 535328 14210
rect 532148 14146 532200 14152
rect 535276 14146 535328 14152
rect 531594 12880 531650 12889
rect 531594 12815 531650 12824
rect 531608 12714 531636 12815
rect 531596 12708 531648 12714
rect 531596 12650 531648 12656
rect 531962 11520 532018 11529
rect 531962 11455 532018 11464
rect 531976 11354 532004 11455
rect 535288 11393 535316 14146
rect 535380 12889 535408 15506
rect 535366 12880 535422 12889
rect 535366 12815 535422 12824
rect 535368 12708 535420 12714
rect 535368 12650 535420 12656
rect 535274 11384 535330 11393
rect 531964 11348 532016 11354
rect 531964 11290 532016 11296
rect 535184 11348 535236 11354
rect 535274 11319 535330 11328
rect 535184 11290 535236 11296
rect 127716 10940 127768 10946
rect 127716 10882 127768 10888
rect 127714 10704 127770 10713
rect 127714 10639 127770 10648
rect 127624 3528 127676 3534
rect 127624 3470 127676 3476
rect 126428 2984 126480 2990
rect 126428 2926 126480 2932
rect 127728 2854 127756 10639
rect 531778 10160 531834 10169
rect 531778 10095 531834 10104
rect 531792 9722 531820 10095
rect 531780 9716 531832 9722
rect 531780 9658 531832 9664
rect 535000 9716 535052 9722
rect 535000 9658 535052 9664
rect 127806 8800 127862 8809
rect 127806 8735 127862 8744
rect 532238 8800 532294 8809
rect 532238 8735 532294 8744
rect 127820 3466 127848 8735
rect 532252 8362 532280 8735
rect 532240 8356 532292 8362
rect 532240 8298 532292 8304
rect 531962 7440 532018 7449
rect 531962 7375 532018 7384
rect 531976 7138 532004 7375
rect 531964 7132 532016 7138
rect 531964 7074 532016 7080
rect 535012 6769 535040 9658
rect 535196 8265 535224 11290
rect 535380 9897 535408 12650
rect 535366 9888 535422 9897
rect 535366 9823 535422 9832
rect 535276 8356 535328 8362
rect 535276 8298 535328 8304
rect 535182 8256 535238 8265
rect 535182 8191 535238 8200
rect 535184 7132 535236 7138
rect 535184 7074 535236 7080
rect 534998 6760 535054 6769
rect 534998 6695 535054 6704
rect 531594 6080 531650 6089
rect 531594 6015 531650 6024
rect 531608 5914 531636 6015
rect 531596 5908 531648 5914
rect 531596 5850 531648 5856
rect 532606 4720 532662 4729
rect 532606 4655 532662 4664
rect 532620 4554 532648 4655
rect 532608 4548 532660 4554
rect 532608 4490 532660 4496
rect 127808 3460 127860 3466
rect 127808 3402 127860 3408
rect 128360 3392 128412 3398
rect 128360 3334 128412 3340
rect 127716 2848 127768 2854
rect 127716 2790 127768 2796
rect 128372 2718 128400 3334
rect 146680 2718 146708 4148
rect 179984 2786 180012 4148
rect 179972 2780 180024 2786
rect 179972 2722 180024 2728
rect 128360 2712 128412 2718
rect 128360 2654 128412 2660
rect 146668 2712 146720 2718
rect 146668 2654 146720 2660
rect 126244 2236 126296 2242
rect 126244 2178 126296 2184
rect 213288 2174 213316 4148
rect 236184 2848 236236 2854
rect 236184 2790 236236 2796
rect 168656 2168 168708 2174
rect 168656 2110 168708 2116
rect 213276 2168 213328 2174
rect 213276 2110 213328 2116
rect 124312 2100 124364 2106
rect 124312 2042 124364 2048
rect 118056 2032 118108 2038
rect 118056 1974 118108 1980
rect 106004 1964 106056 1970
rect 106004 1906 106056 1912
rect 115296 1964 115348 1970
rect 115296 1906 115348 1912
rect 168668 800 168696 2110
rect 183468 2100 183520 2106
rect 183468 2042 183520 2048
rect 183480 1358 183508 2042
rect 183468 1352 183520 1358
rect 183468 1294 183520 1300
rect 236196 800 236224 2790
rect 246684 2786 246712 4148
rect 279988 2854 280016 4148
rect 313292 2922 313320 4148
rect 313280 2916 313332 2922
rect 313280 2858 313332 2864
rect 346688 2854 346716 4148
rect 371148 2916 371200 2922
rect 371148 2858 371200 2864
rect 279976 2848 280028 2854
rect 279976 2790 280028 2796
rect 303712 2848 303764 2854
rect 303712 2790 303764 2796
rect 346676 2848 346728 2854
rect 346676 2790 346728 2796
rect 246672 2780 246724 2786
rect 246672 2722 246724 2728
rect 303724 800 303752 2790
rect 371160 800 371188 2858
rect 379992 2106 380020 4148
rect 535196 3777 535224 7074
rect 535288 5273 535316 8298
rect 535368 5908 535420 5914
rect 535368 5850 535420 5856
rect 535274 5264 535330 5273
rect 535274 5199 535330 5208
rect 535182 3768 535238 3777
rect 535182 3703 535238 3712
rect 438676 2848 438728 2854
rect 438676 2790 438728 2796
rect 379980 2100 380032 2106
rect 379980 2042 380032 2048
rect 438688 800 438716 2790
rect 535380 2281 535408 5850
rect 535460 4548 535512 4554
rect 535460 4490 535512 4496
rect 535366 2272 535422 2281
rect 535366 2207 535422 2216
rect 506204 2100 506256 2106
rect 506204 2042 506256 2048
rect 506216 800 506244 2042
rect 33690 0 33746 800
rect 101126 0 101182 800
rect 168654 0 168710 800
rect 236182 0 236238 800
rect 303710 0 303766 800
rect 371146 0 371202 800
rect 438674 0 438730 800
rect 506202 0 506258 800
rect 535472 785 535500 4490
rect 535458 776 535514 785
rect 535458 711 535514 720
<< via2 >>
rect 8114 160656 8170 160712
rect 9034 155216 9090 155272
rect 15934 155352 15990 155408
rect 40222 156712 40278 156768
rect 36726 156576 36782 156632
rect 43718 156848 43774 156904
rect 48870 158752 48926 158808
rect 46386 157936 46442 157992
rect 26606 153312 26662 153368
rect 5998 153176 6054 153232
rect 12806 151816 12862 151872
rect 54114 157120 54170 157176
rect 55862 159296 55918 159352
rect 54942 156984 54998 157040
rect 49606 152360 49662 152416
rect 62762 159568 62818 159624
rect 65338 155624 65394 155680
rect 69662 160928 69718 160984
rect 72330 160792 72386 160848
rect 73158 159704 73214 159760
rect 68834 159432 68890 159488
rect 64510 155488 64566 155544
rect 75734 159976 75790 160032
rect 83554 161064 83610 161120
rect 86130 158072 86186 158128
rect 69662 153040 69718 153096
rect 56506 152632 56562 152688
rect 89718 157800 89774 157856
rect 97446 161200 97502 161256
rect 96526 159840 96582 159896
rect 100022 159160 100078 159216
rect 100758 158616 100814 158672
rect 107842 158208 107898 158264
rect 109590 157256 109646 157312
rect 97814 155896 97870 155952
rect 95698 155760 95754 155816
rect 93122 152496 93178 152552
rect 112994 158344 113050 158400
rect 115662 155080 115718 155136
rect 117318 161336 117374 161392
rect 9402 151272 9458 151328
rect 23110 151272 23166 151328
rect 33506 151272 33562 151328
rect 117962 153312 118018 153368
rect 116674 146104 116730 146160
rect 116582 134680 116638 134736
rect 115938 89120 115994 89176
rect 116674 123256 116730 123312
rect 116766 111968 116822 112024
rect 119342 151816 119398 151872
rect 116950 100544 117006 100600
rect 119434 150728 119490 150784
rect 120722 153176 120778 153232
rect 126886 158480 126942 158536
rect 122102 150592 122158 150648
rect 126242 150456 126298 150512
rect 128634 152904 128690 152960
rect 130842 157800 130898 157856
rect 132406 152768 132462 152824
rect 134798 156440 134854 156496
rect 135994 160656 136050 160712
rect 136638 155216 136694 155272
rect 138018 155216 138074 155272
rect 141790 155352 141846 155408
rect 154026 153040 154082 153096
rect 154670 152360 154726 152416
rect 157246 156576 157302 156632
rect 156694 152360 156750 152416
rect 161018 157936 161074 157992
rect 159822 156712 159878 156768
rect 160466 152632 160522 152688
rect 162306 156848 162362 156904
rect 164882 158616 164938 158672
rect 166170 157392 166226 157448
rect 171046 159296 171102 159352
rect 170034 157120 170090 157176
rect 170678 156984 170734 157040
rect 172058 156576 172114 156632
rect 174082 159568 174138 159624
rect 173346 153856 173402 153912
rect 175830 159976 175886 160032
rect 176290 153720 176346 153776
rect 178406 155624 178462 155680
rect 177762 155488 177818 155544
rect 180982 159432 181038 159488
rect 181626 160928 181682 160984
rect 183650 160792 183706 160848
rect 183282 153992 183338 154048
rect 184202 159704 184258 159760
rect 187606 160656 187662 160712
rect 191838 161064 191894 161120
rect 190182 154128 190238 154184
rect 194506 159296 194562 159352
rect 193770 158072 193826 158128
rect 193678 154264 193734 154320
rect 197358 159160 197414 159216
rect 197082 154400 197138 154456
rect 200210 155896 200266 155952
rect 198922 152496 198978 152552
rect 201314 159840 201370 159896
rect 200854 155760 200910 155816
rect 202142 161200 202198 161256
rect 201406 159432 201462 159488
rect 203154 155352 203210 155408
rect 203430 155216 203486 155272
rect 209870 158208 209926 158264
rect 211158 157256 211214 157312
rect 213734 158344 213790 158400
rect 216954 161336 217010 161392
rect 215666 155080 215722 155136
rect 223946 158480 224002 158536
rect 225234 152904 225290 152960
rect 227810 152768 227866 152824
rect 229742 156440 229798 156496
rect 245842 152360 245898 152416
rect 251086 155352 251142 155408
rect 257342 156576 257398 156632
rect 257986 153856 258042 153912
rect 260562 153720 260618 153776
rect 264702 157936 264758 157992
rect 265714 153992 265770 154048
rect 268934 160656 268990 160712
rect 270406 159432 270462 159488
rect 270866 154128 270922 154184
rect 271694 156576 271750 156632
rect 274086 159296 274142 159352
rect 273442 154264 273498 154320
rect 276018 154400 276074 154456
rect 280342 159296 280398 159352
rect 280526 155216 280582 155272
rect 284666 158072 284722 158128
rect 291106 155216 291162 155272
rect 292486 156712 292542 156768
rect 313922 155352 313978 155408
rect 322938 155352 322994 155408
rect 326066 157936 326122 157992
rect 329286 155216 329342 155272
rect 331218 156576 331274 156632
rect 337658 159296 337714 159352
rect 340878 158072 340934 158128
rect 346582 156712 346638 156768
rect 347226 155352 347282 155408
rect 531594 151136 531650 151192
rect 126978 150864 127034 150920
rect 126978 148996 126980 149016
rect 126980 148996 127032 149016
rect 127032 148996 127034 149016
rect 126978 148960 127034 148996
rect 126978 147056 127034 147112
rect 126978 145152 127034 145208
rect 126978 143248 127034 143304
rect 126978 139440 127034 139496
rect 126978 137400 127034 137456
rect 126978 135496 127034 135552
rect 126978 133592 127034 133648
rect 126978 131688 127034 131744
rect 126978 129784 127034 129840
rect 126978 127880 127034 127936
rect 126978 125976 127034 126032
rect 126334 124072 126390 124128
rect 126978 122032 127034 122088
rect 126978 120128 127034 120184
rect 126978 118224 127034 118280
rect 126978 116320 127034 116376
rect 126978 112512 127034 112568
rect 126978 110608 127034 110664
rect 126978 108704 127034 108760
rect 126978 106664 127034 106720
rect 126978 104796 126980 104816
rect 126980 104796 127032 104816
rect 127032 104796 127034 104816
rect 126978 104760 127034 104796
rect 126978 102856 127034 102912
rect 126978 100952 127034 101008
rect 126978 99048 127034 99104
rect 126978 97144 127034 97200
rect 126978 95240 127034 95296
rect 126242 93200 126298 93256
rect 534722 163104 534778 163160
rect 535458 158616 535514 158672
rect 535366 157120 535422 157176
rect 535274 153992 535330 154048
rect 534906 152496 534962 152552
rect 532606 149776 532662 149832
rect 534722 149504 534778 149560
rect 532330 148416 532386 148472
rect 531962 147056 532018 147112
rect 532146 145696 532202 145752
rect 531778 144336 531834 144392
rect 531686 142976 531742 143032
rect 531962 141616 532018 141672
rect 127898 141344 127954 141400
rect 531962 140256 532018 140312
rect 534814 148008 534870 148064
rect 531594 138896 531650 138952
rect 535182 151000 535238 151056
rect 535090 146512 535146 146568
rect 534998 144880 535054 144936
rect 531410 137536 531466 137592
rect 532146 136176 532202 136232
rect 536102 161608 536158 161664
rect 536194 160112 536250 160168
rect 536286 155624 536342 155680
rect 536194 143384 536250 143440
rect 536010 141888 536066 141944
rect 531778 134852 531780 134872
rect 531780 134852 531832 134872
rect 531832 134852 531834 134872
rect 531778 134816 531834 134852
rect 531778 133320 531834 133376
rect 536746 140392 536802 140448
rect 536654 138896 536710 138952
rect 536562 137400 536618 137456
rect 536470 135768 536526 135824
rect 536378 134272 536434 134328
rect 536102 132776 536158 132832
rect 531410 131996 531412 132016
rect 531412 131996 531464 132016
rect 531464 131996 531466 132016
rect 531410 131960 531466 131996
rect 532606 130636 532608 130656
rect 532608 130636 532660 130656
rect 532660 130636 532662 130656
rect 532606 130600 532662 130636
rect 531594 129240 531650 129296
rect 531962 127880 532018 127936
rect 531870 126556 531872 126576
rect 531872 126556 531924 126576
rect 531924 126556 531926 126576
rect 531870 126520 531926 126556
rect 532606 125196 532608 125216
rect 532608 125196 532660 125216
rect 532660 125196 532662 125216
rect 532606 125160 532662 125196
rect 535458 125160 535514 125216
rect 531778 123836 531780 123856
rect 531780 123836 531832 123856
rect 531832 123836 531834 123856
rect 531778 123800 531834 123836
rect 532606 122476 532608 122496
rect 532608 122476 532660 122496
rect 532660 122476 532662 122496
rect 532606 122440 532662 122476
rect 532146 121116 532148 121136
rect 532148 121116 532200 121136
rect 532200 121116 532202 121136
rect 532146 121080 532202 121116
rect 532514 119720 532570 119776
rect 532606 118396 532608 118416
rect 532608 118396 532660 118416
rect 532660 118396 532662 118416
rect 532606 118360 532662 118396
rect 536286 131280 536342 131336
rect 536194 129784 536250 129840
rect 535642 122168 535698 122224
rect 532330 117036 532332 117056
rect 532332 117036 532384 117056
rect 532384 117036 532386 117056
rect 532330 117000 532386 117036
rect 532606 115676 532608 115696
rect 532608 115676 532660 115696
rect 532660 115676 532662 115696
rect 532606 115640 532662 115676
rect 535550 114552 535606 114608
rect 127714 114416 127770 114472
rect 531686 114144 531742 114200
rect 535458 113056 535514 113112
rect 531778 112784 531834 112840
rect 531962 110100 531964 110120
rect 531964 110100 532016 110120
rect 532016 110100 532018 110120
rect 531962 110064 532018 110100
rect 531778 108704 531834 108760
rect 531778 107380 531780 107400
rect 531780 107380 531832 107400
rect 531832 107380 531834 107400
rect 531778 107344 531834 107380
rect 535458 111560 535514 111616
rect 532606 111460 532608 111480
rect 532608 111460 532660 111480
rect 532660 111460 532662 111480
rect 532606 111424 532662 111460
rect 532514 105984 532570 106040
rect 532422 103264 532478 103320
rect 532238 101904 532294 101960
rect 535458 110064 535514 110120
rect 535458 108432 535514 108488
rect 536654 128288 536710 128344
rect 536378 123664 536434 123720
rect 536286 120672 536342 120728
rect 536194 117544 536250 117600
rect 536746 126656 536802 126712
rect 536470 119176 536526 119232
rect 536654 116048 536710 116104
rect 535458 106936 535514 106992
rect 535458 105440 535514 105496
rect 532606 104624 532662 104680
rect 535458 103944 535514 104000
rect 532146 100544 532202 100600
rect 535458 102448 535514 102504
rect 535458 100952 535514 101008
rect 532238 99184 532294 99240
rect 532054 96328 532110 96384
rect 127622 91296 127678 91352
rect 126978 89392 127034 89448
rect 126978 87488 127034 87544
rect 532422 97824 532478 97880
rect 535458 99320 535514 99376
rect 535458 97824 535514 97880
rect 535458 96328 535514 96384
rect 532606 94968 532662 95024
rect 535458 94832 535514 94888
rect 532238 93608 532294 93664
rect 532146 92248 532202 92304
rect 532054 90888 532110 90944
rect 531962 86808 532018 86864
rect 126978 85584 127034 85640
rect 535458 93336 535514 93392
rect 535458 91840 535514 91896
rect 535458 90208 535514 90264
rect 532514 89528 532570 89584
rect 532422 88168 532478 88224
rect 532054 84088 532110 84144
rect 126978 83680 127034 83736
rect 532330 82728 532386 82784
rect 126978 81776 127034 81832
rect 535458 88712 535514 88768
rect 535458 87216 535514 87272
rect 535458 85720 535514 85776
rect 532606 85448 532662 85504
rect 535458 84244 535514 84280
rect 535458 84224 535460 84244
rect 535460 84224 535512 84244
rect 535512 84224 535514 84244
rect 532514 81368 532570 81424
rect 535642 82728 535698 82784
rect 535550 81096 535606 81152
rect 532606 80008 532662 80064
rect 126978 79872 127034 79928
rect 535458 79600 535514 79656
rect 532146 78684 532148 78704
rect 532148 78684 532200 78704
rect 532200 78684 532202 78704
rect 532146 78648 532202 78684
rect 116122 77832 116178 77888
rect 126978 77832 127034 77888
rect 532606 77188 532608 77208
rect 532608 77188 532660 77208
rect 532660 77188 532662 77208
rect 532606 77152 532662 77188
rect 126978 75948 127034 75984
rect 126978 75928 126980 75948
rect 126980 75928 127032 75948
rect 127032 75928 127034 75948
rect 536286 78104 536342 78160
rect 535550 76608 535606 76664
rect 532606 75828 532608 75848
rect 532608 75828 532660 75848
rect 532660 75828 532662 75848
rect 532606 75792 532662 75828
rect 532606 74468 532608 74488
rect 532608 74468 532660 74488
rect 532660 74468 532662 74488
rect 532606 74432 532662 74468
rect 126978 74024 127034 74080
rect 116582 66408 116638 66464
rect 115938 20848 115994 20904
rect 535642 75112 535698 75168
rect 532422 73108 532424 73128
rect 532424 73108 532476 73128
rect 532476 73108 532478 73128
rect 532422 73072 532478 73108
rect 126978 72120 127034 72176
rect 535550 71984 535606 72040
rect 532422 71732 532478 71768
rect 532422 71712 532424 71732
rect 532424 71712 532476 71732
rect 532476 71712 532478 71732
rect 535458 70488 535514 70544
rect 531778 70352 531834 70408
rect 126978 70216 127034 70272
rect 116766 54984 116822 55040
rect 116674 43696 116730 43752
rect 116858 32272 116914 32328
rect 117226 9560 117282 9616
rect 531962 68992 532018 69048
rect 126978 68312 127034 68368
rect 535734 73616 535790 73672
rect 535550 68992 535606 69048
rect 531962 67632 532018 67688
rect 127438 66408 127494 66464
rect 535458 67496 535514 67552
rect 531962 66272 532018 66328
rect 535458 66000 535514 66056
rect 532146 64912 532202 64968
rect 126978 64504 127034 64560
rect 535458 64504 535514 64560
rect 531318 63552 531374 63608
rect 126978 62464 127034 62520
rect 535458 62872 535514 62928
rect 532146 62192 532202 62248
rect 535458 61376 535514 61432
rect 532330 60832 532386 60888
rect 126978 60560 127034 60616
rect 535458 59880 535514 59936
rect 532514 59336 532570 59392
rect 127806 58656 127862 58712
rect 127622 56752 127678 56808
rect 126978 54848 127034 54904
rect 126978 51076 126980 51096
rect 126980 51076 127032 51096
rect 127032 51076 127034 51096
rect 126978 51040 127034 51076
rect 126242 49000 126298 49056
rect 126978 47096 127034 47152
rect 126978 45192 127034 45248
rect 126978 43288 127034 43344
rect 126978 41420 126980 41440
rect 126980 41420 127032 41440
rect 127032 41420 127034 41440
rect 126978 41384 127034 41420
rect 126978 39480 127034 39536
rect 126978 37576 127034 37632
rect 126334 35672 126390 35728
rect 126978 33632 127034 33688
rect 126978 31764 126980 31784
rect 126980 31764 127032 31784
rect 127032 31764 127034 31784
rect 126978 31728 127034 31764
rect 126978 29824 127034 29880
rect 126978 27920 127034 27976
rect 126978 26016 127034 26072
rect 126426 24112 126482 24168
rect 126978 22208 127034 22264
rect 126978 20304 127034 20360
rect 126978 18264 127034 18320
rect 127254 16360 127310 16416
rect 126978 14456 127034 14512
rect 126978 12552 127034 12608
rect 126978 6840 127034 6896
rect 126978 4936 127034 4992
rect 535458 58384 535514 58440
rect 532606 57976 532662 58032
rect 535458 56888 535514 56944
rect 532422 56616 532478 56672
rect 535458 55392 535514 55448
rect 532606 55256 532662 55312
rect 531318 53896 531374 53952
rect 535458 53760 535514 53816
rect 127714 52944 127770 53000
rect 532146 52536 532202 52592
rect 535458 52264 535514 52320
rect 532606 51176 532662 51232
rect 535458 50768 535514 50824
rect 532514 49816 532570 49872
rect 535458 49272 535514 49328
rect 531962 48456 532018 48512
rect 535458 47776 535514 47832
rect 532606 47096 532662 47152
rect 535458 46280 535514 46336
rect 532606 45772 532608 45792
rect 532608 45772 532660 45792
rect 532660 45772 532662 45792
rect 532606 45736 532662 45772
rect 535458 44648 535514 44704
rect 532514 44376 532570 44432
rect 535458 43152 535514 43208
rect 532606 43052 532608 43072
rect 532608 43052 532660 43072
rect 532660 43052 532662 43072
rect 532606 43016 532662 43052
rect 532606 41692 532608 41712
rect 532608 41692 532660 41712
rect 532660 41692 532662 41712
rect 532606 41656 532662 41692
rect 535458 41692 535460 41712
rect 535460 41692 535512 41712
rect 535512 41692 535514 41712
rect 535458 41656 535514 41692
rect 532606 40180 532662 40216
rect 532606 40160 532608 40180
rect 532608 40160 532660 40180
rect 532660 40160 532662 40180
rect 535458 40180 535514 40216
rect 535458 40160 535460 40180
rect 535460 40160 535512 40180
rect 535512 40160 535514 40180
rect 532606 38820 532662 38856
rect 532606 38800 532608 38820
rect 532608 38800 532660 38820
rect 532660 38800 532662 38820
rect 535458 38664 535514 38720
rect 532606 37460 532662 37496
rect 532606 37440 532608 37460
rect 532608 37440 532660 37460
rect 532660 37440 532662 37460
rect 535366 37168 535422 37224
rect 532330 36100 532386 36136
rect 532330 36080 532332 36100
rect 532332 36080 532384 36100
rect 532384 36080 532386 36100
rect 535366 35536 535422 35592
rect 532606 34740 532662 34776
rect 532606 34720 532608 34740
rect 532608 34720 532660 34740
rect 532660 34720 532662 34740
rect 535366 34040 535422 34096
rect 531962 33380 532018 33416
rect 531962 33360 531964 33380
rect 531964 33360 532016 33380
rect 532016 33360 532018 33380
rect 535366 32544 535422 32600
rect 532606 32020 532662 32056
rect 532606 32000 532608 32020
rect 532608 32000 532660 32020
rect 532660 32000 532662 32020
rect 535366 31048 535422 31104
rect 532606 30660 532662 30696
rect 532606 30640 532608 30660
rect 532608 30640 532660 30660
rect 532660 30640 532662 30660
rect 535366 29552 535422 29608
rect 532606 29300 532662 29336
rect 532606 29280 532608 29300
rect 532608 29280 532660 29300
rect 532660 29280 532662 29300
rect 535366 28056 535422 28112
rect 532606 27920 532662 27976
rect 532330 26580 532386 26616
rect 532330 26560 532332 26580
rect 532332 26560 532384 26580
rect 532384 26560 532386 26580
rect 532606 25200 532662 25256
rect 535458 26424 535514 26480
rect 535366 24928 535422 24984
rect 532054 23840 532110 23896
rect 531962 22364 532018 22400
rect 531962 22344 531964 22364
rect 531964 22344 532016 22364
rect 532016 22344 532018 22364
rect 535366 23432 535422 23488
rect 535274 21936 535330 21992
rect 531962 21004 532018 21040
rect 531962 20984 531964 21004
rect 531964 20984 532016 21004
rect 532016 20984 532018 21004
rect 531962 19644 532018 19680
rect 531962 19624 531964 19644
rect 531964 19624 532016 19644
rect 532016 19624 532018 19644
rect 532330 18264 532386 18320
rect 535366 20440 535422 20496
rect 535274 18944 535330 19000
rect 535182 17312 535238 17368
rect 532238 16924 532294 16960
rect 532238 16904 532240 16924
rect 532240 16904 532292 16924
rect 532292 16904 532294 16924
rect 532606 15564 532662 15600
rect 532606 15544 532608 15564
rect 532608 15544 532660 15564
rect 532660 15544 532662 15564
rect 535366 15816 535422 15872
rect 535274 14320 535330 14376
rect 532146 14204 532202 14240
rect 532146 14184 532148 14204
rect 532148 14184 532200 14204
rect 532200 14184 532202 14204
rect 531594 12824 531650 12880
rect 531962 11464 532018 11520
rect 535366 12824 535422 12880
rect 535274 11328 535330 11384
rect 127714 10648 127770 10704
rect 531778 10104 531834 10160
rect 127806 8744 127862 8800
rect 532238 8744 532294 8800
rect 531962 7384 532018 7440
rect 535366 9832 535422 9888
rect 535182 8200 535238 8256
rect 534998 6704 535054 6760
rect 531594 6024 531650 6080
rect 532606 4664 532662 4720
rect 535274 5208 535330 5264
rect 535182 3712 535238 3768
rect 535366 2216 535422 2272
rect 535458 720 535514 776
<< metal3 >>
rect 534717 163162 534783 163165
rect 539200 163162 540000 163192
rect 534717 163160 540000 163162
rect 534717 163104 534722 163160
rect 534778 163104 540000 163160
rect 534717 163102 540000 163104
rect 534717 163099 534783 163102
rect 539200 163072 540000 163102
rect 536097 161666 536163 161669
rect 539200 161666 540000 161696
rect 536097 161664 540000 161666
rect 536097 161608 536102 161664
rect 536158 161608 540000 161664
rect 536097 161606 540000 161608
rect 536097 161603 536163 161606
rect 539200 161576 540000 161606
rect 117313 161394 117379 161397
rect 216949 161394 217015 161397
rect 117313 161392 217015 161394
rect 117313 161336 117318 161392
rect 117374 161336 216954 161392
rect 217010 161336 217015 161392
rect 117313 161334 217015 161336
rect 117313 161331 117379 161334
rect 216949 161331 217015 161334
rect 97441 161258 97507 161261
rect 202137 161258 202203 161261
rect 97441 161256 202203 161258
rect 97441 161200 97446 161256
rect 97502 161200 202142 161256
rect 202198 161200 202203 161256
rect 97441 161198 202203 161200
rect 97441 161195 97507 161198
rect 202137 161195 202203 161198
rect 83549 161122 83615 161125
rect 191833 161122 191899 161125
rect 83549 161120 191899 161122
rect 83549 161064 83554 161120
rect 83610 161064 191838 161120
rect 191894 161064 191899 161120
rect 83549 161062 191899 161064
rect 83549 161059 83615 161062
rect 191833 161059 191899 161062
rect 69657 160986 69723 160989
rect 181621 160986 181687 160989
rect 69657 160984 181687 160986
rect 69657 160928 69662 160984
rect 69718 160928 181626 160984
rect 181682 160928 181687 160984
rect 69657 160926 181687 160928
rect 69657 160923 69723 160926
rect 181621 160923 181687 160926
rect 72325 160850 72391 160853
rect 183645 160850 183711 160853
rect 72325 160848 183711 160850
rect 72325 160792 72330 160848
rect 72386 160792 183650 160848
rect 183706 160792 183711 160848
rect 72325 160790 183711 160792
rect 72325 160787 72391 160790
rect 183645 160787 183711 160790
rect 8109 160714 8175 160717
rect 135989 160714 136055 160717
rect 8109 160712 136055 160714
rect 8109 160656 8114 160712
rect 8170 160656 135994 160712
rect 136050 160656 136055 160712
rect 8109 160654 136055 160656
rect 8109 160651 8175 160654
rect 135989 160651 136055 160654
rect 187601 160714 187667 160717
rect 268929 160714 268995 160717
rect 187601 160712 268995 160714
rect 187601 160656 187606 160712
rect 187662 160656 268934 160712
rect 268990 160656 268995 160712
rect 187601 160654 268995 160656
rect 187601 160651 187667 160654
rect 268929 160651 268995 160654
rect 536189 160170 536255 160173
rect 539200 160170 540000 160200
rect 536189 160168 540000 160170
rect 536189 160112 536194 160168
rect 536250 160112 540000 160168
rect 536189 160110 540000 160112
rect 536189 160107 536255 160110
rect 539200 160080 540000 160110
rect 75729 160034 75795 160037
rect 175825 160034 175891 160037
rect 75729 160032 175891 160034
rect 75729 159976 75734 160032
rect 75790 159976 175830 160032
rect 175886 159976 175891 160032
rect 75729 159974 175891 159976
rect 75729 159971 75795 159974
rect 175825 159971 175891 159974
rect 96521 159898 96587 159901
rect 201309 159898 201375 159901
rect 96521 159896 201375 159898
rect 96521 159840 96526 159896
rect 96582 159840 201314 159896
rect 201370 159840 201375 159896
rect 96521 159838 201375 159840
rect 96521 159835 96587 159838
rect 201309 159835 201375 159838
rect 73153 159762 73219 159765
rect 184197 159762 184263 159765
rect 73153 159760 184263 159762
rect 73153 159704 73158 159760
rect 73214 159704 184202 159760
rect 184258 159704 184263 159760
rect 73153 159702 184263 159704
rect 73153 159699 73219 159702
rect 184197 159699 184263 159702
rect 62757 159626 62823 159629
rect 174077 159626 174143 159629
rect 62757 159624 174143 159626
rect 62757 159568 62762 159624
rect 62818 159568 174082 159624
rect 174138 159568 174143 159624
rect 62757 159566 174143 159568
rect 62757 159563 62823 159566
rect 174077 159563 174143 159566
rect 68829 159490 68895 159493
rect 180977 159490 181043 159493
rect 68829 159488 181043 159490
rect 68829 159432 68834 159488
rect 68890 159432 180982 159488
rect 181038 159432 181043 159488
rect 68829 159430 181043 159432
rect 68829 159427 68895 159430
rect 180977 159427 181043 159430
rect 201401 159490 201467 159493
rect 270401 159490 270467 159493
rect 201401 159488 270467 159490
rect 201401 159432 201406 159488
rect 201462 159432 270406 159488
rect 270462 159432 270467 159488
rect 201401 159430 270467 159432
rect 201401 159427 201467 159430
rect 270401 159427 270467 159430
rect 55857 159354 55923 159357
rect 171041 159354 171107 159357
rect 55857 159352 171107 159354
rect 55857 159296 55862 159352
rect 55918 159296 171046 159352
rect 171102 159296 171107 159352
rect 55857 159294 171107 159296
rect 55857 159291 55923 159294
rect 171041 159291 171107 159294
rect 194501 159354 194567 159357
rect 274081 159354 274147 159357
rect 194501 159352 274147 159354
rect 194501 159296 194506 159352
rect 194562 159296 274086 159352
rect 274142 159296 274147 159352
rect 194501 159294 274147 159296
rect 194501 159291 194567 159294
rect 274081 159291 274147 159294
rect 280337 159354 280403 159357
rect 337653 159354 337719 159357
rect 280337 159352 337719 159354
rect 280337 159296 280342 159352
rect 280398 159296 337658 159352
rect 337714 159296 337719 159352
rect 280337 159294 337719 159296
rect 280337 159291 280403 159294
rect 337653 159291 337719 159294
rect 100017 159218 100083 159221
rect 197353 159218 197419 159221
rect 100017 159216 197419 159218
rect 100017 159160 100022 159216
rect 100078 159160 197358 159216
rect 197414 159160 197419 159216
rect 100017 159158 197419 159160
rect 100017 159155 100083 159158
rect 197353 159155 197419 159158
rect 48865 158810 48931 158813
rect 48998 158810 49004 158812
rect 48865 158808 49004 158810
rect 48865 158752 48870 158808
rect 48926 158752 49004 158808
rect 48865 158750 49004 158752
rect 48865 158747 48931 158750
rect 48998 158748 49004 158750
rect 49068 158748 49074 158812
rect 100753 158674 100819 158677
rect 164877 158674 164943 158677
rect 100753 158672 164943 158674
rect 100753 158616 100758 158672
rect 100814 158616 164882 158672
rect 164938 158616 164943 158672
rect 100753 158614 164943 158616
rect 100753 158611 100819 158614
rect 164877 158611 164943 158614
rect 535453 158674 535519 158677
rect 539200 158674 540000 158704
rect 535453 158672 540000 158674
rect 535453 158616 535458 158672
rect 535514 158616 540000 158672
rect 535453 158614 540000 158616
rect 535453 158611 535519 158614
rect 539200 158584 540000 158614
rect 126881 158538 126947 158541
rect 223941 158538 224007 158541
rect 126881 158536 224007 158538
rect 126881 158480 126886 158536
rect 126942 158480 223946 158536
rect 224002 158480 224007 158536
rect 126881 158478 224007 158480
rect 126881 158475 126947 158478
rect 223941 158475 224007 158478
rect 112989 158402 113055 158405
rect 213729 158402 213795 158405
rect 112989 158400 213795 158402
rect 112989 158344 112994 158400
rect 113050 158344 213734 158400
rect 213790 158344 213795 158400
rect 112989 158342 213795 158344
rect 112989 158339 113055 158342
rect 213729 158339 213795 158342
rect 107837 158266 107903 158269
rect 209865 158266 209931 158269
rect 107837 158264 209931 158266
rect 107837 158208 107842 158264
rect 107898 158208 209870 158264
rect 209926 158208 209931 158264
rect 107837 158206 209931 158208
rect 107837 158203 107903 158206
rect 209865 158203 209931 158206
rect 86125 158130 86191 158133
rect 193765 158130 193831 158133
rect 86125 158128 193831 158130
rect 86125 158072 86130 158128
rect 86186 158072 193770 158128
rect 193826 158072 193831 158128
rect 86125 158070 193831 158072
rect 86125 158067 86191 158070
rect 193765 158067 193831 158070
rect 284661 158130 284727 158133
rect 340873 158130 340939 158133
rect 284661 158128 340939 158130
rect 284661 158072 284666 158128
rect 284722 158072 340878 158128
rect 340934 158072 340939 158128
rect 284661 158070 340939 158072
rect 284661 158067 284727 158070
rect 340873 158067 340939 158070
rect 46381 157994 46447 157997
rect 161013 157994 161079 157997
rect 46381 157992 161079 157994
rect 46381 157936 46386 157992
rect 46442 157936 161018 157992
rect 161074 157936 161079 157992
rect 46381 157934 161079 157936
rect 46381 157931 46447 157934
rect 161013 157931 161079 157934
rect 264697 157994 264763 157997
rect 326061 157994 326127 157997
rect 264697 157992 326127 157994
rect 264697 157936 264702 157992
rect 264758 157936 326066 157992
rect 326122 157936 326127 157992
rect 264697 157934 326127 157936
rect 264697 157931 264763 157934
rect 326061 157931 326127 157934
rect 89713 157858 89779 157861
rect 130837 157858 130903 157861
rect 89713 157856 130903 157858
rect 89713 157800 89718 157856
rect 89774 157800 130842 157856
rect 130898 157800 130903 157856
rect 89713 157798 130903 157800
rect 89713 157795 89779 157798
rect 130837 157795 130903 157798
rect 164182 157388 164188 157452
rect 164252 157450 164258 157452
rect 166165 157450 166231 157453
rect 164252 157448 166231 157450
rect 164252 157392 166170 157448
rect 166226 157392 166231 157448
rect 164252 157390 166231 157392
rect 164252 157388 164258 157390
rect 166165 157387 166231 157390
rect 109585 157314 109651 157317
rect 211153 157314 211219 157317
rect 109585 157312 211219 157314
rect 109585 157256 109590 157312
rect 109646 157256 211158 157312
rect 211214 157256 211219 157312
rect 109585 157254 211219 157256
rect 109585 157251 109651 157254
rect 211153 157251 211219 157254
rect 54109 157178 54175 157181
rect 170029 157178 170095 157181
rect 54109 157176 170095 157178
rect 54109 157120 54114 157176
rect 54170 157120 170034 157176
rect 170090 157120 170095 157176
rect 54109 157118 170095 157120
rect 54109 157115 54175 157118
rect 170029 157115 170095 157118
rect 535361 157178 535427 157181
rect 539200 157178 540000 157208
rect 535361 157176 540000 157178
rect 535361 157120 535366 157176
rect 535422 157120 540000 157176
rect 535361 157118 540000 157120
rect 535361 157115 535427 157118
rect 539200 157088 540000 157118
rect 54937 157042 55003 157045
rect 170673 157042 170739 157045
rect 54937 157040 170739 157042
rect 54937 156984 54942 157040
rect 54998 156984 170678 157040
rect 170734 156984 170739 157040
rect 54937 156982 170739 156984
rect 54937 156979 55003 156982
rect 170673 156979 170739 156982
rect 43713 156906 43779 156909
rect 162301 156906 162367 156909
rect 43713 156904 162367 156906
rect 43713 156848 43718 156904
rect 43774 156848 162306 156904
rect 162362 156848 162367 156904
rect 43713 156846 162367 156848
rect 43713 156843 43779 156846
rect 162301 156843 162367 156846
rect 40217 156770 40283 156773
rect 159817 156770 159883 156773
rect 40217 156768 159883 156770
rect 40217 156712 40222 156768
rect 40278 156712 159822 156768
rect 159878 156712 159883 156768
rect 40217 156710 159883 156712
rect 40217 156707 40283 156710
rect 159817 156707 159883 156710
rect 292481 156770 292547 156773
rect 346577 156770 346643 156773
rect 292481 156768 346643 156770
rect 292481 156712 292486 156768
rect 292542 156712 346582 156768
rect 346638 156712 346643 156768
rect 292481 156710 346643 156712
rect 292481 156707 292547 156710
rect 346577 156707 346643 156710
rect 36721 156634 36787 156637
rect 157241 156634 157307 156637
rect 36721 156632 157307 156634
rect 36721 156576 36726 156632
rect 36782 156576 157246 156632
rect 157302 156576 157307 156632
rect 36721 156574 157307 156576
rect 36721 156571 36787 156574
rect 157241 156571 157307 156574
rect 172053 156634 172119 156637
rect 257337 156634 257403 156637
rect 172053 156632 257403 156634
rect 172053 156576 172058 156632
rect 172114 156576 257342 156632
rect 257398 156576 257403 156632
rect 172053 156574 257403 156576
rect 172053 156571 172119 156574
rect 257337 156571 257403 156574
rect 271689 156634 271755 156637
rect 331213 156634 331279 156637
rect 271689 156632 331279 156634
rect 271689 156576 271694 156632
rect 271750 156576 331218 156632
rect 331274 156576 331279 156632
rect 271689 156574 331279 156576
rect 271689 156571 271755 156574
rect 331213 156571 331279 156574
rect 134793 156498 134859 156501
rect 229737 156498 229803 156501
rect 134793 156496 229803 156498
rect 134793 156440 134798 156496
rect 134854 156440 229742 156496
rect 229798 156440 229803 156496
rect 134793 156438 229803 156440
rect 134793 156435 134859 156438
rect 229737 156435 229803 156438
rect 97809 155954 97875 155957
rect 200205 155954 200271 155957
rect 97809 155952 200271 155954
rect 97809 155896 97814 155952
rect 97870 155896 200210 155952
rect 200266 155896 200271 155952
rect 97809 155894 200271 155896
rect 97809 155891 97875 155894
rect 200205 155891 200271 155894
rect 95693 155818 95759 155821
rect 200849 155818 200915 155821
rect 95693 155816 200915 155818
rect 95693 155760 95698 155816
rect 95754 155760 200854 155816
rect 200910 155760 200915 155816
rect 95693 155758 200915 155760
rect 95693 155755 95759 155758
rect 200849 155755 200915 155758
rect 65333 155682 65399 155685
rect 178401 155682 178467 155685
rect 65333 155680 178467 155682
rect 65333 155624 65338 155680
rect 65394 155624 178406 155680
rect 178462 155624 178467 155680
rect 65333 155622 178467 155624
rect 65333 155619 65399 155622
rect 178401 155619 178467 155622
rect 536281 155682 536347 155685
rect 539200 155682 540000 155712
rect 536281 155680 540000 155682
rect 536281 155624 536286 155680
rect 536342 155624 540000 155680
rect 536281 155622 540000 155624
rect 536281 155619 536347 155622
rect 539200 155592 540000 155622
rect 64505 155546 64571 155549
rect 177757 155546 177823 155549
rect 64505 155544 177823 155546
rect 64505 155488 64510 155544
rect 64566 155488 177762 155544
rect 177818 155488 177823 155544
rect 64505 155486 177823 155488
rect 64505 155483 64571 155486
rect 177757 155483 177823 155486
rect 15929 155410 15995 155413
rect 141785 155410 141851 155413
rect 15929 155408 141851 155410
rect 15929 155352 15934 155408
rect 15990 155352 141790 155408
rect 141846 155352 141851 155408
rect 15929 155350 141851 155352
rect 15929 155347 15995 155350
rect 141785 155347 141851 155350
rect 203149 155410 203215 155413
rect 251081 155410 251147 155413
rect 313917 155410 313983 155413
rect 203149 155408 209790 155410
rect 203149 155352 203154 155408
rect 203210 155352 209790 155408
rect 203149 155350 209790 155352
rect 203149 155347 203215 155350
rect 9029 155274 9095 155277
rect 136633 155274 136699 155277
rect 9029 155272 136699 155274
rect 9029 155216 9034 155272
rect 9090 155216 136638 155272
rect 136694 155216 136699 155272
rect 9029 155214 136699 155216
rect 9029 155211 9095 155214
rect 136633 155211 136699 155214
rect 138013 155274 138079 155277
rect 203425 155274 203491 155277
rect 138013 155272 203491 155274
rect 138013 155216 138018 155272
rect 138074 155216 203430 155272
rect 203486 155216 203491 155272
rect 138013 155214 203491 155216
rect 209730 155274 209790 155350
rect 251081 155408 313983 155410
rect 251081 155352 251086 155408
rect 251142 155352 313922 155408
rect 313978 155352 313983 155408
rect 251081 155350 313983 155352
rect 251081 155347 251147 155350
rect 313917 155347 313983 155350
rect 322933 155410 322999 155413
rect 347221 155410 347287 155413
rect 322933 155408 347287 155410
rect 322933 155352 322938 155408
rect 322994 155352 347226 155408
rect 347282 155352 347287 155408
rect 322933 155350 347287 155352
rect 322933 155347 322999 155350
rect 347221 155347 347287 155350
rect 280521 155274 280587 155277
rect 209730 155272 280587 155274
rect 209730 155216 280526 155272
rect 280582 155216 280587 155272
rect 209730 155214 280587 155216
rect 138013 155211 138079 155214
rect 203425 155211 203491 155214
rect 280521 155211 280587 155214
rect 291101 155274 291167 155277
rect 329281 155274 329347 155277
rect 291101 155272 329347 155274
rect 291101 155216 291106 155272
rect 291162 155216 329286 155272
rect 329342 155216 329347 155272
rect 291101 155214 329347 155216
rect 291101 155211 291167 155214
rect 329281 155211 329347 155214
rect 115657 155138 115723 155141
rect 215661 155138 215727 155141
rect 115657 155136 215727 155138
rect 115657 155080 115662 155136
rect 115718 155080 215666 155136
rect 215722 155080 215727 155136
rect 115657 155078 215727 155080
rect 115657 155075 115723 155078
rect 215661 155075 215727 155078
rect 197077 154458 197143 154461
rect 276013 154458 276079 154461
rect 197077 154456 276079 154458
rect 197077 154400 197082 154456
rect 197138 154400 276018 154456
rect 276074 154400 276079 154456
rect 197077 154398 276079 154400
rect 197077 154395 197143 154398
rect 276013 154395 276079 154398
rect 193673 154322 193739 154325
rect 273437 154322 273503 154325
rect 193673 154320 273503 154322
rect 193673 154264 193678 154320
rect 193734 154264 273442 154320
rect 273498 154264 273503 154320
rect 193673 154262 273503 154264
rect 193673 154259 193739 154262
rect 273437 154259 273503 154262
rect 190177 154186 190243 154189
rect 270861 154186 270927 154189
rect 190177 154184 270927 154186
rect 190177 154128 190182 154184
rect 190238 154128 270866 154184
rect 270922 154128 270927 154184
rect 190177 154126 270927 154128
rect 190177 154123 190243 154126
rect 270861 154123 270927 154126
rect 183277 154050 183343 154053
rect 265709 154050 265775 154053
rect 183277 154048 265775 154050
rect 183277 153992 183282 154048
rect 183338 153992 265714 154048
rect 265770 153992 265775 154048
rect 183277 153990 265775 153992
rect 183277 153987 183343 153990
rect 265709 153987 265775 153990
rect 535269 154050 535335 154053
rect 539200 154050 540000 154080
rect 535269 154048 540000 154050
rect 535269 153992 535274 154048
rect 535330 153992 540000 154048
rect 535269 153990 540000 153992
rect 535269 153987 535335 153990
rect 539200 153960 540000 153990
rect 173341 153914 173407 153917
rect 257981 153914 258047 153917
rect 173341 153912 258047 153914
rect 173341 153856 173346 153912
rect 173402 153856 257986 153912
rect 258042 153856 258047 153912
rect 173341 153854 258047 153856
rect 173341 153851 173407 153854
rect 257981 153851 258047 153854
rect 176285 153778 176351 153781
rect 260557 153778 260623 153781
rect 176285 153776 260623 153778
rect 176285 153720 176290 153776
rect 176346 153720 260562 153776
rect 260618 153720 260623 153776
rect 176285 153718 260623 153720
rect 176285 153715 176351 153718
rect 260557 153715 260623 153718
rect 26601 153370 26667 153373
rect 117957 153370 118023 153373
rect 26601 153368 118023 153370
rect 26601 153312 26606 153368
rect 26662 153312 117962 153368
rect 118018 153312 118023 153368
rect 26601 153310 118023 153312
rect 26601 153307 26667 153310
rect 117957 153307 118023 153310
rect 5993 153234 6059 153237
rect 120717 153234 120783 153237
rect 5993 153232 120783 153234
rect 5993 153176 5998 153232
rect 6054 153176 120722 153232
rect 120778 153176 120783 153232
rect 5993 153174 120783 153176
rect 5993 153171 6059 153174
rect 120717 153171 120783 153174
rect 69657 153098 69723 153101
rect 154021 153098 154087 153101
rect 69657 153096 154087 153098
rect 69657 153040 69662 153096
rect 69718 153040 154026 153096
rect 154082 153040 154087 153096
rect 69657 153038 154087 153040
rect 69657 153035 69723 153038
rect 154021 153035 154087 153038
rect 128629 152962 128695 152965
rect 225229 152962 225295 152965
rect 128629 152960 225295 152962
rect 128629 152904 128634 152960
rect 128690 152904 225234 152960
rect 225290 152904 225295 152960
rect 128629 152902 225295 152904
rect 128629 152899 128695 152902
rect 225229 152899 225295 152902
rect 132401 152826 132467 152829
rect 227805 152826 227871 152829
rect 132401 152824 227871 152826
rect 132401 152768 132406 152824
rect 132462 152768 227810 152824
rect 227866 152768 227871 152824
rect 132401 152766 227871 152768
rect 132401 152763 132467 152766
rect 227805 152763 227871 152766
rect 56501 152690 56567 152693
rect 160461 152690 160527 152693
rect 56501 152688 160527 152690
rect 56501 152632 56506 152688
rect 56562 152632 160466 152688
rect 160522 152632 160527 152688
rect 56501 152630 160527 152632
rect 56501 152627 56567 152630
rect 160461 152627 160527 152630
rect 93117 152554 93183 152557
rect 198917 152554 198983 152557
rect 93117 152552 198983 152554
rect 93117 152496 93122 152552
rect 93178 152496 198922 152552
rect 198978 152496 198983 152552
rect 93117 152494 198983 152496
rect 93117 152491 93183 152494
rect 198917 152491 198983 152494
rect 534901 152554 534967 152557
rect 539200 152554 540000 152584
rect 534901 152552 540000 152554
rect 534901 152496 534906 152552
rect 534962 152496 540000 152552
rect 534901 152494 540000 152496
rect 534901 152491 534967 152494
rect 539200 152464 540000 152494
rect 49601 152418 49667 152421
rect 154665 152418 154731 152421
rect 49601 152416 154731 152418
rect 49601 152360 49606 152416
rect 49662 152360 154670 152416
rect 154726 152360 154731 152416
rect 49601 152358 154731 152360
rect 49601 152355 49667 152358
rect 154665 152355 154731 152358
rect 156689 152418 156755 152421
rect 245837 152418 245903 152421
rect 156689 152416 245903 152418
rect 156689 152360 156694 152416
rect 156750 152360 245842 152416
rect 245898 152360 245903 152416
rect 156689 152358 245903 152360
rect 156689 152355 156755 152358
rect 245837 152355 245903 152358
rect 12801 151874 12867 151877
rect 119337 151874 119403 151877
rect 12801 151872 119403 151874
rect 12801 151816 12806 151872
rect 12862 151816 119342 151872
rect 119398 151816 119403 151872
rect 12801 151814 119403 151816
rect 12801 151811 12867 151814
rect 119337 151811 119403 151814
rect 9397 151330 9463 151333
rect 23105 151330 23171 151333
rect 33501 151330 33567 151333
rect 9397 151328 16590 151330
rect 9397 151272 9402 151328
rect 9458 151272 16590 151328
rect 9397 151270 16590 151272
rect 9397 151267 9463 151270
rect 16530 150514 16590 151270
rect 23105 151328 26250 151330
rect 23105 151272 23110 151328
rect 23166 151272 26250 151328
rect 23105 151270 26250 151272
rect 23105 151267 23171 151270
rect 26190 150650 26250 151270
rect 33501 151328 35910 151330
rect 33501 151272 33506 151328
rect 33562 151272 35910 151328
rect 33501 151270 35910 151272
rect 33501 151267 33567 151270
rect 35850 150786 35910 151270
rect 531589 151194 531655 151197
rect 529828 151192 531655 151194
rect 529828 151136 531594 151192
rect 531650 151136 531655 151192
rect 529828 151134 531655 151136
rect 531589 151131 531655 151134
rect 535177 151058 535243 151061
rect 539200 151058 540000 151088
rect 535177 151056 540000 151058
rect 535177 151000 535182 151056
rect 535238 151000 540000 151056
rect 535177 150998 540000 151000
rect 535177 150995 535243 150998
rect 539200 150968 540000 150998
rect 126973 150922 127039 150925
rect 126973 150920 130180 150922
rect 126973 150864 126978 150920
rect 127034 150864 130180 150920
rect 126973 150862 130180 150864
rect 126973 150859 127039 150862
rect 119429 150786 119495 150789
rect 35850 150784 119495 150786
rect 35850 150728 119434 150784
rect 119490 150728 119495 150784
rect 35850 150726 119495 150728
rect 119429 150723 119495 150726
rect 122097 150650 122163 150653
rect 26190 150648 122163 150650
rect 26190 150592 122102 150648
rect 122158 150592 122163 150648
rect 26190 150590 122163 150592
rect 122097 150587 122163 150590
rect 126237 150514 126303 150517
rect 16530 150512 126303 150514
rect 16530 150456 126242 150512
rect 126298 150456 126303 150512
rect 16530 150454 126303 150456
rect 126237 150451 126303 150454
rect 532601 149834 532667 149837
rect 529828 149832 532667 149834
rect 529828 149776 532606 149832
rect 532662 149776 532667 149832
rect 529828 149774 532667 149776
rect 532601 149771 532667 149774
rect 534717 149562 534783 149565
rect 539200 149562 540000 149592
rect 534717 149560 540000 149562
rect 534717 149504 534722 149560
rect 534778 149504 540000 149560
rect 534717 149502 540000 149504
rect 534717 149499 534783 149502
rect 539200 149472 540000 149502
rect 126973 149018 127039 149021
rect 126973 149016 130180 149018
rect 126973 148960 126978 149016
rect 127034 148960 130180 149016
rect 126973 148958 130180 148960
rect 126973 148955 127039 148958
rect 532325 148474 532391 148477
rect 529828 148472 532391 148474
rect 529828 148416 532330 148472
rect 532386 148416 532391 148472
rect 529828 148414 532391 148416
rect 532325 148411 532391 148414
rect 534809 148066 534875 148069
rect 539200 148066 540000 148096
rect 534809 148064 540000 148066
rect 534809 148008 534814 148064
rect 534870 148008 540000 148064
rect 534809 148006 540000 148008
rect 534809 148003 534875 148006
rect 539200 147976 540000 148006
rect 126973 147114 127039 147117
rect 531957 147114 532023 147117
rect 126973 147112 130180 147114
rect 126973 147056 126978 147112
rect 127034 147056 130180 147112
rect 126973 147054 130180 147056
rect 529828 147112 532023 147114
rect 529828 147056 531962 147112
rect 532018 147056 532023 147112
rect 529828 147054 532023 147056
rect 126973 147051 127039 147054
rect 531957 147051 532023 147054
rect 535085 146570 535151 146573
rect 539200 146570 540000 146600
rect 535085 146568 540000 146570
rect 535085 146512 535090 146568
rect 535146 146512 540000 146568
rect 535085 146510 540000 146512
rect 535085 146507 535151 146510
rect 539200 146480 540000 146510
rect 116669 146162 116735 146165
rect 113804 146160 116735 146162
rect 113804 146104 116674 146160
rect 116730 146104 116735 146160
rect 113804 146102 116735 146104
rect 116669 146099 116735 146102
rect 532141 145754 532207 145757
rect 529828 145752 532207 145754
rect 529828 145696 532146 145752
rect 532202 145696 532207 145752
rect 529828 145694 532207 145696
rect 532141 145691 532207 145694
rect 126973 145210 127039 145213
rect 126973 145208 130180 145210
rect 126973 145152 126978 145208
rect 127034 145152 130180 145208
rect 126973 145150 130180 145152
rect 126973 145147 127039 145150
rect 534993 144938 535059 144941
rect 539200 144938 540000 144968
rect 534993 144936 540000 144938
rect 534993 144880 534998 144936
rect 535054 144880 540000 144936
rect 534993 144878 540000 144880
rect 534993 144875 535059 144878
rect 539200 144848 540000 144878
rect 531773 144394 531839 144397
rect 529828 144392 531839 144394
rect 529828 144336 531778 144392
rect 531834 144336 531839 144392
rect 529828 144334 531839 144336
rect 531773 144331 531839 144334
rect 536189 143442 536255 143445
rect 539200 143442 540000 143472
rect 536189 143440 540000 143442
rect 536189 143384 536194 143440
rect 536250 143384 540000 143440
rect 536189 143382 540000 143384
rect 536189 143379 536255 143382
rect 539200 143352 540000 143382
rect 126973 143306 127039 143309
rect 126973 143304 130180 143306
rect 126973 143248 126978 143304
rect 127034 143248 130180 143304
rect 126973 143246 130180 143248
rect 126973 143243 127039 143246
rect 531681 143034 531747 143037
rect 529828 143032 531747 143034
rect 529828 142976 531686 143032
rect 531742 142976 531747 143032
rect 529828 142974 531747 142976
rect 531681 142971 531747 142974
rect 536005 141946 536071 141949
rect 539200 141946 540000 141976
rect 536005 141944 540000 141946
rect 536005 141888 536010 141944
rect 536066 141888 540000 141944
rect 536005 141886 540000 141888
rect 536005 141883 536071 141886
rect 539200 141856 540000 141886
rect 531957 141674 532023 141677
rect 529828 141672 532023 141674
rect 529828 141616 531962 141672
rect 532018 141616 532023 141672
rect 529828 141614 532023 141616
rect 531957 141611 532023 141614
rect 127893 141402 127959 141405
rect 127893 141400 130180 141402
rect 127893 141344 127898 141400
rect 127954 141344 130180 141400
rect 127893 141342 130180 141344
rect 127893 141339 127959 141342
rect 536741 140450 536807 140453
rect 539200 140450 540000 140480
rect 536741 140448 540000 140450
rect 536741 140392 536746 140448
rect 536802 140392 540000 140448
rect 536741 140390 540000 140392
rect 536741 140387 536807 140390
rect 539200 140360 540000 140390
rect 531957 140314 532023 140317
rect 529828 140312 532023 140314
rect 529828 140256 531962 140312
rect 532018 140256 532023 140312
rect 529828 140254 532023 140256
rect 531957 140251 532023 140254
rect 126973 139498 127039 139501
rect 126973 139496 130180 139498
rect 126973 139440 126978 139496
rect 127034 139440 130180 139496
rect 126973 139438 130180 139440
rect 126973 139435 127039 139438
rect 531589 138954 531655 138957
rect 529828 138952 531655 138954
rect 529828 138896 531594 138952
rect 531650 138896 531655 138952
rect 529828 138894 531655 138896
rect 531589 138891 531655 138894
rect 536649 138954 536715 138957
rect 539200 138954 540000 138984
rect 536649 138952 540000 138954
rect 536649 138896 536654 138952
rect 536710 138896 540000 138952
rect 536649 138894 540000 138896
rect 536649 138891 536715 138894
rect 539200 138864 540000 138894
rect 531405 137594 531471 137597
rect 529828 137592 531471 137594
rect 529828 137536 531410 137592
rect 531466 137536 531471 137592
rect 529828 137534 531471 137536
rect 531405 137531 531471 137534
rect 126973 137458 127039 137461
rect 536557 137458 536623 137461
rect 539200 137458 540000 137488
rect 126973 137456 130180 137458
rect 126973 137400 126978 137456
rect 127034 137400 130180 137456
rect 126973 137398 130180 137400
rect 536557 137456 540000 137458
rect 536557 137400 536562 137456
rect 536618 137400 540000 137456
rect 536557 137398 540000 137400
rect 126973 137395 127039 137398
rect 536557 137395 536623 137398
rect 539200 137368 540000 137398
rect 532141 136234 532207 136237
rect 529828 136232 532207 136234
rect 529828 136176 532146 136232
rect 532202 136176 532207 136232
rect 529828 136174 532207 136176
rect 532141 136171 532207 136174
rect 536465 135826 536531 135829
rect 539200 135826 540000 135856
rect 536465 135824 540000 135826
rect 536465 135768 536470 135824
rect 536526 135768 540000 135824
rect 536465 135766 540000 135768
rect 536465 135763 536531 135766
rect 539200 135736 540000 135766
rect 126973 135554 127039 135557
rect 126973 135552 130180 135554
rect 126973 135496 126978 135552
rect 127034 135496 130180 135552
rect 126973 135494 130180 135496
rect 126973 135491 127039 135494
rect 531773 134874 531839 134877
rect 529828 134872 531839 134874
rect 529828 134816 531778 134872
rect 531834 134816 531839 134872
rect 529828 134814 531839 134816
rect 531773 134811 531839 134814
rect 116577 134738 116643 134741
rect 113804 134736 116643 134738
rect 113804 134680 116582 134736
rect 116638 134680 116643 134736
rect 113804 134678 116643 134680
rect 116577 134675 116643 134678
rect 536373 134330 536439 134333
rect 539200 134330 540000 134360
rect 536373 134328 540000 134330
rect 536373 134272 536378 134328
rect 536434 134272 540000 134328
rect 536373 134270 540000 134272
rect 536373 134267 536439 134270
rect 539200 134240 540000 134270
rect 126973 133650 127039 133653
rect 126973 133648 130180 133650
rect 126973 133592 126978 133648
rect 127034 133592 130180 133648
rect 126973 133590 130180 133592
rect 126973 133587 127039 133590
rect 531773 133378 531839 133381
rect 529828 133376 531839 133378
rect 529828 133320 531778 133376
rect 531834 133320 531839 133376
rect 529828 133318 531839 133320
rect 531773 133315 531839 133318
rect 536097 132834 536163 132837
rect 539200 132834 540000 132864
rect 536097 132832 540000 132834
rect 536097 132776 536102 132832
rect 536158 132776 540000 132832
rect 536097 132774 540000 132776
rect 536097 132771 536163 132774
rect 539200 132744 540000 132774
rect 531405 132018 531471 132021
rect 529828 132016 531471 132018
rect 529828 131960 531410 132016
rect 531466 131960 531471 132016
rect 529828 131958 531471 131960
rect 531405 131955 531471 131958
rect 126973 131746 127039 131749
rect 126973 131744 130180 131746
rect 126973 131688 126978 131744
rect 127034 131688 130180 131744
rect 126973 131686 130180 131688
rect 126973 131683 127039 131686
rect 536281 131338 536347 131341
rect 539200 131338 540000 131368
rect 536281 131336 540000 131338
rect 536281 131280 536286 131336
rect 536342 131280 540000 131336
rect 536281 131278 540000 131280
rect 536281 131275 536347 131278
rect 539200 131248 540000 131278
rect 532601 130658 532667 130661
rect 529828 130656 532667 130658
rect 529828 130600 532606 130656
rect 532662 130600 532667 130656
rect 529828 130598 532667 130600
rect 532601 130595 532667 130598
rect 126973 129842 127039 129845
rect 536189 129842 536255 129845
rect 539200 129842 540000 129872
rect 126973 129840 130180 129842
rect 126973 129784 126978 129840
rect 127034 129784 130180 129840
rect 126973 129782 130180 129784
rect 536189 129840 540000 129842
rect 536189 129784 536194 129840
rect 536250 129784 540000 129840
rect 536189 129782 540000 129784
rect 126973 129779 127039 129782
rect 536189 129779 536255 129782
rect 539200 129752 540000 129782
rect 531589 129298 531655 129301
rect 529828 129296 531655 129298
rect 529828 129240 531594 129296
rect 531650 129240 531655 129296
rect 529828 129238 531655 129240
rect 531589 129235 531655 129238
rect 536649 128346 536715 128349
rect 539200 128346 540000 128376
rect 536649 128344 540000 128346
rect 536649 128288 536654 128344
rect 536710 128288 540000 128344
rect 536649 128286 540000 128288
rect 536649 128283 536715 128286
rect 539200 128256 540000 128286
rect 126973 127938 127039 127941
rect 531957 127938 532023 127941
rect 126973 127936 130180 127938
rect 126973 127880 126978 127936
rect 127034 127880 130180 127936
rect 126973 127878 130180 127880
rect 529828 127936 532023 127938
rect 529828 127880 531962 127936
rect 532018 127880 532023 127936
rect 529828 127878 532023 127880
rect 126973 127875 127039 127878
rect 531957 127875 532023 127878
rect 536741 126714 536807 126717
rect 539200 126714 540000 126744
rect 536741 126712 540000 126714
rect 536741 126656 536746 126712
rect 536802 126656 540000 126712
rect 536741 126654 540000 126656
rect 536741 126651 536807 126654
rect 539200 126624 540000 126654
rect 531865 126578 531931 126581
rect 529828 126576 531931 126578
rect 529828 126520 531870 126576
rect 531926 126520 531931 126576
rect 529828 126518 531931 126520
rect 531865 126515 531931 126518
rect 126973 126034 127039 126037
rect 126973 126032 130180 126034
rect 126973 125976 126978 126032
rect 127034 125976 130180 126032
rect 126973 125974 130180 125976
rect 126973 125971 127039 125974
rect 532601 125218 532667 125221
rect 529828 125216 532667 125218
rect 529828 125160 532606 125216
rect 532662 125160 532667 125216
rect 529828 125158 532667 125160
rect 532601 125155 532667 125158
rect 535453 125218 535519 125221
rect 539200 125218 540000 125248
rect 535453 125216 540000 125218
rect 535453 125160 535458 125216
rect 535514 125160 540000 125216
rect 535453 125158 540000 125160
rect 535453 125155 535519 125158
rect 539200 125128 540000 125158
rect 126329 124130 126395 124133
rect 126329 124128 130180 124130
rect 126329 124072 126334 124128
rect 126390 124072 130180 124128
rect 126329 124070 130180 124072
rect 126329 124067 126395 124070
rect 531773 123858 531839 123861
rect 529828 123856 531839 123858
rect 529828 123800 531778 123856
rect 531834 123800 531839 123856
rect 529828 123798 531839 123800
rect 531773 123795 531839 123798
rect 536373 123722 536439 123725
rect 539200 123722 540000 123752
rect 536373 123720 540000 123722
rect 536373 123664 536378 123720
rect 536434 123664 540000 123720
rect 536373 123662 540000 123664
rect 536373 123659 536439 123662
rect 539200 123632 540000 123662
rect 116669 123314 116735 123317
rect 113804 123312 116735 123314
rect 113804 123256 116674 123312
rect 116730 123256 116735 123312
rect 113804 123254 116735 123256
rect 116669 123251 116735 123254
rect 532601 122498 532667 122501
rect 529828 122496 532667 122498
rect 529828 122440 532606 122496
rect 532662 122440 532667 122496
rect 529828 122438 532667 122440
rect 532601 122435 532667 122438
rect 535637 122226 535703 122229
rect 539200 122226 540000 122256
rect 535637 122224 540000 122226
rect 535637 122168 535642 122224
rect 535698 122168 540000 122224
rect 535637 122166 540000 122168
rect 535637 122163 535703 122166
rect 539200 122136 540000 122166
rect 126973 122090 127039 122093
rect 126973 122088 130180 122090
rect 126973 122032 126978 122088
rect 127034 122032 130180 122088
rect 126973 122030 130180 122032
rect 126973 122027 127039 122030
rect 532141 121138 532207 121141
rect 529828 121136 532207 121138
rect 529828 121080 532146 121136
rect 532202 121080 532207 121136
rect 529828 121078 532207 121080
rect 532141 121075 532207 121078
rect 536281 120730 536347 120733
rect 539200 120730 540000 120760
rect 536281 120728 540000 120730
rect 536281 120672 536286 120728
rect 536342 120672 540000 120728
rect 536281 120670 540000 120672
rect 536281 120667 536347 120670
rect 539200 120640 540000 120670
rect 126973 120186 127039 120189
rect 126973 120184 130180 120186
rect 126973 120128 126978 120184
rect 127034 120128 130180 120184
rect 126973 120126 130180 120128
rect 126973 120123 127039 120126
rect 532509 119778 532575 119781
rect 529828 119776 532575 119778
rect 529828 119720 532514 119776
rect 532570 119720 532575 119776
rect 529828 119718 532575 119720
rect 532509 119715 532575 119718
rect 536465 119234 536531 119237
rect 539200 119234 540000 119264
rect 536465 119232 540000 119234
rect 536465 119176 536470 119232
rect 536526 119176 540000 119232
rect 536465 119174 540000 119176
rect 536465 119171 536531 119174
rect 539200 119144 540000 119174
rect 532601 118418 532667 118421
rect 529828 118416 532667 118418
rect 529828 118360 532606 118416
rect 532662 118360 532667 118416
rect 529828 118358 532667 118360
rect 532601 118355 532667 118358
rect 126973 118282 127039 118285
rect 126973 118280 130180 118282
rect 126973 118224 126978 118280
rect 127034 118224 130180 118280
rect 126973 118222 130180 118224
rect 126973 118219 127039 118222
rect 536189 117602 536255 117605
rect 539200 117602 540000 117632
rect 536189 117600 540000 117602
rect 536189 117544 536194 117600
rect 536250 117544 540000 117600
rect 536189 117542 540000 117544
rect 536189 117539 536255 117542
rect 539200 117512 540000 117542
rect 532325 117058 532391 117061
rect 529828 117056 532391 117058
rect 529828 117000 532330 117056
rect 532386 117000 532391 117056
rect 529828 116998 532391 117000
rect 532325 116995 532391 116998
rect 126973 116378 127039 116381
rect 126973 116376 130180 116378
rect 126973 116320 126978 116376
rect 127034 116320 130180 116376
rect 126973 116318 130180 116320
rect 126973 116315 127039 116318
rect 536649 116106 536715 116109
rect 539200 116106 540000 116136
rect 536649 116104 540000 116106
rect 536649 116048 536654 116104
rect 536710 116048 540000 116104
rect 536649 116046 540000 116048
rect 536649 116043 536715 116046
rect 539200 116016 540000 116046
rect 532601 115698 532667 115701
rect 529828 115696 532667 115698
rect 529828 115640 532606 115696
rect 532662 115640 532667 115696
rect 529828 115638 532667 115640
rect 532601 115635 532667 115638
rect 535545 114610 535611 114613
rect 539200 114610 540000 114640
rect 535545 114608 540000 114610
rect 535545 114552 535550 114608
rect 535606 114552 540000 114608
rect 535545 114550 540000 114552
rect 535545 114547 535611 114550
rect 539200 114520 540000 114550
rect 127709 114474 127775 114477
rect 127709 114472 130180 114474
rect 127709 114416 127714 114472
rect 127770 114416 130180 114472
rect 127709 114414 130180 114416
rect 127709 114411 127775 114414
rect 531681 114202 531747 114205
rect 529828 114200 531747 114202
rect 529828 114144 531686 114200
rect 531742 114144 531747 114200
rect 529828 114142 531747 114144
rect 531681 114139 531747 114142
rect 535453 113114 535519 113117
rect 539200 113114 540000 113144
rect 535453 113112 540000 113114
rect 535453 113056 535458 113112
rect 535514 113056 540000 113112
rect 535453 113054 540000 113056
rect 535453 113051 535519 113054
rect 539200 113024 540000 113054
rect 531773 112842 531839 112845
rect 529828 112840 531839 112842
rect 529828 112784 531778 112840
rect 531834 112784 531839 112840
rect 529828 112782 531839 112784
rect 531773 112779 531839 112782
rect 126973 112570 127039 112573
rect 126973 112568 130180 112570
rect 126973 112512 126978 112568
rect 127034 112512 130180 112568
rect 126973 112510 130180 112512
rect 126973 112507 127039 112510
rect 116761 112026 116827 112029
rect 113804 112024 116827 112026
rect 113804 111968 116766 112024
rect 116822 111968 116827 112024
rect 113804 111966 116827 111968
rect 116761 111963 116827 111966
rect 535453 111618 535519 111621
rect 539200 111618 540000 111648
rect 535453 111616 540000 111618
rect 535453 111560 535458 111616
rect 535514 111560 540000 111616
rect 535453 111558 540000 111560
rect 535453 111555 535519 111558
rect 539200 111528 540000 111558
rect 532601 111482 532667 111485
rect 529828 111480 532667 111482
rect 529828 111424 532606 111480
rect 532662 111424 532667 111480
rect 529828 111422 532667 111424
rect 532601 111419 532667 111422
rect 126973 110666 127039 110669
rect 126973 110664 130180 110666
rect 126973 110608 126978 110664
rect 127034 110608 130180 110664
rect 126973 110606 130180 110608
rect 126973 110603 127039 110606
rect 531957 110122 532023 110125
rect 529828 110120 532023 110122
rect 529828 110064 531962 110120
rect 532018 110064 532023 110120
rect 529828 110062 532023 110064
rect 531957 110059 532023 110062
rect 535453 110122 535519 110125
rect 539200 110122 540000 110152
rect 535453 110120 540000 110122
rect 535453 110064 535458 110120
rect 535514 110064 540000 110120
rect 535453 110062 540000 110064
rect 535453 110059 535519 110062
rect 539200 110032 540000 110062
rect 126973 108762 127039 108765
rect 531773 108762 531839 108765
rect 126973 108760 130180 108762
rect 126973 108704 126978 108760
rect 127034 108704 130180 108760
rect 126973 108702 130180 108704
rect 529828 108760 531839 108762
rect 529828 108704 531778 108760
rect 531834 108704 531839 108760
rect 529828 108702 531839 108704
rect 126973 108699 127039 108702
rect 531773 108699 531839 108702
rect 535453 108490 535519 108493
rect 539200 108490 540000 108520
rect 535453 108488 540000 108490
rect 535453 108432 535458 108488
rect 535514 108432 540000 108488
rect 535453 108430 540000 108432
rect 535453 108427 535519 108430
rect 539200 108400 540000 108430
rect 531773 107402 531839 107405
rect 529828 107400 531839 107402
rect 529828 107344 531778 107400
rect 531834 107344 531839 107400
rect 529828 107342 531839 107344
rect 531773 107339 531839 107342
rect 535453 106994 535519 106997
rect 539200 106994 540000 107024
rect 535453 106992 540000 106994
rect 535453 106936 535458 106992
rect 535514 106936 540000 106992
rect 535453 106934 540000 106936
rect 535453 106931 535519 106934
rect 539200 106904 540000 106934
rect 126973 106722 127039 106725
rect 126973 106720 130180 106722
rect 126973 106664 126978 106720
rect 127034 106664 130180 106720
rect 126973 106662 130180 106664
rect 126973 106659 127039 106662
rect 532509 106042 532575 106045
rect 529828 106040 532575 106042
rect 529828 105984 532514 106040
rect 532570 105984 532575 106040
rect 529828 105982 532575 105984
rect 532509 105979 532575 105982
rect 535453 105498 535519 105501
rect 539200 105498 540000 105528
rect 535453 105496 540000 105498
rect 535453 105440 535458 105496
rect 535514 105440 540000 105496
rect 535453 105438 540000 105440
rect 535453 105435 535519 105438
rect 539200 105408 540000 105438
rect 126973 104818 127039 104821
rect 126973 104816 130180 104818
rect 126973 104760 126978 104816
rect 127034 104760 130180 104816
rect 126973 104758 130180 104760
rect 126973 104755 127039 104758
rect 532601 104682 532667 104685
rect 529828 104680 532667 104682
rect 529828 104624 532606 104680
rect 532662 104624 532667 104680
rect 529828 104622 532667 104624
rect 532601 104619 532667 104622
rect 535453 104002 535519 104005
rect 539200 104002 540000 104032
rect 535453 104000 540000 104002
rect 535453 103944 535458 104000
rect 535514 103944 540000 104000
rect 535453 103942 540000 103944
rect 535453 103939 535519 103942
rect 539200 103912 540000 103942
rect 532417 103322 532483 103325
rect 529828 103320 532483 103322
rect 529828 103264 532422 103320
rect 532478 103264 532483 103320
rect 529828 103262 532483 103264
rect 532417 103259 532483 103262
rect 126973 102914 127039 102917
rect 126973 102912 130180 102914
rect 126973 102856 126978 102912
rect 127034 102856 130180 102912
rect 126973 102854 130180 102856
rect 126973 102851 127039 102854
rect 535453 102506 535519 102509
rect 539200 102506 540000 102536
rect 535453 102504 540000 102506
rect 535453 102448 535458 102504
rect 535514 102448 540000 102504
rect 535453 102446 540000 102448
rect 535453 102443 535519 102446
rect 539200 102416 540000 102446
rect 532233 101962 532299 101965
rect 529828 101960 532299 101962
rect 529828 101904 532238 101960
rect 532294 101904 532299 101960
rect 529828 101902 532299 101904
rect 532233 101899 532299 101902
rect 126973 101010 127039 101013
rect 535453 101010 535519 101013
rect 539200 101010 540000 101040
rect 126973 101008 130180 101010
rect 126973 100952 126978 101008
rect 127034 100952 130180 101008
rect 126973 100950 130180 100952
rect 535453 101008 540000 101010
rect 535453 100952 535458 101008
rect 535514 100952 540000 101008
rect 535453 100950 540000 100952
rect 126973 100947 127039 100950
rect 535453 100947 535519 100950
rect 539200 100920 540000 100950
rect 116945 100602 117011 100605
rect 532141 100602 532207 100605
rect 113804 100600 117011 100602
rect 113804 100544 116950 100600
rect 117006 100544 117011 100600
rect 113804 100542 117011 100544
rect 529828 100600 532207 100602
rect 529828 100544 532146 100600
rect 532202 100544 532207 100600
rect 529828 100542 532207 100544
rect 116945 100539 117011 100542
rect 532141 100539 532207 100542
rect 535453 99378 535519 99381
rect 539200 99378 540000 99408
rect 535453 99376 540000 99378
rect 535453 99320 535458 99376
rect 535514 99320 540000 99376
rect 535453 99318 540000 99320
rect 535453 99315 535519 99318
rect 539200 99288 540000 99318
rect 532233 99242 532299 99245
rect 529828 99240 532299 99242
rect 529828 99184 532238 99240
rect 532294 99184 532299 99240
rect 529828 99182 532299 99184
rect 532233 99179 532299 99182
rect 126973 99106 127039 99109
rect 126973 99104 130180 99106
rect 126973 99048 126978 99104
rect 127034 99048 130180 99104
rect 126973 99046 130180 99048
rect 126973 99043 127039 99046
rect 532417 97882 532483 97885
rect 529828 97880 532483 97882
rect 529828 97824 532422 97880
rect 532478 97824 532483 97880
rect 529828 97822 532483 97824
rect 532417 97819 532483 97822
rect 535453 97882 535519 97885
rect 539200 97882 540000 97912
rect 535453 97880 540000 97882
rect 535453 97824 535458 97880
rect 535514 97824 540000 97880
rect 535453 97822 540000 97824
rect 535453 97819 535519 97822
rect 539200 97792 540000 97822
rect 126973 97202 127039 97205
rect 126973 97200 130180 97202
rect 126973 97144 126978 97200
rect 127034 97144 130180 97200
rect 126973 97142 130180 97144
rect 126973 97139 127039 97142
rect 532049 96386 532115 96389
rect 529828 96384 532115 96386
rect 529828 96328 532054 96384
rect 532110 96328 532115 96384
rect 529828 96326 532115 96328
rect 532049 96323 532115 96326
rect 535453 96386 535519 96389
rect 539200 96386 540000 96416
rect 535453 96384 540000 96386
rect 535453 96328 535458 96384
rect 535514 96328 540000 96384
rect 535453 96326 540000 96328
rect 535453 96323 535519 96326
rect 539200 96296 540000 96326
rect 126973 95298 127039 95301
rect 126973 95296 130180 95298
rect 126973 95240 126978 95296
rect 127034 95240 130180 95296
rect 126973 95238 130180 95240
rect 126973 95235 127039 95238
rect 532601 95026 532667 95029
rect 529828 95024 532667 95026
rect 529828 94968 532606 95024
rect 532662 94968 532667 95024
rect 529828 94966 532667 94968
rect 532601 94963 532667 94966
rect 535453 94890 535519 94893
rect 539200 94890 540000 94920
rect 535453 94888 540000 94890
rect 535453 94832 535458 94888
rect 535514 94832 540000 94888
rect 535453 94830 540000 94832
rect 535453 94827 535519 94830
rect 539200 94800 540000 94830
rect 532233 93666 532299 93669
rect 529828 93664 532299 93666
rect 529828 93608 532238 93664
rect 532294 93608 532299 93664
rect 529828 93606 532299 93608
rect 532233 93603 532299 93606
rect 535453 93394 535519 93397
rect 539200 93394 540000 93424
rect 535453 93392 540000 93394
rect 535453 93336 535458 93392
rect 535514 93336 540000 93392
rect 535453 93334 540000 93336
rect 535453 93331 535519 93334
rect 539200 93304 540000 93334
rect 126237 93258 126303 93261
rect 126237 93256 130180 93258
rect 126237 93200 126242 93256
rect 126298 93200 130180 93256
rect 126237 93198 130180 93200
rect 126237 93195 126303 93198
rect 532141 92306 532207 92309
rect 529828 92304 532207 92306
rect 529828 92248 532146 92304
rect 532202 92248 532207 92304
rect 529828 92246 532207 92248
rect 532141 92243 532207 92246
rect 535453 91898 535519 91901
rect 539200 91898 540000 91928
rect 535453 91896 540000 91898
rect 535453 91840 535458 91896
rect 535514 91840 540000 91896
rect 535453 91838 540000 91840
rect 535453 91835 535519 91838
rect 539200 91808 540000 91838
rect 127617 91354 127683 91357
rect 127617 91352 130180 91354
rect 127617 91296 127622 91352
rect 127678 91296 130180 91352
rect 127617 91294 130180 91296
rect 127617 91291 127683 91294
rect 532049 90946 532115 90949
rect 529828 90944 532115 90946
rect 529828 90888 532054 90944
rect 532110 90888 532115 90944
rect 529828 90886 532115 90888
rect 532049 90883 532115 90886
rect 535453 90266 535519 90269
rect 539200 90266 540000 90296
rect 535453 90264 540000 90266
rect 535453 90208 535458 90264
rect 535514 90208 540000 90264
rect 535453 90206 540000 90208
rect 535453 90203 535519 90206
rect 539200 90176 540000 90206
rect 532509 89586 532575 89589
rect 529828 89584 532575 89586
rect 529828 89528 532514 89584
rect 532570 89528 532575 89584
rect 529828 89526 532575 89528
rect 532509 89523 532575 89526
rect 126973 89450 127039 89453
rect 126973 89448 130180 89450
rect 126973 89392 126978 89448
rect 127034 89392 130180 89448
rect 126973 89390 130180 89392
rect 126973 89387 127039 89390
rect 115933 89178 115999 89181
rect 113804 89176 115999 89178
rect 113804 89120 115938 89176
rect 115994 89120 115999 89176
rect 113804 89118 115999 89120
rect 115933 89115 115999 89118
rect 535453 88770 535519 88773
rect 539200 88770 540000 88800
rect 535453 88768 540000 88770
rect 535453 88712 535458 88768
rect 535514 88712 540000 88768
rect 535453 88710 540000 88712
rect 535453 88707 535519 88710
rect 539200 88680 540000 88710
rect 532417 88226 532483 88229
rect 529828 88224 532483 88226
rect 529828 88168 532422 88224
rect 532478 88168 532483 88224
rect 529828 88166 532483 88168
rect 532417 88163 532483 88166
rect 126973 87546 127039 87549
rect 126973 87544 130180 87546
rect 126973 87488 126978 87544
rect 127034 87488 130180 87544
rect 126973 87486 130180 87488
rect 126973 87483 127039 87486
rect 535453 87274 535519 87277
rect 539200 87274 540000 87304
rect 535453 87272 540000 87274
rect 535453 87216 535458 87272
rect 535514 87216 540000 87272
rect 535453 87214 540000 87216
rect 535453 87211 535519 87214
rect 539200 87184 540000 87214
rect 531957 86866 532023 86869
rect 529828 86864 532023 86866
rect 529828 86808 531962 86864
rect 532018 86808 532023 86864
rect 529828 86806 532023 86808
rect 531957 86803 532023 86806
rect 535453 85778 535519 85781
rect 539200 85778 540000 85808
rect 535453 85776 540000 85778
rect 535453 85720 535458 85776
rect 535514 85720 540000 85776
rect 535453 85718 540000 85720
rect 535453 85715 535519 85718
rect 539200 85688 540000 85718
rect 126973 85642 127039 85645
rect 126973 85640 130180 85642
rect 126973 85584 126978 85640
rect 127034 85584 130180 85640
rect 126973 85582 130180 85584
rect 126973 85579 127039 85582
rect 532601 85506 532667 85509
rect 529828 85504 532667 85506
rect 529828 85448 532606 85504
rect 532662 85448 532667 85504
rect 529828 85446 532667 85448
rect 532601 85443 532667 85446
rect 535453 84282 535519 84285
rect 539200 84282 540000 84312
rect 535453 84280 540000 84282
rect 535453 84224 535458 84280
rect 535514 84224 540000 84280
rect 535453 84222 540000 84224
rect 535453 84219 535519 84222
rect 539200 84192 540000 84222
rect 532049 84146 532115 84149
rect 529828 84144 532115 84146
rect 529828 84088 532054 84144
rect 532110 84088 532115 84144
rect 529828 84086 532115 84088
rect 532049 84083 532115 84086
rect 126973 83738 127039 83741
rect 126973 83736 130180 83738
rect 126973 83680 126978 83736
rect 127034 83680 130180 83736
rect 126973 83678 130180 83680
rect 126973 83675 127039 83678
rect 532325 82786 532391 82789
rect 529828 82784 532391 82786
rect 529828 82728 532330 82784
rect 532386 82728 532391 82784
rect 529828 82726 532391 82728
rect 532325 82723 532391 82726
rect 535637 82786 535703 82789
rect 539200 82786 540000 82816
rect 535637 82784 540000 82786
rect 535637 82728 535642 82784
rect 535698 82728 540000 82784
rect 535637 82726 540000 82728
rect 535637 82723 535703 82726
rect 539200 82696 540000 82726
rect 126973 81834 127039 81837
rect 126973 81832 130180 81834
rect 126973 81776 126978 81832
rect 127034 81776 130180 81832
rect 126973 81774 130180 81776
rect 126973 81771 127039 81774
rect 532509 81426 532575 81429
rect 529828 81424 532575 81426
rect 529828 81368 532514 81424
rect 532570 81368 532575 81424
rect 529828 81366 532575 81368
rect 532509 81363 532575 81366
rect 535545 81154 535611 81157
rect 539200 81154 540000 81184
rect 535545 81152 540000 81154
rect 535545 81096 535550 81152
rect 535606 81096 540000 81152
rect 535545 81094 540000 81096
rect 535545 81091 535611 81094
rect 539200 81064 540000 81094
rect 532601 80066 532667 80069
rect 529828 80064 532667 80066
rect 529828 80008 532606 80064
rect 532662 80008 532667 80064
rect 529828 80006 532667 80008
rect 532601 80003 532667 80006
rect 126973 79930 127039 79933
rect 126973 79928 130180 79930
rect 126973 79872 126978 79928
rect 127034 79872 130180 79928
rect 126973 79870 130180 79872
rect 126973 79867 127039 79870
rect 535453 79658 535519 79661
rect 539200 79658 540000 79688
rect 535453 79656 540000 79658
rect 535453 79600 535458 79656
rect 535514 79600 540000 79656
rect 535453 79598 540000 79600
rect 535453 79595 535519 79598
rect 539200 79568 540000 79598
rect 532141 78706 532207 78709
rect 529828 78704 532207 78706
rect 529828 78648 532146 78704
rect 532202 78648 532207 78704
rect 529828 78646 532207 78648
rect 532141 78643 532207 78646
rect 536281 78162 536347 78165
rect 539200 78162 540000 78192
rect 536281 78160 540000 78162
rect 536281 78104 536286 78160
rect 536342 78104 540000 78160
rect 536281 78102 540000 78104
rect 536281 78099 536347 78102
rect 539200 78072 540000 78102
rect 116117 77890 116183 77893
rect 113804 77888 116183 77890
rect 113804 77832 116122 77888
rect 116178 77832 116183 77888
rect 113804 77830 116183 77832
rect 116117 77827 116183 77830
rect 126973 77890 127039 77893
rect 126973 77888 130180 77890
rect 126973 77832 126978 77888
rect 127034 77832 130180 77888
rect 126973 77830 130180 77832
rect 126973 77827 127039 77830
rect 532601 77210 532667 77213
rect 529828 77208 532667 77210
rect 529828 77152 532606 77208
rect 532662 77152 532667 77208
rect 529828 77150 532667 77152
rect 532601 77147 532667 77150
rect 535545 76666 535611 76669
rect 539200 76666 540000 76696
rect 535545 76664 540000 76666
rect 535545 76608 535550 76664
rect 535606 76608 540000 76664
rect 535545 76606 540000 76608
rect 535545 76603 535611 76606
rect 539200 76576 540000 76606
rect 126973 75986 127039 75989
rect 126973 75984 130180 75986
rect 126973 75928 126978 75984
rect 127034 75928 130180 75984
rect 126973 75926 130180 75928
rect 126973 75923 127039 75926
rect 532601 75850 532667 75853
rect 529828 75848 532667 75850
rect 529828 75792 532606 75848
rect 532662 75792 532667 75848
rect 529828 75790 532667 75792
rect 532601 75787 532667 75790
rect 535637 75170 535703 75173
rect 539200 75170 540000 75200
rect 535637 75168 540000 75170
rect 535637 75112 535642 75168
rect 535698 75112 540000 75168
rect 535637 75110 540000 75112
rect 535637 75107 535703 75110
rect 539200 75080 540000 75110
rect 532601 74490 532667 74493
rect 529828 74488 532667 74490
rect 529828 74432 532606 74488
rect 532662 74432 532667 74488
rect 529828 74430 532667 74432
rect 532601 74427 532667 74430
rect 126973 74082 127039 74085
rect 126973 74080 130180 74082
rect 126973 74024 126978 74080
rect 127034 74024 130180 74080
rect 126973 74022 130180 74024
rect 126973 74019 127039 74022
rect 535729 73674 535795 73677
rect 539200 73674 540000 73704
rect 535729 73672 540000 73674
rect 535729 73616 535734 73672
rect 535790 73616 540000 73672
rect 535729 73614 540000 73616
rect 535729 73611 535795 73614
rect 539200 73584 540000 73614
rect 532417 73130 532483 73133
rect 529828 73128 532483 73130
rect 529828 73072 532422 73128
rect 532478 73072 532483 73128
rect 529828 73070 532483 73072
rect 532417 73067 532483 73070
rect 126973 72178 127039 72181
rect 126973 72176 130180 72178
rect 126973 72120 126978 72176
rect 127034 72120 130180 72176
rect 126973 72118 130180 72120
rect 126973 72115 127039 72118
rect 535545 72042 535611 72045
rect 539200 72042 540000 72072
rect 535545 72040 540000 72042
rect 535545 71984 535550 72040
rect 535606 71984 540000 72040
rect 535545 71982 540000 71984
rect 535545 71979 535611 71982
rect 539200 71952 540000 71982
rect 532417 71770 532483 71773
rect 529828 71768 532483 71770
rect 529828 71712 532422 71768
rect 532478 71712 532483 71768
rect 529828 71710 532483 71712
rect 532417 71707 532483 71710
rect 535453 70546 535519 70549
rect 539200 70546 540000 70576
rect 535453 70544 540000 70546
rect 535453 70488 535458 70544
rect 535514 70488 540000 70544
rect 535453 70486 540000 70488
rect 535453 70483 535519 70486
rect 539200 70456 540000 70486
rect 531773 70410 531839 70413
rect 529828 70408 531839 70410
rect 529828 70352 531778 70408
rect 531834 70352 531839 70408
rect 529828 70350 531839 70352
rect 531773 70347 531839 70350
rect 126973 70274 127039 70277
rect 126973 70272 130180 70274
rect 126973 70216 126978 70272
rect 127034 70216 130180 70272
rect 126973 70214 130180 70216
rect 126973 70211 127039 70214
rect 531957 69050 532023 69053
rect 529828 69048 532023 69050
rect 529828 68992 531962 69048
rect 532018 68992 532023 69048
rect 529828 68990 532023 68992
rect 531957 68987 532023 68990
rect 535545 69050 535611 69053
rect 539200 69050 540000 69080
rect 535545 69048 540000 69050
rect 535545 68992 535550 69048
rect 535606 68992 540000 69048
rect 535545 68990 540000 68992
rect 535545 68987 535611 68990
rect 539200 68960 540000 68990
rect 126973 68370 127039 68373
rect 126973 68368 130180 68370
rect 126973 68312 126978 68368
rect 127034 68312 130180 68368
rect 126973 68310 130180 68312
rect 126973 68307 127039 68310
rect 531957 67690 532023 67693
rect 529828 67688 532023 67690
rect 529828 67632 531962 67688
rect 532018 67632 532023 67688
rect 529828 67630 532023 67632
rect 531957 67627 532023 67630
rect 535453 67554 535519 67557
rect 539200 67554 540000 67584
rect 535453 67552 540000 67554
rect 535453 67496 535458 67552
rect 535514 67496 540000 67552
rect 535453 67494 540000 67496
rect 535453 67491 535519 67494
rect 539200 67464 540000 67494
rect 116577 66466 116643 66469
rect 113804 66464 116643 66466
rect 113804 66408 116582 66464
rect 116638 66408 116643 66464
rect 113804 66406 116643 66408
rect 116577 66403 116643 66406
rect 127433 66466 127499 66469
rect 127433 66464 130180 66466
rect 127433 66408 127438 66464
rect 127494 66408 130180 66464
rect 127433 66406 130180 66408
rect 127433 66403 127499 66406
rect 531957 66330 532023 66333
rect 529828 66328 532023 66330
rect 529828 66272 531962 66328
rect 532018 66272 532023 66328
rect 529828 66270 532023 66272
rect 531957 66267 532023 66270
rect 535453 66058 535519 66061
rect 539200 66058 540000 66088
rect 535453 66056 540000 66058
rect 535453 66000 535458 66056
rect 535514 66000 540000 66056
rect 535453 65998 540000 66000
rect 535453 65995 535519 65998
rect 539200 65968 540000 65998
rect 532141 64970 532207 64973
rect 529828 64968 532207 64970
rect 529828 64912 532146 64968
rect 532202 64912 532207 64968
rect 529828 64910 532207 64912
rect 532141 64907 532207 64910
rect 126973 64562 127039 64565
rect 535453 64562 535519 64565
rect 539200 64562 540000 64592
rect 126973 64560 130180 64562
rect 126973 64504 126978 64560
rect 127034 64504 130180 64560
rect 126973 64502 130180 64504
rect 535453 64560 540000 64562
rect 535453 64504 535458 64560
rect 535514 64504 540000 64560
rect 535453 64502 540000 64504
rect 126973 64499 127039 64502
rect 535453 64499 535519 64502
rect 539200 64472 540000 64502
rect 531313 63610 531379 63613
rect 529828 63608 531379 63610
rect 529828 63552 531318 63608
rect 531374 63552 531379 63608
rect 529828 63550 531379 63552
rect 531313 63547 531379 63550
rect 535453 62930 535519 62933
rect 539200 62930 540000 62960
rect 535453 62928 540000 62930
rect 535453 62872 535458 62928
rect 535514 62872 540000 62928
rect 535453 62870 540000 62872
rect 535453 62867 535519 62870
rect 539200 62840 540000 62870
rect 126973 62522 127039 62525
rect 126973 62520 130180 62522
rect 126973 62464 126978 62520
rect 127034 62464 130180 62520
rect 126973 62462 130180 62464
rect 126973 62459 127039 62462
rect 532141 62250 532207 62253
rect 529828 62248 532207 62250
rect 529828 62192 532146 62248
rect 532202 62192 532207 62248
rect 529828 62190 532207 62192
rect 532141 62187 532207 62190
rect 535453 61434 535519 61437
rect 539200 61434 540000 61464
rect 535453 61432 540000 61434
rect 535453 61376 535458 61432
rect 535514 61376 540000 61432
rect 535453 61374 540000 61376
rect 535453 61371 535519 61374
rect 539200 61344 540000 61374
rect 532325 60890 532391 60893
rect 529828 60888 532391 60890
rect 529828 60832 532330 60888
rect 532386 60832 532391 60888
rect 529828 60830 532391 60832
rect 532325 60827 532391 60830
rect 126973 60618 127039 60621
rect 126973 60616 130180 60618
rect 126973 60560 126978 60616
rect 127034 60560 130180 60616
rect 126973 60558 130180 60560
rect 126973 60555 127039 60558
rect 535453 59938 535519 59941
rect 539200 59938 540000 59968
rect 535453 59936 540000 59938
rect 535453 59880 535458 59936
rect 535514 59880 540000 59936
rect 535453 59878 540000 59880
rect 535453 59875 535519 59878
rect 539200 59848 540000 59878
rect 532509 59394 532575 59397
rect 529828 59392 532575 59394
rect 529828 59336 532514 59392
rect 532570 59336 532575 59392
rect 529828 59334 532575 59336
rect 532509 59331 532575 59334
rect 127801 58714 127867 58717
rect 127801 58712 130180 58714
rect 127801 58656 127806 58712
rect 127862 58656 130180 58712
rect 127801 58654 130180 58656
rect 127801 58651 127867 58654
rect 535453 58442 535519 58445
rect 539200 58442 540000 58472
rect 535453 58440 540000 58442
rect 535453 58384 535458 58440
rect 535514 58384 540000 58440
rect 535453 58382 540000 58384
rect 535453 58379 535519 58382
rect 539200 58352 540000 58382
rect 532601 58034 532667 58037
rect 529828 58032 532667 58034
rect 529828 57976 532606 58032
rect 532662 57976 532667 58032
rect 529828 57974 532667 57976
rect 532601 57971 532667 57974
rect 535453 56946 535519 56949
rect 539200 56946 540000 56976
rect 535453 56944 540000 56946
rect 535453 56888 535458 56944
rect 535514 56888 540000 56944
rect 535453 56886 540000 56888
rect 535453 56883 535519 56886
rect 539200 56856 540000 56886
rect 127617 56810 127683 56813
rect 127617 56808 130180 56810
rect 127617 56752 127622 56808
rect 127678 56752 130180 56808
rect 127617 56750 130180 56752
rect 127617 56747 127683 56750
rect 532417 56674 532483 56677
rect 529828 56672 532483 56674
rect 529828 56616 532422 56672
rect 532478 56616 532483 56672
rect 529828 56614 532483 56616
rect 532417 56611 532483 56614
rect 535453 55450 535519 55453
rect 539200 55450 540000 55480
rect 535453 55448 540000 55450
rect 535453 55392 535458 55448
rect 535514 55392 540000 55448
rect 535453 55390 540000 55392
rect 535453 55387 535519 55390
rect 539200 55360 540000 55390
rect 532601 55314 532667 55317
rect 529828 55312 532667 55314
rect 529828 55256 532606 55312
rect 532662 55256 532667 55312
rect 529828 55254 532667 55256
rect 532601 55251 532667 55254
rect 116761 55042 116827 55045
rect 113804 55040 116827 55042
rect 113804 54984 116766 55040
rect 116822 54984 116827 55040
rect 113804 54982 116827 54984
rect 116761 54979 116827 54982
rect 126973 54906 127039 54909
rect 126973 54904 130180 54906
rect 126973 54848 126978 54904
rect 127034 54848 130180 54904
rect 126973 54846 130180 54848
rect 126973 54843 127039 54846
rect 531313 53954 531379 53957
rect 529828 53952 531379 53954
rect 529828 53896 531318 53952
rect 531374 53896 531379 53952
rect 529828 53894 531379 53896
rect 531313 53891 531379 53894
rect 535453 53818 535519 53821
rect 539200 53818 540000 53848
rect 535453 53816 540000 53818
rect 535453 53760 535458 53816
rect 535514 53760 540000 53816
rect 535453 53758 540000 53760
rect 535453 53755 535519 53758
rect 539200 53728 540000 53758
rect 127709 53002 127775 53005
rect 127709 53000 130180 53002
rect 127709 52944 127714 53000
rect 127770 52944 130180 53000
rect 127709 52942 130180 52944
rect 127709 52939 127775 52942
rect 532141 52594 532207 52597
rect 529828 52592 532207 52594
rect 529828 52536 532146 52592
rect 532202 52536 532207 52592
rect 529828 52534 532207 52536
rect 532141 52531 532207 52534
rect 535453 52322 535519 52325
rect 539200 52322 540000 52352
rect 535453 52320 540000 52322
rect 535453 52264 535458 52320
rect 535514 52264 540000 52320
rect 535453 52262 540000 52264
rect 535453 52259 535519 52262
rect 539200 52232 540000 52262
rect 532601 51234 532667 51237
rect 529828 51232 532667 51234
rect 529828 51176 532606 51232
rect 532662 51176 532667 51232
rect 529828 51174 532667 51176
rect 532601 51171 532667 51174
rect 126973 51098 127039 51101
rect 126973 51096 130180 51098
rect 126973 51040 126978 51096
rect 127034 51040 130180 51096
rect 126973 51038 130180 51040
rect 126973 51035 127039 51038
rect 535453 50826 535519 50829
rect 539200 50826 540000 50856
rect 535453 50824 540000 50826
rect 535453 50768 535458 50824
rect 535514 50768 540000 50824
rect 535453 50766 540000 50768
rect 535453 50763 535519 50766
rect 539200 50736 540000 50766
rect 532509 49874 532575 49877
rect 529828 49872 532575 49874
rect 529828 49816 532514 49872
rect 532570 49816 532575 49872
rect 529828 49814 532575 49816
rect 532509 49811 532575 49814
rect 535453 49330 535519 49333
rect 539200 49330 540000 49360
rect 535453 49328 540000 49330
rect 535453 49272 535458 49328
rect 535514 49272 540000 49328
rect 535453 49270 540000 49272
rect 535453 49267 535519 49270
rect 539200 49240 540000 49270
rect 126237 49058 126303 49061
rect 126237 49056 130180 49058
rect 126237 49000 126242 49056
rect 126298 49000 130180 49056
rect 126237 48998 130180 49000
rect 126237 48995 126303 48998
rect 531957 48514 532023 48517
rect 529828 48512 532023 48514
rect 529828 48456 531962 48512
rect 532018 48456 532023 48512
rect 529828 48454 532023 48456
rect 531957 48451 532023 48454
rect 535453 47834 535519 47837
rect 539200 47834 540000 47864
rect 535453 47832 540000 47834
rect 535453 47776 535458 47832
rect 535514 47776 540000 47832
rect 535453 47774 540000 47776
rect 535453 47771 535519 47774
rect 539200 47744 540000 47774
rect 126973 47154 127039 47157
rect 532601 47154 532667 47157
rect 126973 47152 130180 47154
rect 126973 47096 126978 47152
rect 127034 47096 130180 47152
rect 126973 47094 130180 47096
rect 529828 47152 532667 47154
rect 529828 47096 532606 47152
rect 532662 47096 532667 47152
rect 529828 47094 532667 47096
rect 126973 47091 127039 47094
rect 532601 47091 532667 47094
rect 535453 46338 535519 46341
rect 539200 46338 540000 46368
rect 535453 46336 540000 46338
rect 535453 46280 535458 46336
rect 535514 46280 540000 46336
rect 535453 46278 540000 46280
rect 535453 46275 535519 46278
rect 539200 46248 540000 46278
rect 532601 45794 532667 45797
rect 529828 45792 532667 45794
rect 529828 45736 532606 45792
rect 532662 45736 532667 45792
rect 529828 45734 532667 45736
rect 532601 45731 532667 45734
rect 126973 45250 127039 45253
rect 126973 45248 130180 45250
rect 126973 45192 126978 45248
rect 127034 45192 130180 45248
rect 126973 45190 130180 45192
rect 126973 45187 127039 45190
rect 535453 44706 535519 44709
rect 539200 44706 540000 44736
rect 535453 44704 540000 44706
rect 535453 44648 535458 44704
rect 535514 44648 540000 44704
rect 535453 44646 540000 44648
rect 535453 44643 535519 44646
rect 539200 44616 540000 44646
rect 532509 44434 532575 44437
rect 529828 44432 532575 44434
rect 529828 44376 532514 44432
rect 532570 44376 532575 44432
rect 529828 44374 532575 44376
rect 532509 44371 532575 44374
rect 116669 43754 116735 43757
rect 113804 43752 116735 43754
rect 113804 43696 116674 43752
rect 116730 43696 116735 43752
rect 113804 43694 116735 43696
rect 116669 43691 116735 43694
rect 126973 43346 127039 43349
rect 126973 43344 130180 43346
rect 126973 43288 126978 43344
rect 127034 43288 130180 43344
rect 126973 43286 130180 43288
rect 126973 43283 127039 43286
rect 535453 43210 535519 43213
rect 539200 43210 540000 43240
rect 535453 43208 540000 43210
rect 535453 43152 535458 43208
rect 535514 43152 540000 43208
rect 535453 43150 540000 43152
rect 535453 43147 535519 43150
rect 539200 43120 540000 43150
rect 532601 43074 532667 43077
rect 529828 43072 532667 43074
rect 529828 43016 532606 43072
rect 532662 43016 532667 43072
rect 529828 43014 532667 43016
rect 532601 43011 532667 43014
rect 532601 41714 532667 41717
rect 529828 41712 532667 41714
rect 529828 41656 532606 41712
rect 532662 41656 532667 41712
rect 529828 41654 532667 41656
rect 532601 41651 532667 41654
rect 535453 41714 535519 41717
rect 539200 41714 540000 41744
rect 535453 41712 540000 41714
rect 535453 41656 535458 41712
rect 535514 41656 540000 41712
rect 535453 41654 540000 41656
rect 535453 41651 535519 41654
rect 539200 41624 540000 41654
rect 126973 41442 127039 41445
rect 126973 41440 130180 41442
rect 126973 41384 126978 41440
rect 127034 41384 130180 41440
rect 126973 41382 130180 41384
rect 126973 41379 127039 41382
rect 532601 40218 532667 40221
rect 529828 40216 532667 40218
rect 529828 40160 532606 40216
rect 532662 40160 532667 40216
rect 529828 40158 532667 40160
rect 532601 40155 532667 40158
rect 535453 40218 535519 40221
rect 539200 40218 540000 40248
rect 535453 40216 540000 40218
rect 535453 40160 535458 40216
rect 535514 40160 540000 40216
rect 535453 40158 540000 40160
rect 535453 40155 535519 40158
rect 539200 40128 540000 40158
rect 126973 39538 127039 39541
rect 126973 39536 130180 39538
rect 126973 39480 126978 39536
rect 127034 39480 130180 39536
rect 126973 39478 130180 39480
rect 126973 39475 127039 39478
rect 532601 38858 532667 38861
rect 529828 38856 532667 38858
rect 529828 38800 532606 38856
rect 532662 38800 532667 38856
rect 529828 38798 532667 38800
rect 532601 38795 532667 38798
rect 535453 38722 535519 38725
rect 539200 38722 540000 38752
rect 535453 38720 540000 38722
rect 535453 38664 535458 38720
rect 535514 38664 540000 38720
rect 535453 38662 540000 38664
rect 535453 38659 535519 38662
rect 539200 38632 540000 38662
rect 126973 37634 127039 37637
rect 126973 37632 130180 37634
rect 126973 37576 126978 37632
rect 127034 37576 130180 37632
rect 126973 37574 130180 37576
rect 126973 37571 127039 37574
rect 532601 37498 532667 37501
rect 529828 37496 532667 37498
rect 529828 37440 532606 37496
rect 532662 37440 532667 37496
rect 529828 37438 532667 37440
rect 532601 37435 532667 37438
rect 535361 37226 535427 37229
rect 539200 37226 540000 37256
rect 535361 37224 540000 37226
rect 535361 37168 535366 37224
rect 535422 37168 540000 37224
rect 535361 37166 540000 37168
rect 535361 37163 535427 37166
rect 539200 37136 540000 37166
rect 532325 36138 532391 36141
rect 529828 36136 532391 36138
rect 529828 36080 532330 36136
rect 532386 36080 532391 36136
rect 529828 36078 532391 36080
rect 532325 36075 532391 36078
rect 126329 35730 126395 35733
rect 126329 35728 130180 35730
rect 126329 35672 126334 35728
rect 126390 35672 130180 35728
rect 126329 35670 130180 35672
rect 126329 35667 126395 35670
rect 535361 35594 535427 35597
rect 539200 35594 540000 35624
rect 535361 35592 540000 35594
rect 535361 35536 535366 35592
rect 535422 35536 540000 35592
rect 535361 35534 540000 35536
rect 535361 35531 535427 35534
rect 539200 35504 540000 35534
rect 532601 34778 532667 34781
rect 529828 34776 532667 34778
rect 529828 34720 532606 34776
rect 532662 34720 532667 34776
rect 529828 34718 532667 34720
rect 532601 34715 532667 34718
rect 535361 34098 535427 34101
rect 539200 34098 540000 34128
rect 535361 34096 540000 34098
rect 535361 34040 535366 34096
rect 535422 34040 540000 34096
rect 535361 34038 540000 34040
rect 535361 34035 535427 34038
rect 539200 34008 540000 34038
rect 126973 33690 127039 33693
rect 126973 33688 130180 33690
rect 126973 33632 126978 33688
rect 127034 33632 130180 33688
rect 126973 33630 130180 33632
rect 126973 33627 127039 33630
rect 531957 33418 532023 33421
rect 529828 33416 532023 33418
rect 529828 33360 531962 33416
rect 532018 33360 532023 33416
rect 529828 33358 532023 33360
rect 531957 33355 532023 33358
rect 535361 32602 535427 32605
rect 539200 32602 540000 32632
rect 535361 32600 540000 32602
rect 535361 32544 535366 32600
rect 535422 32544 540000 32600
rect 535361 32542 540000 32544
rect 535361 32539 535427 32542
rect 539200 32512 540000 32542
rect 116853 32330 116919 32333
rect 113804 32328 116919 32330
rect 113804 32272 116858 32328
rect 116914 32272 116919 32328
rect 113804 32270 116919 32272
rect 116853 32267 116919 32270
rect 532601 32058 532667 32061
rect 529828 32056 532667 32058
rect 529828 32000 532606 32056
rect 532662 32000 532667 32056
rect 529828 31998 532667 32000
rect 532601 31995 532667 31998
rect 126973 31786 127039 31789
rect 126973 31784 130180 31786
rect 126973 31728 126978 31784
rect 127034 31728 130180 31784
rect 126973 31726 130180 31728
rect 126973 31723 127039 31726
rect 535361 31106 535427 31109
rect 539200 31106 540000 31136
rect 535361 31104 540000 31106
rect 535361 31048 535366 31104
rect 535422 31048 540000 31104
rect 535361 31046 540000 31048
rect 535361 31043 535427 31046
rect 539200 31016 540000 31046
rect 532601 30698 532667 30701
rect 529828 30696 532667 30698
rect 529828 30640 532606 30696
rect 532662 30640 532667 30696
rect 529828 30638 532667 30640
rect 532601 30635 532667 30638
rect 126973 29882 127039 29885
rect 126973 29880 130180 29882
rect 126973 29824 126978 29880
rect 127034 29824 130180 29880
rect 126973 29822 130180 29824
rect 126973 29819 127039 29822
rect 535361 29610 535427 29613
rect 539200 29610 540000 29640
rect 535361 29608 540000 29610
rect 535361 29552 535366 29608
rect 535422 29552 540000 29608
rect 535361 29550 540000 29552
rect 535361 29547 535427 29550
rect 539200 29520 540000 29550
rect 532601 29338 532667 29341
rect 529828 29336 532667 29338
rect 529828 29280 532606 29336
rect 532662 29280 532667 29336
rect 529828 29278 532667 29280
rect 532601 29275 532667 29278
rect 535361 28114 535427 28117
rect 539200 28114 540000 28144
rect 535361 28112 540000 28114
rect 535361 28056 535366 28112
rect 535422 28056 540000 28112
rect 535361 28054 540000 28056
rect 535361 28051 535427 28054
rect 539200 28024 540000 28054
rect 126973 27978 127039 27981
rect 532601 27978 532667 27981
rect 126973 27976 130180 27978
rect 126973 27920 126978 27976
rect 127034 27920 130180 27976
rect 126973 27918 130180 27920
rect 529828 27976 532667 27978
rect 529828 27920 532606 27976
rect 532662 27920 532667 27976
rect 529828 27918 532667 27920
rect 126973 27915 127039 27918
rect 532601 27915 532667 27918
rect 532325 26618 532391 26621
rect 529828 26616 532391 26618
rect 529828 26560 532330 26616
rect 532386 26560 532391 26616
rect 529828 26558 532391 26560
rect 532325 26555 532391 26558
rect 535453 26482 535519 26485
rect 539200 26482 540000 26512
rect 535453 26480 540000 26482
rect 535453 26424 535458 26480
rect 535514 26424 540000 26480
rect 535453 26422 540000 26424
rect 535453 26419 535519 26422
rect 539200 26392 540000 26422
rect 126973 26074 127039 26077
rect 126973 26072 130180 26074
rect 126973 26016 126978 26072
rect 127034 26016 130180 26072
rect 126973 26014 130180 26016
rect 126973 26011 127039 26014
rect 532601 25258 532667 25261
rect 529828 25256 532667 25258
rect 529828 25200 532606 25256
rect 532662 25200 532667 25256
rect 529828 25198 532667 25200
rect 532601 25195 532667 25198
rect 535361 24986 535427 24989
rect 539200 24986 540000 25016
rect 535361 24984 540000 24986
rect 535361 24928 535366 24984
rect 535422 24928 540000 24984
rect 535361 24926 540000 24928
rect 535361 24923 535427 24926
rect 539200 24896 540000 24926
rect 126421 24170 126487 24173
rect 126421 24168 130180 24170
rect 126421 24112 126426 24168
rect 126482 24112 130180 24168
rect 126421 24110 130180 24112
rect 126421 24107 126487 24110
rect 532049 23898 532115 23901
rect 529828 23896 532115 23898
rect 529828 23840 532054 23896
rect 532110 23840 532115 23896
rect 529828 23838 532115 23840
rect 532049 23835 532115 23838
rect 535361 23490 535427 23493
rect 539200 23490 540000 23520
rect 535361 23488 540000 23490
rect 535361 23432 535366 23488
rect 535422 23432 540000 23488
rect 535361 23430 540000 23432
rect 535361 23427 535427 23430
rect 539200 23400 540000 23430
rect 531957 22402 532023 22405
rect 529828 22400 532023 22402
rect 529828 22344 531962 22400
rect 532018 22344 532023 22400
rect 529828 22342 532023 22344
rect 531957 22339 532023 22342
rect 126973 22266 127039 22269
rect 126973 22264 130180 22266
rect 126973 22208 126978 22264
rect 127034 22208 130180 22264
rect 126973 22206 130180 22208
rect 126973 22203 127039 22206
rect 535269 21994 535335 21997
rect 539200 21994 540000 22024
rect 535269 21992 540000 21994
rect 535269 21936 535274 21992
rect 535330 21936 540000 21992
rect 535269 21934 540000 21936
rect 535269 21931 535335 21934
rect 539200 21904 540000 21934
rect 531957 21042 532023 21045
rect 529828 21040 532023 21042
rect 529828 20984 531962 21040
rect 532018 20984 532023 21040
rect 529828 20982 532023 20984
rect 531957 20979 532023 20982
rect 115933 20906 115999 20909
rect 113804 20904 115999 20906
rect 113804 20848 115938 20904
rect 115994 20848 115999 20904
rect 113804 20846 115999 20848
rect 115933 20843 115999 20846
rect 535361 20498 535427 20501
rect 539200 20498 540000 20528
rect 535361 20496 540000 20498
rect 535361 20440 535366 20496
rect 535422 20440 540000 20496
rect 535361 20438 540000 20440
rect 535361 20435 535427 20438
rect 539200 20408 540000 20438
rect 126973 20362 127039 20365
rect 126973 20360 130180 20362
rect 126973 20304 126978 20360
rect 127034 20304 130180 20360
rect 126973 20302 130180 20304
rect 126973 20299 127039 20302
rect 531957 19682 532023 19685
rect 529828 19680 532023 19682
rect 529828 19624 531962 19680
rect 532018 19624 532023 19680
rect 529828 19622 532023 19624
rect 531957 19619 532023 19622
rect 535269 19002 535335 19005
rect 539200 19002 540000 19032
rect 535269 19000 540000 19002
rect 535269 18944 535274 19000
rect 535330 18944 540000 19000
rect 535269 18942 540000 18944
rect 535269 18939 535335 18942
rect 539200 18912 540000 18942
rect 126973 18322 127039 18325
rect 532325 18322 532391 18325
rect 126973 18320 130180 18322
rect 126973 18264 126978 18320
rect 127034 18264 130180 18320
rect 126973 18262 130180 18264
rect 529828 18320 532391 18322
rect 529828 18264 532330 18320
rect 532386 18264 532391 18320
rect 529828 18262 532391 18264
rect 126973 18259 127039 18262
rect 532325 18259 532391 18262
rect 535177 17370 535243 17373
rect 539200 17370 540000 17400
rect 535177 17368 540000 17370
rect 535177 17312 535182 17368
rect 535238 17312 540000 17368
rect 535177 17310 540000 17312
rect 535177 17307 535243 17310
rect 539200 17280 540000 17310
rect 532233 16962 532299 16965
rect 529828 16960 532299 16962
rect 529828 16904 532238 16960
rect 532294 16904 532299 16960
rect 529828 16902 532299 16904
rect 532233 16899 532299 16902
rect 127249 16418 127315 16421
rect 127249 16416 130180 16418
rect 127249 16360 127254 16416
rect 127310 16360 130180 16416
rect 127249 16358 130180 16360
rect 127249 16355 127315 16358
rect 535361 15874 535427 15877
rect 539200 15874 540000 15904
rect 535361 15872 540000 15874
rect 535361 15816 535366 15872
rect 535422 15816 540000 15872
rect 535361 15814 540000 15816
rect 535361 15811 535427 15814
rect 539200 15784 540000 15814
rect 532601 15602 532667 15605
rect 529828 15600 532667 15602
rect 529828 15544 532606 15600
rect 532662 15544 532667 15600
rect 529828 15542 532667 15544
rect 532601 15539 532667 15542
rect 126973 14514 127039 14517
rect 126973 14512 130180 14514
rect 126973 14456 126978 14512
rect 127034 14456 130180 14512
rect 126973 14454 130180 14456
rect 126973 14451 127039 14454
rect 535269 14378 535335 14381
rect 539200 14378 540000 14408
rect 535269 14376 540000 14378
rect 535269 14320 535274 14376
rect 535330 14320 540000 14376
rect 535269 14318 540000 14320
rect 535269 14315 535335 14318
rect 539200 14288 540000 14318
rect 532141 14242 532207 14245
rect 529828 14240 532207 14242
rect 529828 14184 532146 14240
rect 532202 14184 532207 14240
rect 529828 14182 532207 14184
rect 532141 14179 532207 14182
rect 531589 12882 531655 12885
rect 529828 12880 531655 12882
rect 529828 12824 531594 12880
rect 531650 12824 531655 12880
rect 529828 12822 531655 12824
rect 531589 12819 531655 12822
rect 535361 12882 535427 12885
rect 539200 12882 540000 12912
rect 535361 12880 540000 12882
rect 535361 12824 535366 12880
rect 535422 12824 540000 12880
rect 535361 12822 540000 12824
rect 535361 12819 535427 12822
rect 539200 12792 540000 12822
rect 126973 12610 127039 12613
rect 126973 12608 130180 12610
rect 126973 12552 126978 12608
rect 127034 12552 130180 12608
rect 126973 12550 130180 12552
rect 126973 12547 127039 12550
rect 531957 11522 532023 11525
rect 529828 11520 532023 11522
rect 529828 11464 531962 11520
rect 532018 11464 532023 11520
rect 529828 11462 532023 11464
rect 531957 11459 532023 11462
rect 535269 11386 535335 11389
rect 539200 11386 540000 11416
rect 535269 11384 540000 11386
rect 535269 11328 535274 11384
rect 535330 11328 540000 11384
rect 535269 11326 540000 11328
rect 535269 11323 535335 11326
rect 539200 11296 540000 11326
rect 127709 10706 127775 10709
rect 127709 10704 130180 10706
rect 127709 10648 127714 10704
rect 127770 10648 130180 10704
rect 127709 10646 130180 10648
rect 127709 10643 127775 10646
rect 531773 10162 531839 10165
rect 529828 10160 531839 10162
rect 529828 10104 531778 10160
rect 531834 10104 531839 10160
rect 529828 10102 531839 10104
rect 531773 10099 531839 10102
rect 535361 9890 535427 9893
rect 539200 9890 540000 9920
rect 535361 9888 540000 9890
rect 535361 9832 535366 9888
rect 535422 9832 540000 9888
rect 535361 9830 540000 9832
rect 535361 9827 535427 9830
rect 539200 9800 540000 9830
rect 117221 9618 117287 9621
rect 113804 9616 117287 9618
rect 113804 9560 117226 9616
rect 117282 9560 117287 9616
rect 113804 9558 117287 9560
rect 117221 9555 117287 9558
rect 127801 8802 127867 8805
rect 532233 8802 532299 8805
rect 127801 8800 130180 8802
rect 127801 8744 127806 8800
rect 127862 8744 130180 8800
rect 127801 8742 130180 8744
rect 529828 8800 532299 8802
rect 529828 8744 532238 8800
rect 532294 8744 532299 8800
rect 529828 8742 532299 8744
rect 127801 8739 127867 8742
rect 532233 8739 532299 8742
rect 535177 8258 535243 8261
rect 539200 8258 540000 8288
rect 535177 8256 540000 8258
rect 535177 8200 535182 8256
rect 535238 8200 540000 8256
rect 535177 8198 540000 8200
rect 535177 8195 535243 8198
rect 539200 8168 540000 8198
rect 531957 7442 532023 7445
rect 529828 7440 532023 7442
rect 529828 7384 531962 7440
rect 532018 7384 532023 7440
rect 529828 7382 532023 7384
rect 531957 7379 532023 7382
rect 126973 6898 127039 6901
rect 126973 6896 130180 6898
rect 126973 6840 126978 6896
rect 127034 6840 130180 6896
rect 126973 6838 130180 6840
rect 126973 6835 127039 6838
rect 534993 6762 535059 6765
rect 539200 6762 540000 6792
rect 534993 6760 540000 6762
rect 534993 6704 534998 6760
rect 535054 6704 540000 6760
rect 534993 6702 540000 6704
rect 534993 6699 535059 6702
rect 539200 6672 540000 6702
rect 531589 6082 531655 6085
rect 529828 6080 531655 6082
rect 529828 6024 531594 6080
rect 531650 6024 531655 6080
rect 529828 6022 531655 6024
rect 531589 6019 531655 6022
rect 535269 5266 535335 5269
rect 539200 5266 540000 5296
rect 535269 5264 540000 5266
rect 535269 5208 535274 5264
rect 535330 5208 540000 5264
rect 535269 5206 540000 5208
rect 535269 5203 535335 5206
rect 539200 5176 540000 5206
rect 126973 4994 127039 4997
rect 126973 4992 130180 4994
rect 126973 4936 126978 4992
rect 127034 4936 130180 4992
rect 126973 4934 130180 4936
rect 126973 4931 127039 4934
rect 532601 4722 532667 4725
rect 529828 4720 532667 4722
rect 529828 4664 532606 4720
rect 532662 4664 532667 4720
rect 529828 4662 532667 4664
rect 532601 4659 532667 4662
rect 535177 3770 535243 3773
rect 539200 3770 540000 3800
rect 535177 3768 540000 3770
rect 535177 3712 535182 3768
rect 535238 3712 540000 3768
rect 535177 3710 540000 3712
rect 535177 3707 535243 3710
rect 539200 3680 540000 3710
rect 535361 2274 535427 2277
rect 539200 2274 540000 2304
rect 535361 2272 540000 2274
rect 535361 2216 535366 2272
rect 535422 2216 540000 2272
rect 535361 2214 540000 2216
rect 535361 2211 535427 2214
rect 539200 2184 540000 2214
rect 535453 778 535519 781
rect 539200 778 540000 808
rect 535453 776 540000 778
rect 535453 720 535458 776
rect 535514 720 540000 776
rect 535453 718 540000 720
rect 535453 715 535519 718
rect 539200 688 540000 718
<< via3 >>
rect 49004 158748 49068 158812
rect 164188 157388 164252 157452
<< metal4 >>
rect 164190 157453 164250 158662
rect 164187 157452 164253 157453
rect 164187 157388 164188 157452
rect 164252 157388 164253 157452
rect 164187 157387 164253 157388
<< via4 >>
rect 48918 158812 49154 158898
rect 48918 158748 49004 158812
rect 49004 158748 49068 158812
rect 49068 158748 49154 158812
rect 48918 158662 49154 158748
rect 164102 158662 164338 158898
<< metal5 >>
rect 48876 158898 164380 158940
rect 48876 158662 48918 158898
rect 49154 158662 164102 158898
rect 164338 158662 164380 158898
rect 48876 158620 164380 158662
rect 1104 148346 2000 148666
rect 116000 148346 128000 148666
rect 532000 148346 538844 148666
rect 1104 135346 2000 135666
rect 116000 135346 128000 135666
rect 532000 135346 538844 135666
rect 1104 122346 2000 122666
rect 116000 122346 128000 122666
rect 532000 122346 538844 122666
rect 1104 109346 2000 109666
rect 116000 109346 128000 109666
rect 532000 109346 538844 109666
rect 1104 96346 2000 96666
rect 116000 96346 128000 96666
rect 532000 96346 538844 96666
rect 1104 83346 2000 83666
rect 116000 83346 128000 83666
rect 532000 83346 538844 83666
rect 1104 70346 2000 70666
rect 116000 70346 128000 70666
rect 532000 70346 538844 70666
rect 1104 57346 2000 57666
rect 116000 57346 128000 57666
rect 532000 57346 538844 57666
rect 1104 44346 2000 44666
rect 116000 44346 128000 44666
rect 532000 44346 538844 44666
rect 1104 31346 2000 31666
rect 116000 31346 128000 31666
rect 532000 31346 538844 31666
rect 1104 18346 2000 18666
rect 116000 18346 128000 18666
rect 532000 18346 538844 18666
rect 1104 5346 2000 5666
rect 116000 5346 128000 5666
rect 532000 5346 538844 5666
use mgmt_core  core
timestamp 1636710816
transform 1 0 130000 0 1 4000
box 0 0 400000 148000
use DFFRAM  DFFRAM
timestamp 1636710816
transform 1 0 4000 0 1 4000
box 4 0 110000 148000
<< labels >>
rlabel metal5 s 1104 18346 2000 18666 6 VGND
port 0 nsew ground input
rlabel metal5 s 116000 18346 128000 18666 6 VGND
port 0 nsew ground input
rlabel metal5 s 532000 18346 538844 18666 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 44346 2000 44666 6 VGND
port 0 nsew ground input
rlabel metal5 s 116000 44346 128000 44666 6 VGND
port 0 nsew ground input
rlabel metal5 s 532000 44346 538844 44666 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 70346 2000 70666 6 VGND
port 0 nsew ground input
rlabel metal5 s 116000 70346 128000 70666 6 VGND
port 0 nsew ground input
rlabel metal5 s 532000 70346 538844 70666 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 96346 2000 96666 6 VGND
port 0 nsew ground input
rlabel metal5 s 116000 96346 128000 96666 6 VGND
port 0 nsew ground input
rlabel metal5 s 532000 96346 538844 96666 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 122346 2000 122666 6 VGND
port 0 nsew ground input
rlabel metal5 s 116000 122346 128000 122666 6 VGND
port 0 nsew ground input
rlabel metal5 s 532000 122346 538844 122666 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 148346 2000 148666 6 VGND
port 0 nsew ground input
rlabel metal5 s 116000 148346 128000 148666 6 VGND
port 0 nsew ground input
rlabel metal5 s 532000 148346 538844 148666 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 5346 2000 5666 6 VPWR
port 1 nsew power input
rlabel metal5 s 116000 5346 128000 5666 6 VPWR
port 1 nsew power input
rlabel metal5 s 532000 5346 538844 5666 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 31346 2000 31666 6 VPWR
port 1 nsew power input
rlabel metal5 s 116000 31346 128000 31666 6 VPWR
port 1 nsew power input
rlabel metal5 s 532000 31346 538844 31666 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 57346 2000 57666 6 VPWR
port 1 nsew power input
rlabel metal5 s 116000 57346 128000 57666 6 VPWR
port 1 nsew power input
rlabel metal5 s 532000 57346 538844 57666 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 83346 2000 83666 6 VPWR
port 1 nsew power input
rlabel metal5 s 116000 83346 128000 83666 6 VPWR
port 1 nsew power input
rlabel metal5 s 532000 83346 538844 83666 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 109346 2000 109666 6 VPWR
port 1 nsew power input
rlabel metal5 s 116000 109346 128000 109666 6 VPWR
port 1 nsew power input
rlabel metal5 s 532000 109346 538844 109666 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 135346 2000 135666 6 VPWR
port 1 nsew power input
rlabel metal5 s 116000 135346 128000 135666 6 VPWR
port 1 nsew power input
rlabel metal5 s 532000 135346 538844 135666 6 VPWR
port 1 nsew power input
rlabel metal2 s 506202 0 506258 800 6 core_clk
port 2 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 core_rstn
port 3 nsew signal input
rlabel metal3 s 539200 64472 540000 64592 6 debug_in
port 4 nsew signal input
rlabel metal3 s 539200 65968 540000 66088 6 debug_mode
port 5 nsew signal tristate
rlabel metal3 s 539200 67464 540000 67584 6 debug_oeb
port 6 nsew signal tristate
rlabel metal3 s 539200 68960 540000 69080 6 debug_out
port 7 nsew signal tristate
rlabel metal3 s 539200 144848 540000 144968 6 flash_clk
port 8 nsew signal tristate
rlabel metal3 s 539200 143352 540000 143472 6 flash_csb
port 9 nsew signal tristate
rlabel metal3 s 539200 146480 540000 146600 6 flash_io0_di
port 10 nsew signal input
rlabel metal3 s 539200 147976 540000 148096 6 flash_io0_do
port 11 nsew signal tristate
rlabel metal3 s 539200 149472 540000 149592 6 flash_io0_oeb
port 12 nsew signal tristate
rlabel metal3 s 539200 150968 540000 151088 6 flash_io1_di
port 13 nsew signal input
rlabel metal3 s 539200 152464 540000 152584 6 flash_io1_do
port 14 nsew signal tristate
rlabel metal3 s 539200 153960 540000 154080 6 flash_io1_oeb
port 15 nsew signal tristate
rlabel metal3 s 539200 155592 540000 155712 6 flash_io2_di
port 16 nsew signal input
rlabel metal3 s 539200 157088 540000 157208 6 flash_io2_do
port 17 nsew signal tristate
rlabel metal3 s 539200 158584 540000 158704 6 flash_io2_oeb
port 18 nsew signal tristate
rlabel metal3 s 539200 160080 540000 160200 6 flash_io3_di
port 19 nsew signal input
rlabel metal3 s 539200 161576 540000 161696 6 flash_io3_do
port 20 nsew signal tristate
rlabel metal3 s 539200 163072 540000 163192 6 flash_io3_oeb
port 21 nsew signal tristate
rlabel metal2 s 101126 0 101182 800 6 gpio_in_pad
port 22 nsew signal input
rlabel metal2 s 168654 0 168710 800 6 gpio_inenb_pad
port 23 nsew signal tristate
rlabel metal2 s 236182 0 236238 800 6 gpio_mode0_pad
port 24 nsew signal tristate
rlabel metal2 s 303710 0 303766 800 6 gpio_mode1_pad
port 25 nsew signal tristate
rlabel metal2 s 371146 0 371202 800 6 gpio_out_pad
port 26 nsew signal tristate
rlabel metal2 s 438674 0 438730 800 6 gpio_outenb_pad
port 27 nsew signal tristate
rlabel metal3 s 539200 91808 540000 91928 6 hk_ack_i
port 28 nsew signal input
rlabel metal3 s 539200 94800 540000 94920 6 hk_dat_i[0]
port 29 nsew signal input
rlabel metal3 s 539200 110032 540000 110152 6 hk_dat_i[10]
port 30 nsew signal input
rlabel metal3 s 539200 111528 540000 111648 6 hk_dat_i[11]
port 31 nsew signal input
rlabel metal3 s 539200 113024 540000 113144 6 hk_dat_i[12]
port 32 nsew signal input
rlabel metal3 s 539200 114520 540000 114640 6 hk_dat_i[13]
port 33 nsew signal input
rlabel metal3 s 539200 116016 540000 116136 6 hk_dat_i[14]
port 34 nsew signal input
rlabel metal3 s 539200 117512 540000 117632 6 hk_dat_i[15]
port 35 nsew signal input
rlabel metal3 s 539200 119144 540000 119264 6 hk_dat_i[16]
port 36 nsew signal input
rlabel metal3 s 539200 120640 540000 120760 6 hk_dat_i[17]
port 37 nsew signal input
rlabel metal3 s 539200 122136 540000 122256 6 hk_dat_i[18]
port 38 nsew signal input
rlabel metal3 s 539200 123632 540000 123752 6 hk_dat_i[19]
port 39 nsew signal input
rlabel metal3 s 539200 96296 540000 96416 6 hk_dat_i[1]
port 40 nsew signal input
rlabel metal3 s 539200 125128 540000 125248 6 hk_dat_i[20]
port 41 nsew signal input
rlabel metal3 s 539200 126624 540000 126744 6 hk_dat_i[21]
port 42 nsew signal input
rlabel metal3 s 539200 128256 540000 128376 6 hk_dat_i[22]
port 43 nsew signal input
rlabel metal3 s 539200 129752 540000 129872 6 hk_dat_i[23]
port 44 nsew signal input
rlabel metal3 s 539200 131248 540000 131368 6 hk_dat_i[24]
port 45 nsew signal input
rlabel metal3 s 539200 132744 540000 132864 6 hk_dat_i[25]
port 46 nsew signal input
rlabel metal3 s 539200 134240 540000 134360 6 hk_dat_i[26]
port 47 nsew signal input
rlabel metal3 s 539200 135736 540000 135856 6 hk_dat_i[27]
port 48 nsew signal input
rlabel metal3 s 539200 137368 540000 137488 6 hk_dat_i[28]
port 49 nsew signal input
rlabel metal3 s 539200 138864 540000 138984 6 hk_dat_i[29]
port 50 nsew signal input
rlabel metal3 s 539200 97792 540000 97912 6 hk_dat_i[2]
port 51 nsew signal input
rlabel metal3 s 539200 140360 540000 140480 6 hk_dat_i[30]
port 52 nsew signal input
rlabel metal3 s 539200 141856 540000 141976 6 hk_dat_i[31]
port 53 nsew signal input
rlabel metal3 s 539200 99288 540000 99408 6 hk_dat_i[3]
port 54 nsew signal input
rlabel metal3 s 539200 100920 540000 101040 6 hk_dat_i[4]
port 55 nsew signal input
rlabel metal3 s 539200 102416 540000 102536 6 hk_dat_i[5]
port 56 nsew signal input
rlabel metal3 s 539200 103912 540000 104032 6 hk_dat_i[6]
port 57 nsew signal input
rlabel metal3 s 539200 105408 540000 105528 6 hk_dat_i[7]
port 58 nsew signal input
rlabel metal3 s 539200 106904 540000 107024 6 hk_dat_i[8]
port 59 nsew signal input
rlabel metal3 s 539200 108400 540000 108520 6 hk_dat_i[9]
port 60 nsew signal input
rlabel metal3 s 539200 93304 540000 93424 6 hk_stb_o
port 61 nsew signal tristate
rlabel metal2 s 537758 163200 537814 164000 6 irq[0]
port 62 nsew signal input
rlabel metal2 s 538678 163200 538734 164000 6 irq[1]
port 63 nsew signal input
rlabel metal2 s 539506 163200 539562 164000 6 irq[2]
port 64 nsew signal input
rlabel metal3 s 539200 75080 540000 75200 6 irq[3]
port 65 nsew signal input
rlabel metal3 s 539200 73584 540000 73704 6 irq[4]
port 66 nsew signal input
rlabel metal3 s 539200 71952 540000 72072 6 irq[5]
port 67 nsew signal input
rlabel metal2 s 386 163200 442 164000 6 la_iena[0]
port 68 nsew signal tristate
rlabel metal2 s 347042 163200 347098 164000 6 la_iena[100]
port 69 nsew signal tristate
rlabel metal2 s 350538 163200 350594 164000 6 la_iena[101]
port 70 nsew signal tristate
rlabel metal2 s 354034 163200 354090 164000 6 la_iena[102]
port 71 nsew signal tristate
rlabel metal2 s 357438 163200 357494 164000 6 la_iena[103]
port 72 nsew signal tristate
rlabel metal2 s 360934 163200 360990 164000 6 la_iena[104]
port 73 nsew signal tristate
rlabel metal2 s 364430 163200 364486 164000 6 la_iena[105]
port 74 nsew signal tristate
rlabel metal2 s 367834 163200 367890 164000 6 la_iena[106]
port 75 nsew signal tristate
rlabel metal2 s 371330 163200 371386 164000 6 la_iena[107]
port 76 nsew signal tristate
rlabel metal2 s 374826 163200 374882 164000 6 la_iena[108]
port 77 nsew signal tristate
rlabel metal2 s 378322 163200 378378 164000 6 la_iena[109]
port 78 nsew signal tristate
rlabel metal2 s 34978 163200 35034 164000 6 la_iena[10]
port 79 nsew signal tristate
rlabel metal2 s 381726 163200 381782 164000 6 la_iena[110]
port 80 nsew signal tristate
rlabel metal2 s 385222 163200 385278 164000 6 la_iena[111]
port 81 nsew signal tristate
rlabel metal2 s 388718 163200 388774 164000 6 la_iena[112]
port 82 nsew signal tristate
rlabel metal2 s 392122 163200 392178 164000 6 la_iena[113]
port 83 nsew signal tristate
rlabel metal2 s 395618 163200 395674 164000 6 la_iena[114]
port 84 nsew signal tristate
rlabel metal2 s 399114 163200 399170 164000 6 la_iena[115]
port 85 nsew signal tristate
rlabel metal2 s 402518 163200 402574 164000 6 la_iena[116]
port 86 nsew signal tristate
rlabel metal2 s 406014 163200 406070 164000 6 la_iena[117]
port 87 nsew signal tristate
rlabel metal2 s 409510 163200 409566 164000 6 la_iena[118]
port 88 nsew signal tristate
rlabel metal2 s 412914 163200 412970 164000 6 la_iena[119]
port 89 nsew signal tristate
rlabel metal2 s 38474 163200 38530 164000 6 la_iena[11]
port 90 nsew signal tristate
rlabel metal2 s 416410 163200 416466 164000 6 la_iena[120]
port 91 nsew signal tristate
rlabel metal2 s 419906 163200 419962 164000 6 la_iena[121]
port 92 nsew signal tristate
rlabel metal2 s 423402 163200 423458 164000 6 la_iena[122]
port 93 nsew signal tristate
rlabel metal2 s 426806 163200 426862 164000 6 la_iena[123]
port 94 nsew signal tristate
rlabel metal2 s 430302 163200 430358 164000 6 la_iena[124]
port 95 nsew signal tristate
rlabel metal2 s 433798 163200 433854 164000 6 la_iena[125]
port 96 nsew signal tristate
rlabel metal2 s 437202 163200 437258 164000 6 la_iena[126]
port 97 nsew signal tristate
rlabel metal2 s 440698 163200 440754 164000 6 la_iena[127]
port 98 nsew signal tristate
rlabel metal2 s 41970 163200 42026 164000 6 la_iena[12]
port 99 nsew signal tristate
rlabel metal2 s 45374 163200 45430 164000 6 la_iena[13]
port 100 nsew signal tristate
rlabel metal2 s 48870 163200 48926 164000 6 la_iena[14]
port 101 nsew signal tristate
rlabel metal2 s 52366 163200 52422 164000 6 la_iena[15]
port 102 nsew signal tristate
rlabel metal2 s 55862 163200 55918 164000 6 la_iena[16]
port 103 nsew signal tristate
rlabel metal2 s 59266 163200 59322 164000 6 la_iena[17]
port 104 nsew signal tristate
rlabel metal2 s 62762 163200 62818 164000 6 la_iena[18]
port 105 nsew signal tristate
rlabel metal2 s 66258 163200 66314 164000 6 la_iena[19]
port 106 nsew signal tristate
rlabel metal2 s 3790 163200 3846 164000 6 la_iena[1]
port 107 nsew signal tristate
rlabel metal2 s 69662 163200 69718 164000 6 la_iena[20]
port 108 nsew signal tristate
rlabel metal2 s 73158 163200 73214 164000 6 la_iena[21]
port 109 nsew signal tristate
rlabel metal2 s 76654 163200 76710 164000 6 la_iena[22]
port 110 nsew signal tristate
rlabel metal2 s 80058 163200 80114 164000 6 la_iena[23]
port 111 nsew signal tristate
rlabel metal2 s 83554 163200 83610 164000 6 la_iena[24]
port 112 nsew signal tristate
rlabel metal2 s 87050 163200 87106 164000 6 la_iena[25]
port 113 nsew signal tristate
rlabel metal2 s 90454 163200 90510 164000 6 la_iena[26]
port 114 nsew signal tristate
rlabel metal2 s 93950 163200 94006 164000 6 la_iena[27]
port 115 nsew signal tristate
rlabel metal2 s 97446 163200 97502 164000 6 la_iena[28]
port 116 nsew signal tristate
rlabel metal2 s 100850 163200 100906 164000 6 la_iena[29]
port 117 nsew signal tristate
rlabel metal2 s 7286 163200 7342 164000 6 la_iena[2]
port 118 nsew signal tristate
rlabel metal2 s 104346 163200 104402 164000 6 la_iena[30]
port 119 nsew signal tristate
rlabel metal2 s 107842 163200 107898 164000 6 la_iena[31]
port 120 nsew signal tristate
rlabel metal2 s 111338 163200 111394 164000 6 la_iena[32]
port 121 nsew signal tristate
rlabel metal2 s 114742 163200 114798 164000 6 la_iena[33]
port 122 nsew signal tristate
rlabel metal2 s 118238 163200 118294 164000 6 la_iena[34]
port 123 nsew signal tristate
rlabel metal2 s 121734 163200 121790 164000 6 la_iena[35]
port 124 nsew signal tristate
rlabel metal2 s 125138 163200 125194 164000 6 la_iena[36]
port 125 nsew signal tristate
rlabel metal2 s 128634 163200 128690 164000 6 la_iena[37]
port 126 nsew signal tristate
rlabel metal2 s 132130 163200 132186 164000 6 la_iena[38]
port 127 nsew signal tristate
rlabel metal2 s 135534 163200 135590 164000 6 la_iena[39]
port 128 nsew signal tristate
rlabel metal2 s 10782 163200 10838 164000 6 la_iena[3]
port 129 nsew signal tristate
rlabel metal2 s 139030 163200 139086 164000 6 la_iena[40]
port 130 nsew signal tristate
rlabel metal2 s 142526 163200 142582 164000 6 la_iena[41]
port 131 nsew signal tristate
rlabel metal2 s 145930 163200 145986 164000 6 la_iena[42]
port 132 nsew signal tristate
rlabel metal2 s 149426 163200 149482 164000 6 la_iena[43]
port 133 nsew signal tristate
rlabel metal2 s 152922 163200 152978 164000 6 la_iena[44]
port 134 nsew signal tristate
rlabel metal2 s 156326 163200 156382 164000 6 la_iena[45]
port 135 nsew signal tristate
rlabel metal2 s 159822 163200 159878 164000 6 la_iena[46]
port 136 nsew signal tristate
rlabel metal2 s 163318 163200 163374 164000 6 la_iena[47]
port 137 nsew signal tristate
rlabel metal2 s 166814 163200 166870 164000 6 la_iena[48]
port 138 nsew signal tristate
rlabel metal2 s 170218 163200 170274 164000 6 la_iena[49]
port 139 nsew signal tristate
rlabel metal2 s 14186 163200 14242 164000 6 la_iena[4]
port 140 nsew signal tristate
rlabel metal2 s 173714 163200 173770 164000 6 la_iena[50]
port 141 nsew signal tristate
rlabel metal2 s 177210 163200 177266 164000 6 la_iena[51]
port 142 nsew signal tristate
rlabel metal2 s 180614 163200 180670 164000 6 la_iena[52]
port 143 nsew signal tristate
rlabel metal2 s 184110 163200 184166 164000 6 la_iena[53]
port 144 nsew signal tristate
rlabel metal2 s 187606 163200 187662 164000 6 la_iena[54]
port 145 nsew signal tristate
rlabel metal2 s 191010 163200 191066 164000 6 la_iena[55]
port 146 nsew signal tristate
rlabel metal2 s 194506 163200 194562 164000 6 la_iena[56]
port 147 nsew signal tristate
rlabel metal2 s 198002 163200 198058 164000 6 la_iena[57]
port 148 nsew signal tristate
rlabel metal2 s 201406 163200 201462 164000 6 la_iena[58]
port 149 nsew signal tristate
rlabel metal2 s 204902 163200 204958 164000 6 la_iena[59]
port 150 nsew signal tristate
rlabel metal2 s 17682 163200 17738 164000 6 la_iena[5]
port 151 nsew signal tristate
rlabel metal2 s 208398 163200 208454 164000 6 la_iena[60]
port 152 nsew signal tristate
rlabel metal2 s 211894 163200 211950 164000 6 la_iena[61]
port 153 nsew signal tristate
rlabel metal2 s 215298 163200 215354 164000 6 la_iena[62]
port 154 nsew signal tristate
rlabel metal2 s 218794 163200 218850 164000 6 la_iena[63]
port 155 nsew signal tristate
rlabel metal2 s 222290 163200 222346 164000 6 la_iena[64]
port 156 nsew signal tristate
rlabel metal2 s 225694 163200 225750 164000 6 la_iena[65]
port 157 nsew signal tristate
rlabel metal2 s 229190 163200 229246 164000 6 la_iena[66]
port 158 nsew signal tristate
rlabel metal2 s 232686 163200 232742 164000 6 la_iena[67]
port 159 nsew signal tristate
rlabel metal2 s 236090 163200 236146 164000 6 la_iena[68]
port 160 nsew signal tristate
rlabel metal2 s 239586 163200 239642 164000 6 la_iena[69]
port 161 nsew signal tristate
rlabel metal2 s 21178 163200 21234 164000 6 la_iena[6]
port 162 nsew signal tristate
rlabel metal2 s 243082 163200 243138 164000 6 la_iena[70]
port 163 nsew signal tristate
rlabel metal2 s 246486 163200 246542 164000 6 la_iena[71]
port 164 nsew signal tristate
rlabel metal2 s 249982 163200 250038 164000 6 la_iena[72]
port 165 nsew signal tristate
rlabel metal2 s 253478 163200 253534 164000 6 la_iena[73]
port 166 nsew signal tristate
rlabel metal2 s 256882 163200 256938 164000 6 la_iena[74]
port 167 nsew signal tristate
rlabel metal2 s 260378 163200 260434 164000 6 la_iena[75]
port 168 nsew signal tristate
rlabel metal2 s 263874 163200 263930 164000 6 la_iena[76]
port 169 nsew signal tristate
rlabel metal2 s 267370 163200 267426 164000 6 la_iena[77]
port 170 nsew signal tristate
rlabel metal2 s 270774 163200 270830 164000 6 la_iena[78]
port 171 nsew signal tristate
rlabel metal2 s 274270 163200 274326 164000 6 la_iena[79]
port 172 nsew signal tristate
rlabel metal2 s 24582 163200 24638 164000 6 la_iena[7]
port 173 nsew signal tristate
rlabel metal2 s 277766 163200 277822 164000 6 la_iena[80]
port 174 nsew signal tristate
rlabel metal2 s 281170 163200 281226 164000 6 la_iena[81]
port 175 nsew signal tristate
rlabel metal2 s 284666 163200 284722 164000 6 la_iena[82]
port 176 nsew signal tristate
rlabel metal2 s 288162 163200 288218 164000 6 la_iena[83]
port 177 nsew signal tristate
rlabel metal2 s 291566 163200 291622 164000 6 la_iena[84]
port 178 nsew signal tristate
rlabel metal2 s 295062 163200 295118 164000 6 la_iena[85]
port 179 nsew signal tristate
rlabel metal2 s 298558 163200 298614 164000 6 la_iena[86]
port 180 nsew signal tristate
rlabel metal2 s 301962 163200 302018 164000 6 la_iena[87]
port 181 nsew signal tristate
rlabel metal2 s 305458 163200 305514 164000 6 la_iena[88]
port 182 nsew signal tristate
rlabel metal2 s 308954 163200 309010 164000 6 la_iena[89]
port 183 nsew signal tristate
rlabel metal2 s 28078 163200 28134 164000 6 la_iena[8]
port 184 nsew signal tristate
rlabel metal2 s 312358 163200 312414 164000 6 la_iena[90]
port 185 nsew signal tristate
rlabel metal2 s 315854 163200 315910 164000 6 la_iena[91]
port 186 nsew signal tristate
rlabel metal2 s 319350 163200 319406 164000 6 la_iena[92]
port 187 nsew signal tristate
rlabel metal2 s 322846 163200 322902 164000 6 la_iena[93]
port 188 nsew signal tristate
rlabel metal2 s 326250 163200 326306 164000 6 la_iena[94]
port 189 nsew signal tristate
rlabel metal2 s 329746 163200 329802 164000 6 la_iena[95]
port 190 nsew signal tristate
rlabel metal2 s 333242 163200 333298 164000 6 la_iena[96]
port 191 nsew signal tristate
rlabel metal2 s 336646 163200 336702 164000 6 la_iena[97]
port 192 nsew signal tristate
rlabel metal2 s 340142 163200 340198 164000 6 la_iena[98]
port 193 nsew signal tristate
rlabel metal2 s 343638 163200 343694 164000 6 la_iena[99]
port 194 nsew signal tristate
rlabel metal2 s 31574 163200 31630 164000 6 la_iena[9]
port 195 nsew signal tristate
rlabel metal2 s 1214 163200 1270 164000 6 la_input[0]
port 196 nsew signal input
rlabel metal2 s 347962 163200 348018 164000 6 la_input[100]
port 197 nsew signal input
rlabel metal2 s 351366 163200 351422 164000 6 la_input[101]
port 198 nsew signal input
rlabel metal2 s 354862 163200 354918 164000 6 la_input[102]
port 199 nsew signal input
rlabel metal2 s 358358 163200 358414 164000 6 la_input[103]
port 200 nsew signal input
rlabel metal2 s 361854 163200 361910 164000 6 la_input[104]
port 201 nsew signal input
rlabel metal2 s 365258 163200 365314 164000 6 la_input[105]
port 202 nsew signal input
rlabel metal2 s 368754 163200 368810 164000 6 la_input[106]
port 203 nsew signal input
rlabel metal2 s 372250 163200 372306 164000 6 la_input[107]
port 204 nsew signal input
rlabel metal2 s 375654 163200 375710 164000 6 la_input[108]
port 205 nsew signal input
rlabel metal2 s 379150 163200 379206 164000 6 la_input[109]
port 206 nsew signal input
rlabel metal2 s 35898 163200 35954 164000 6 la_input[10]
port 207 nsew signal input
rlabel metal2 s 382646 163200 382702 164000 6 la_input[110]
port 208 nsew signal input
rlabel metal2 s 386050 163200 386106 164000 6 la_input[111]
port 209 nsew signal input
rlabel metal2 s 389546 163200 389602 164000 6 la_input[112]
port 210 nsew signal input
rlabel metal2 s 393042 163200 393098 164000 6 la_input[113]
port 211 nsew signal input
rlabel metal2 s 396446 163200 396502 164000 6 la_input[114]
port 212 nsew signal input
rlabel metal2 s 399942 163200 399998 164000 6 la_input[115]
port 213 nsew signal input
rlabel metal2 s 403438 163200 403494 164000 6 la_input[116]
port 214 nsew signal input
rlabel metal2 s 406842 163200 406898 164000 6 la_input[117]
port 215 nsew signal input
rlabel metal2 s 410338 163200 410394 164000 6 la_input[118]
port 216 nsew signal input
rlabel metal2 s 413834 163200 413890 164000 6 la_input[119]
port 217 nsew signal input
rlabel metal2 s 39302 163200 39358 164000 6 la_input[11]
port 218 nsew signal input
rlabel metal2 s 417330 163200 417386 164000 6 la_input[120]
port 219 nsew signal input
rlabel metal2 s 420734 163200 420790 164000 6 la_input[121]
port 220 nsew signal input
rlabel metal2 s 424230 163200 424286 164000 6 la_input[122]
port 221 nsew signal input
rlabel metal2 s 427726 163200 427782 164000 6 la_input[123]
port 222 nsew signal input
rlabel metal2 s 431130 163200 431186 164000 6 la_input[124]
port 223 nsew signal input
rlabel metal2 s 434626 163200 434682 164000 6 la_input[125]
port 224 nsew signal input
rlabel metal2 s 438122 163200 438178 164000 6 la_input[126]
port 225 nsew signal input
rlabel metal2 s 441526 163200 441582 164000 6 la_input[127]
port 226 nsew signal input
rlabel metal2 s 42798 163200 42854 164000 6 la_input[12]
port 227 nsew signal input
rlabel metal2 s 46294 163200 46350 164000 6 la_input[13]
port 228 nsew signal input
rlabel metal2 s 49790 163200 49846 164000 6 la_input[14]
port 229 nsew signal input
rlabel metal2 s 53194 163200 53250 164000 6 la_input[15]
port 230 nsew signal input
rlabel metal2 s 56690 163200 56746 164000 6 la_input[16]
port 231 nsew signal input
rlabel metal2 s 60186 163200 60242 164000 6 la_input[17]
port 232 nsew signal input
rlabel metal2 s 63590 163200 63646 164000 6 la_input[18]
port 233 nsew signal input
rlabel metal2 s 67086 163200 67142 164000 6 la_input[19]
port 234 nsew signal input
rlabel metal2 s 4710 163200 4766 164000 6 la_input[1]
port 235 nsew signal input
rlabel metal2 s 70582 163200 70638 164000 6 la_input[20]
port 236 nsew signal input
rlabel metal2 s 73986 163200 74042 164000 6 la_input[21]
port 237 nsew signal input
rlabel metal2 s 77482 163200 77538 164000 6 la_input[22]
port 238 nsew signal input
rlabel metal2 s 80978 163200 81034 164000 6 la_input[23]
port 239 nsew signal input
rlabel metal2 s 84382 163200 84438 164000 6 la_input[24]
port 240 nsew signal input
rlabel metal2 s 87878 163200 87934 164000 6 la_input[25]
port 241 nsew signal input
rlabel metal2 s 91374 163200 91430 164000 6 la_input[26]
port 242 nsew signal input
rlabel metal2 s 94870 163200 94926 164000 6 la_input[27]
port 243 nsew signal input
rlabel metal2 s 98274 163200 98330 164000 6 la_input[28]
port 244 nsew signal input
rlabel metal2 s 101770 163200 101826 164000 6 la_input[29]
port 245 nsew signal input
rlabel metal2 s 8114 163200 8170 164000 6 la_input[2]
port 246 nsew signal input
rlabel metal2 s 105266 163200 105322 164000 6 la_input[30]
port 247 nsew signal input
rlabel metal2 s 108670 163200 108726 164000 6 la_input[31]
port 248 nsew signal input
rlabel metal2 s 112166 163200 112222 164000 6 la_input[32]
port 249 nsew signal input
rlabel metal2 s 115662 163200 115718 164000 6 la_input[33]
port 250 nsew signal input
rlabel metal2 s 119066 163200 119122 164000 6 la_input[34]
port 251 nsew signal input
rlabel metal2 s 122562 163200 122618 164000 6 la_input[35]
port 252 nsew signal input
rlabel metal2 s 126058 163200 126114 164000 6 la_input[36]
port 253 nsew signal input
rlabel metal2 s 129462 163200 129518 164000 6 la_input[37]
port 254 nsew signal input
rlabel metal2 s 132958 163200 133014 164000 6 la_input[38]
port 255 nsew signal input
rlabel metal2 s 136454 163200 136510 164000 6 la_input[39]
port 256 nsew signal input
rlabel metal2 s 11610 163200 11666 164000 6 la_input[3]
port 257 nsew signal input
rlabel metal2 s 139858 163200 139914 164000 6 la_input[40]
port 258 nsew signal input
rlabel metal2 s 143354 163200 143410 164000 6 la_input[41]
port 259 nsew signal input
rlabel metal2 s 146850 163200 146906 164000 6 la_input[42]
port 260 nsew signal input
rlabel metal2 s 150346 163200 150402 164000 6 la_input[43]
port 261 nsew signal input
rlabel metal2 s 153750 163200 153806 164000 6 la_input[44]
port 262 nsew signal input
rlabel metal2 s 157246 163200 157302 164000 6 la_input[45]
port 263 nsew signal input
rlabel metal2 s 160742 163200 160798 164000 6 la_input[46]
port 264 nsew signal input
rlabel metal2 s 164146 163200 164202 164000 6 la_input[47]
port 265 nsew signal input
rlabel metal2 s 167642 163200 167698 164000 6 la_input[48]
port 266 nsew signal input
rlabel metal2 s 171138 163200 171194 164000 6 la_input[49]
port 267 nsew signal input
rlabel metal2 s 15106 163200 15162 164000 6 la_input[4]
port 268 nsew signal input
rlabel metal2 s 174542 163200 174598 164000 6 la_input[50]
port 269 nsew signal input
rlabel metal2 s 178038 163200 178094 164000 6 la_input[51]
port 270 nsew signal input
rlabel metal2 s 181534 163200 181590 164000 6 la_input[52]
port 271 nsew signal input
rlabel metal2 s 184938 163200 184994 164000 6 la_input[53]
port 272 nsew signal input
rlabel metal2 s 188434 163200 188490 164000 6 la_input[54]
port 273 nsew signal input
rlabel metal2 s 191930 163200 191986 164000 6 la_input[55]
port 274 nsew signal input
rlabel metal2 s 195334 163200 195390 164000 6 la_input[56]
port 275 nsew signal input
rlabel metal2 s 198830 163200 198886 164000 6 la_input[57]
port 276 nsew signal input
rlabel metal2 s 202326 163200 202382 164000 6 la_input[58]
port 277 nsew signal input
rlabel metal2 s 205822 163200 205878 164000 6 la_input[59]
port 278 nsew signal input
rlabel metal2 s 18510 163200 18566 164000 6 la_input[5]
port 279 nsew signal input
rlabel metal2 s 209226 163200 209282 164000 6 la_input[60]
port 280 nsew signal input
rlabel metal2 s 212722 163200 212778 164000 6 la_input[61]
port 281 nsew signal input
rlabel metal2 s 216218 163200 216274 164000 6 la_input[62]
port 282 nsew signal input
rlabel metal2 s 219622 163200 219678 164000 6 la_input[63]
port 283 nsew signal input
rlabel metal2 s 223118 163200 223174 164000 6 la_input[64]
port 284 nsew signal input
rlabel metal2 s 226614 163200 226670 164000 6 la_input[65]
port 285 nsew signal input
rlabel metal2 s 230018 163200 230074 164000 6 la_input[66]
port 286 nsew signal input
rlabel metal2 s 233514 163200 233570 164000 6 la_input[67]
port 287 nsew signal input
rlabel metal2 s 237010 163200 237066 164000 6 la_input[68]
port 288 nsew signal input
rlabel metal2 s 240414 163200 240470 164000 6 la_input[69]
port 289 nsew signal input
rlabel metal2 s 22006 163200 22062 164000 6 la_input[6]
port 290 nsew signal input
rlabel metal2 s 243910 163200 243966 164000 6 la_input[70]
port 291 nsew signal input
rlabel metal2 s 247406 163200 247462 164000 6 la_input[71]
port 292 nsew signal input
rlabel metal2 s 250902 163200 250958 164000 6 la_input[72]
port 293 nsew signal input
rlabel metal2 s 254306 163200 254362 164000 6 la_input[73]
port 294 nsew signal input
rlabel metal2 s 257802 163200 257858 164000 6 la_input[74]
port 295 nsew signal input
rlabel metal2 s 261298 163200 261354 164000 6 la_input[75]
port 296 nsew signal input
rlabel metal2 s 264702 163200 264758 164000 6 la_input[76]
port 297 nsew signal input
rlabel metal2 s 268198 163200 268254 164000 6 la_input[77]
port 298 nsew signal input
rlabel metal2 s 271694 163200 271750 164000 6 la_input[78]
port 299 nsew signal input
rlabel metal2 s 275098 163200 275154 164000 6 la_input[79]
port 300 nsew signal input
rlabel metal2 s 25502 163200 25558 164000 6 la_input[7]
port 301 nsew signal input
rlabel metal2 s 278594 163200 278650 164000 6 la_input[80]
port 302 nsew signal input
rlabel metal2 s 282090 163200 282146 164000 6 la_input[81]
port 303 nsew signal input
rlabel metal2 s 285494 163200 285550 164000 6 la_input[82]
port 304 nsew signal input
rlabel metal2 s 288990 163200 289046 164000 6 la_input[83]
port 305 nsew signal input
rlabel metal2 s 292486 163200 292542 164000 6 la_input[84]
port 306 nsew signal input
rlabel metal2 s 295890 163200 295946 164000 6 la_input[85]
port 307 nsew signal input
rlabel metal2 s 299386 163200 299442 164000 6 la_input[86]
port 308 nsew signal input
rlabel metal2 s 302882 163200 302938 164000 6 la_input[87]
port 309 nsew signal input
rlabel metal2 s 306378 163200 306434 164000 6 la_input[88]
port 310 nsew signal input
rlabel metal2 s 309782 163200 309838 164000 6 la_input[89]
port 311 nsew signal input
rlabel metal2 s 28906 163200 28962 164000 6 la_input[8]
port 312 nsew signal input
rlabel metal2 s 313278 163200 313334 164000 6 la_input[90]
port 313 nsew signal input
rlabel metal2 s 316774 163200 316830 164000 6 la_input[91]
port 314 nsew signal input
rlabel metal2 s 320178 163200 320234 164000 6 la_input[92]
port 315 nsew signal input
rlabel metal2 s 323674 163200 323730 164000 6 la_input[93]
port 316 nsew signal input
rlabel metal2 s 327170 163200 327226 164000 6 la_input[94]
port 317 nsew signal input
rlabel metal2 s 330574 163200 330630 164000 6 la_input[95]
port 318 nsew signal input
rlabel metal2 s 334070 163200 334126 164000 6 la_input[96]
port 319 nsew signal input
rlabel metal2 s 337566 163200 337622 164000 6 la_input[97]
port 320 nsew signal input
rlabel metal2 s 340970 163200 341026 164000 6 la_input[98]
port 321 nsew signal input
rlabel metal2 s 344466 163200 344522 164000 6 la_input[99]
port 322 nsew signal input
rlabel metal2 s 32402 163200 32458 164000 6 la_input[9]
port 323 nsew signal input
rlabel metal2 s 2042 163200 2098 164000 6 la_oenb[0]
port 324 nsew signal tristate
rlabel metal2 s 348790 163200 348846 164000 6 la_oenb[100]
port 325 nsew signal tristate
rlabel metal2 s 352286 163200 352342 164000 6 la_oenb[101]
port 326 nsew signal tristate
rlabel metal2 s 355782 163200 355838 164000 6 la_oenb[102]
port 327 nsew signal tristate
rlabel metal2 s 359186 163200 359242 164000 6 la_oenb[103]
port 328 nsew signal tristate
rlabel metal2 s 362682 163200 362738 164000 6 la_oenb[104]
port 329 nsew signal tristate
rlabel metal2 s 366178 163200 366234 164000 6 la_oenb[105]
port 330 nsew signal tristate
rlabel metal2 s 369582 163200 369638 164000 6 la_oenb[106]
port 331 nsew signal tristate
rlabel metal2 s 373078 163200 373134 164000 6 la_oenb[107]
port 332 nsew signal tristate
rlabel metal2 s 376574 163200 376630 164000 6 la_oenb[108]
port 333 nsew signal tristate
rlabel metal2 s 379978 163200 380034 164000 6 la_oenb[109]
port 334 nsew signal tristate
rlabel metal2 s 36726 163200 36782 164000 6 la_oenb[10]
port 335 nsew signal tristate
rlabel metal2 s 383474 163200 383530 164000 6 la_oenb[110]
port 336 nsew signal tristate
rlabel metal2 s 386970 163200 387026 164000 6 la_oenb[111]
port 337 nsew signal tristate
rlabel metal2 s 390374 163200 390430 164000 6 la_oenb[112]
port 338 nsew signal tristate
rlabel metal2 s 393870 163200 393926 164000 6 la_oenb[113]
port 339 nsew signal tristate
rlabel metal2 s 397366 163200 397422 164000 6 la_oenb[114]
port 340 nsew signal tristate
rlabel metal2 s 400862 163200 400918 164000 6 la_oenb[115]
port 341 nsew signal tristate
rlabel metal2 s 404266 163200 404322 164000 6 la_oenb[116]
port 342 nsew signal tristate
rlabel metal2 s 407762 163200 407818 164000 6 la_oenb[117]
port 343 nsew signal tristate
rlabel metal2 s 411258 163200 411314 164000 6 la_oenb[118]
port 344 nsew signal tristate
rlabel metal2 s 414662 163200 414718 164000 6 la_oenb[119]
port 345 nsew signal tristate
rlabel metal2 s 40222 163200 40278 164000 6 la_oenb[11]
port 346 nsew signal tristate
rlabel metal2 s 418158 163200 418214 164000 6 la_oenb[120]
port 347 nsew signal tristate
rlabel metal2 s 421654 163200 421710 164000 6 la_oenb[121]
port 348 nsew signal tristate
rlabel metal2 s 425058 163200 425114 164000 6 la_oenb[122]
port 349 nsew signal tristate
rlabel metal2 s 428554 163200 428610 164000 6 la_oenb[123]
port 350 nsew signal tristate
rlabel metal2 s 432050 163200 432106 164000 6 la_oenb[124]
port 351 nsew signal tristate
rlabel metal2 s 435454 163200 435510 164000 6 la_oenb[125]
port 352 nsew signal tristate
rlabel metal2 s 438950 163200 439006 164000 6 la_oenb[126]
port 353 nsew signal tristate
rlabel metal2 s 442446 163200 442502 164000 6 la_oenb[127]
port 354 nsew signal tristate
rlabel metal2 s 43718 163200 43774 164000 6 la_oenb[12]
port 355 nsew signal tristate
rlabel metal2 s 47122 163200 47178 164000 6 la_oenb[13]
port 356 nsew signal tristate
rlabel metal2 s 50618 163200 50674 164000 6 la_oenb[14]
port 357 nsew signal tristate
rlabel metal2 s 54114 163200 54170 164000 6 la_oenb[15]
port 358 nsew signal tristate
rlabel metal2 s 57518 163200 57574 164000 6 la_oenb[16]
port 359 nsew signal tristate
rlabel metal2 s 61014 163200 61070 164000 6 la_oenb[17]
port 360 nsew signal tristate
rlabel metal2 s 64510 163200 64566 164000 6 la_oenb[18]
port 361 nsew signal tristate
rlabel metal2 s 67914 163200 67970 164000 6 la_oenb[19]
port 362 nsew signal tristate
rlabel metal2 s 5538 163200 5594 164000 6 la_oenb[1]
port 363 nsew signal tristate
rlabel metal2 s 71410 163200 71466 164000 6 la_oenb[20]
port 364 nsew signal tristate
rlabel metal2 s 74906 163200 74962 164000 6 la_oenb[21]
port 365 nsew signal tristate
rlabel metal2 s 78310 163200 78366 164000 6 la_oenb[22]
port 366 nsew signal tristate
rlabel metal2 s 81806 163200 81862 164000 6 la_oenb[23]
port 367 nsew signal tristate
rlabel metal2 s 85302 163200 85358 164000 6 la_oenb[24]
port 368 nsew signal tristate
rlabel metal2 s 88798 163200 88854 164000 6 la_oenb[25]
port 369 nsew signal tristate
rlabel metal2 s 92202 163200 92258 164000 6 la_oenb[26]
port 370 nsew signal tristate
rlabel metal2 s 95698 163200 95754 164000 6 la_oenb[27]
port 371 nsew signal tristate
rlabel metal2 s 99194 163200 99250 164000 6 la_oenb[28]
port 372 nsew signal tristate
rlabel metal2 s 102598 163200 102654 164000 6 la_oenb[29]
port 373 nsew signal tristate
rlabel metal2 s 9034 163200 9090 164000 6 la_oenb[2]
port 374 nsew signal tristate
rlabel metal2 s 106094 163200 106150 164000 6 la_oenb[30]
port 375 nsew signal tristate
rlabel metal2 s 109590 163200 109646 164000 6 la_oenb[31]
port 376 nsew signal tristate
rlabel metal2 s 112994 163200 113050 164000 6 la_oenb[32]
port 377 nsew signal tristate
rlabel metal2 s 116490 163200 116546 164000 6 la_oenb[33]
port 378 nsew signal tristate
rlabel metal2 s 119986 163200 120042 164000 6 la_oenb[34]
port 379 nsew signal tristate
rlabel metal2 s 123390 163200 123446 164000 6 la_oenb[35]
port 380 nsew signal tristate
rlabel metal2 s 126886 163200 126942 164000 6 la_oenb[36]
port 381 nsew signal tristate
rlabel metal2 s 130382 163200 130438 164000 6 la_oenb[37]
port 382 nsew signal tristate
rlabel metal2 s 133878 163200 133934 164000 6 la_oenb[38]
port 383 nsew signal tristate
rlabel metal2 s 137282 163200 137338 164000 6 la_oenb[39]
port 384 nsew signal tristate
rlabel metal2 s 12438 163200 12494 164000 6 la_oenb[3]
port 385 nsew signal tristate
rlabel metal2 s 140778 163200 140834 164000 6 la_oenb[40]
port 386 nsew signal tristate
rlabel metal2 s 144274 163200 144330 164000 6 la_oenb[41]
port 387 nsew signal tristate
rlabel metal2 s 147678 163200 147734 164000 6 la_oenb[42]
port 388 nsew signal tristate
rlabel metal2 s 151174 163200 151230 164000 6 la_oenb[43]
port 389 nsew signal tristate
rlabel metal2 s 154670 163200 154726 164000 6 la_oenb[44]
port 390 nsew signal tristate
rlabel metal2 s 158074 163200 158130 164000 6 la_oenb[45]
port 391 nsew signal tristate
rlabel metal2 s 161570 163200 161626 164000 6 la_oenb[46]
port 392 nsew signal tristate
rlabel metal2 s 165066 163200 165122 164000 6 la_oenb[47]
port 393 nsew signal tristate
rlabel metal2 s 168470 163200 168526 164000 6 la_oenb[48]
port 394 nsew signal tristate
rlabel metal2 s 171966 163200 172022 164000 6 la_oenb[49]
port 395 nsew signal tristate
rlabel metal2 s 15934 163200 15990 164000 6 la_oenb[4]
port 396 nsew signal tristate
rlabel metal2 s 175462 163200 175518 164000 6 la_oenb[50]
port 397 nsew signal tristate
rlabel metal2 s 178866 163200 178922 164000 6 la_oenb[51]
port 398 nsew signal tristate
rlabel metal2 s 182362 163200 182418 164000 6 la_oenb[52]
port 399 nsew signal tristate
rlabel metal2 s 185858 163200 185914 164000 6 la_oenb[53]
port 400 nsew signal tristate
rlabel metal2 s 189354 163200 189410 164000 6 la_oenb[54]
port 401 nsew signal tristate
rlabel metal2 s 192758 163200 192814 164000 6 la_oenb[55]
port 402 nsew signal tristate
rlabel metal2 s 196254 163200 196310 164000 6 la_oenb[56]
port 403 nsew signal tristate
rlabel metal2 s 199750 163200 199806 164000 6 la_oenb[57]
port 404 nsew signal tristate
rlabel metal2 s 203154 163200 203210 164000 6 la_oenb[58]
port 405 nsew signal tristate
rlabel metal2 s 206650 163200 206706 164000 6 la_oenb[59]
port 406 nsew signal tristate
rlabel metal2 s 19430 163200 19486 164000 6 la_oenb[5]
port 407 nsew signal tristate
rlabel metal2 s 210146 163200 210202 164000 6 la_oenb[60]
port 408 nsew signal tristate
rlabel metal2 s 213550 163200 213606 164000 6 la_oenb[61]
port 409 nsew signal tristate
rlabel metal2 s 217046 163200 217102 164000 6 la_oenb[62]
port 410 nsew signal tristate
rlabel metal2 s 220542 163200 220598 164000 6 la_oenb[63]
port 411 nsew signal tristate
rlabel metal2 s 223946 163200 224002 164000 6 la_oenb[64]
port 412 nsew signal tristate
rlabel metal2 s 227442 163200 227498 164000 6 la_oenb[65]
port 413 nsew signal tristate
rlabel metal2 s 230938 163200 230994 164000 6 la_oenb[66]
port 414 nsew signal tristate
rlabel metal2 s 234342 163200 234398 164000 6 la_oenb[67]
port 415 nsew signal tristate
rlabel metal2 s 237838 163200 237894 164000 6 la_oenb[68]
port 416 nsew signal tristate
rlabel metal2 s 241334 163200 241390 164000 6 la_oenb[69]
port 417 nsew signal tristate
rlabel metal2 s 22834 163200 22890 164000 6 la_oenb[6]
port 418 nsew signal tristate
rlabel metal2 s 244830 163200 244886 164000 6 la_oenb[70]
port 419 nsew signal tristate
rlabel metal2 s 248234 163200 248290 164000 6 la_oenb[71]
port 420 nsew signal tristate
rlabel metal2 s 251730 163200 251786 164000 6 la_oenb[72]
port 421 nsew signal tristate
rlabel metal2 s 255226 163200 255282 164000 6 la_oenb[73]
port 422 nsew signal tristate
rlabel metal2 s 258630 163200 258686 164000 6 la_oenb[74]
port 423 nsew signal tristate
rlabel metal2 s 262126 163200 262182 164000 6 la_oenb[75]
port 424 nsew signal tristate
rlabel metal2 s 265622 163200 265678 164000 6 la_oenb[76]
port 425 nsew signal tristate
rlabel metal2 s 269026 163200 269082 164000 6 la_oenb[77]
port 426 nsew signal tristate
rlabel metal2 s 272522 163200 272578 164000 6 la_oenb[78]
port 427 nsew signal tristate
rlabel metal2 s 276018 163200 276074 164000 6 la_oenb[79]
port 428 nsew signal tristate
rlabel metal2 s 26330 163200 26386 164000 6 la_oenb[7]
port 429 nsew signal tristate
rlabel metal2 s 279422 163200 279478 164000 6 la_oenb[80]
port 430 nsew signal tristate
rlabel metal2 s 282918 163200 282974 164000 6 la_oenb[81]
port 431 nsew signal tristate
rlabel metal2 s 286414 163200 286470 164000 6 la_oenb[82]
port 432 nsew signal tristate
rlabel metal2 s 289818 163200 289874 164000 6 la_oenb[83]
port 433 nsew signal tristate
rlabel metal2 s 293314 163200 293370 164000 6 la_oenb[84]
port 434 nsew signal tristate
rlabel metal2 s 296810 163200 296866 164000 6 la_oenb[85]
port 435 nsew signal tristate
rlabel metal2 s 300306 163200 300362 164000 6 la_oenb[86]
port 436 nsew signal tristate
rlabel metal2 s 303710 163200 303766 164000 6 la_oenb[87]
port 437 nsew signal tristate
rlabel metal2 s 307206 163200 307262 164000 6 la_oenb[88]
port 438 nsew signal tristate
rlabel metal2 s 310702 163200 310758 164000 6 la_oenb[89]
port 439 nsew signal tristate
rlabel metal2 s 29826 163200 29882 164000 6 la_oenb[8]
port 440 nsew signal tristate
rlabel metal2 s 314106 163200 314162 164000 6 la_oenb[90]
port 441 nsew signal tristate
rlabel metal2 s 317602 163200 317658 164000 6 la_oenb[91]
port 442 nsew signal tristate
rlabel metal2 s 321098 163200 321154 164000 6 la_oenb[92]
port 443 nsew signal tristate
rlabel metal2 s 324502 163200 324558 164000 6 la_oenb[93]
port 444 nsew signal tristate
rlabel metal2 s 327998 163200 328054 164000 6 la_oenb[94]
port 445 nsew signal tristate
rlabel metal2 s 331494 163200 331550 164000 6 la_oenb[95]
port 446 nsew signal tristate
rlabel metal2 s 334898 163200 334954 164000 6 la_oenb[96]
port 447 nsew signal tristate
rlabel metal2 s 338394 163200 338450 164000 6 la_oenb[97]
port 448 nsew signal tristate
rlabel metal2 s 341890 163200 341946 164000 6 la_oenb[98]
port 449 nsew signal tristate
rlabel metal2 s 345386 163200 345442 164000 6 la_oenb[99]
port 450 nsew signal tristate
rlabel metal2 s 33322 163200 33378 164000 6 la_oenb[9]
port 451 nsew signal tristate
rlabel metal2 s 2962 163200 3018 164000 6 la_output[0]
port 452 nsew signal tristate
rlabel metal2 s 349710 163200 349766 164000 6 la_output[100]
port 453 nsew signal tristate
rlabel metal2 s 353114 163200 353170 164000 6 la_output[101]
port 454 nsew signal tristate
rlabel metal2 s 356610 163200 356666 164000 6 la_output[102]
port 455 nsew signal tristate
rlabel metal2 s 360106 163200 360162 164000 6 la_output[103]
port 456 nsew signal tristate
rlabel metal2 s 363510 163200 363566 164000 6 la_output[104]
port 457 nsew signal tristate
rlabel metal2 s 367006 163200 367062 164000 6 la_output[105]
port 458 nsew signal tristate
rlabel metal2 s 370502 163200 370558 164000 6 la_output[106]
port 459 nsew signal tristate
rlabel metal2 s 373906 163200 373962 164000 6 la_output[107]
port 460 nsew signal tristate
rlabel metal2 s 377402 163200 377458 164000 6 la_output[108]
port 461 nsew signal tristate
rlabel metal2 s 380898 163200 380954 164000 6 la_output[109]
port 462 nsew signal tristate
rlabel metal2 s 37646 163200 37702 164000 6 la_output[10]
port 463 nsew signal tristate
rlabel metal2 s 384394 163200 384450 164000 6 la_output[110]
port 464 nsew signal tristate
rlabel metal2 s 387798 163200 387854 164000 6 la_output[111]
port 465 nsew signal tristate
rlabel metal2 s 391294 163200 391350 164000 6 la_output[112]
port 466 nsew signal tristate
rlabel metal2 s 394790 163200 394846 164000 6 la_output[113]
port 467 nsew signal tristate
rlabel metal2 s 398194 163200 398250 164000 6 la_output[114]
port 468 nsew signal tristate
rlabel metal2 s 401690 163200 401746 164000 6 la_output[115]
port 469 nsew signal tristate
rlabel metal2 s 405186 163200 405242 164000 6 la_output[116]
port 470 nsew signal tristate
rlabel metal2 s 408590 163200 408646 164000 6 la_output[117]
port 471 nsew signal tristate
rlabel metal2 s 412086 163200 412142 164000 6 la_output[118]
port 472 nsew signal tristate
rlabel metal2 s 415582 163200 415638 164000 6 la_output[119]
port 473 nsew signal tristate
rlabel metal2 s 41050 163200 41106 164000 6 la_output[11]
port 474 nsew signal tristate
rlabel metal2 s 418986 163200 419042 164000 6 la_output[120]
port 475 nsew signal tristate
rlabel metal2 s 422482 163200 422538 164000 6 la_output[121]
port 476 nsew signal tristate
rlabel metal2 s 425978 163200 426034 164000 6 la_output[122]
port 477 nsew signal tristate
rlabel metal2 s 429382 163200 429438 164000 6 la_output[123]
port 478 nsew signal tristate
rlabel metal2 s 432878 163200 432934 164000 6 la_output[124]
port 479 nsew signal tristate
rlabel metal2 s 436374 163200 436430 164000 6 la_output[125]
port 480 nsew signal tristate
rlabel metal2 s 439870 163200 439926 164000 6 la_output[126]
port 481 nsew signal tristate
rlabel metal2 s 443274 163200 443330 164000 6 la_output[127]
port 482 nsew signal tristate
rlabel metal2 s 44546 163200 44602 164000 6 la_output[12]
port 483 nsew signal tristate
rlabel metal2 s 48042 163200 48098 164000 6 la_output[13]
port 484 nsew signal tristate
rlabel metal2 s 51446 163200 51502 164000 6 la_output[14]
port 485 nsew signal tristate
rlabel metal2 s 54942 163200 54998 164000 6 la_output[15]
port 486 nsew signal tristate
rlabel metal2 s 58438 163200 58494 164000 6 la_output[16]
port 487 nsew signal tristate
rlabel metal2 s 61842 163200 61898 164000 6 la_output[17]
port 488 nsew signal tristate
rlabel metal2 s 65338 163200 65394 164000 6 la_output[18]
port 489 nsew signal tristate
rlabel metal2 s 68834 163200 68890 164000 6 la_output[19]
port 490 nsew signal tristate
rlabel metal2 s 6366 163200 6422 164000 6 la_output[1]
port 491 nsew signal tristate
rlabel metal2 s 72330 163200 72386 164000 6 la_output[20]
port 492 nsew signal tristate
rlabel metal2 s 75734 163200 75790 164000 6 la_output[21]
port 493 nsew signal tristate
rlabel metal2 s 79230 163200 79286 164000 6 la_output[22]
port 494 nsew signal tristate
rlabel metal2 s 82726 163200 82782 164000 6 la_output[23]
port 495 nsew signal tristate
rlabel metal2 s 86130 163200 86186 164000 6 la_output[24]
port 496 nsew signal tristate
rlabel metal2 s 89626 163200 89682 164000 6 la_output[25]
port 497 nsew signal tristate
rlabel metal2 s 93122 163200 93178 164000 6 la_output[26]
port 498 nsew signal tristate
rlabel metal2 s 96526 163200 96582 164000 6 la_output[27]
port 499 nsew signal tristate
rlabel metal2 s 100022 163200 100078 164000 6 la_output[28]
port 500 nsew signal tristate
rlabel metal2 s 103518 163200 103574 164000 6 la_output[29]
port 501 nsew signal tristate
rlabel metal2 s 9862 163200 9918 164000 6 la_output[2]
port 502 nsew signal tristate
rlabel metal2 s 106922 163200 106978 164000 6 la_output[30]
port 503 nsew signal tristate
rlabel metal2 s 110418 163200 110474 164000 6 la_output[31]
port 504 nsew signal tristate
rlabel metal2 s 113914 163200 113970 164000 6 la_output[32]
port 505 nsew signal tristate
rlabel metal2 s 117318 163200 117374 164000 6 la_output[33]
port 506 nsew signal tristate
rlabel metal2 s 120814 163200 120870 164000 6 la_output[34]
port 507 nsew signal tristate
rlabel metal2 s 124310 163200 124366 164000 6 la_output[35]
port 508 nsew signal tristate
rlabel metal2 s 127806 163200 127862 164000 6 la_output[36]
port 509 nsew signal tristate
rlabel metal2 s 131210 163200 131266 164000 6 la_output[37]
port 510 nsew signal tristate
rlabel metal2 s 134706 163200 134762 164000 6 la_output[38]
port 511 nsew signal tristate
rlabel metal2 s 138202 163200 138258 164000 6 la_output[39]
port 512 nsew signal tristate
rlabel metal2 s 13358 163200 13414 164000 6 la_output[3]
port 513 nsew signal tristate
rlabel metal2 s 141606 163200 141662 164000 6 la_output[40]
port 514 nsew signal tristate
rlabel metal2 s 145102 163200 145158 164000 6 la_output[41]
port 515 nsew signal tristate
rlabel metal2 s 148598 163200 148654 164000 6 la_output[42]
port 516 nsew signal tristate
rlabel metal2 s 152002 163200 152058 164000 6 la_output[43]
port 517 nsew signal tristate
rlabel metal2 s 155498 163200 155554 164000 6 la_output[44]
port 518 nsew signal tristate
rlabel metal2 s 158994 163200 159050 164000 6 la_output[45]
port 519 nsew signal tristate
rlabel metal2 s 162398 163200 162454 164000 6 la_output[46]
port 520 nsew signal tristate
rlabel metal2 s 165894 163200 165950 164000 6 la_output[47]
port 521 nsew signal tristate
rlabel metal2 s 169390 163200 169446 164000 6 la_output[48]
port 522 nsew signal tristate
rlabel metal2 s 172886 163200 172942 164000 6 la_output[49]
port 523 nsew signal tristate
rlabel metal2 s 16854 163200 16910 164000 6 la_output[4]
port 524 nsew signal tristate
rlabel metal2 s 176290 163200 176346 164000 6 la_output[50]
port 525 nsew signal tristate
rlabel metal2 s 179786 163200 179842 164000 6 la_output[51]
port 526 nsew signal tristate
rlabel metal2 s 183282 163200 183338 164000 6 la_output[52]
port 527 nsew signal tristate
rlabel metal2 s 186686 163200 186742 164000 6 la_output[53]
port 528 nsew signal tristate
rlabel metal2 s 190182 163200 190238 164000 6 la_output[54]
port 529 nsew signal tristate
rlabel metal2 s 193678 163200 193734 164000 6 la_output[55]
port 530 nsew signal tristate
rlabel metal2 s 197082 163200 197138 164000 6 la_output[56]
port 531 nsew signal tristate
rlabel metal2 s 200578 163200 200634 164000 6 la_output[57]
port 532 nsew signal tristate
rlabel metal2 s 204074 163200 204130 164000 6 la_output[58]
port 533 nsew signal tristate
rlabel metal2 s 207478 163200 207534 164000 6 la_output[59]
port 534 nsew signal tristate
rlabel metal2 s 20258 163200 20314 164000 6 la_output[5]
port 535 nsew signal tristate
rlabel metal2 s 210974 163200 211030 164000 6 la_output[60]
port 536 nsew signal tristate
rlabel metal2 s 214470 163200 214526 164000 6 la_output[61]
port 537 nsew signal tristate
rlabel metal2 s 217874 163200 217930 164000 6 la_output[62]
port 538 nsew signal tristate
rlabel metal2 s 221370 163200 221426 164000 6 la_output[63]
port 539 nsew signal tristate
rlabel metal2 s 224866 163200 224922 164000 6 la_output[64]
port 540 nsew signal tristate
rlabel metal2 s 228362 163200 228418 164000 6 la_output[65]
port 541 nsew signal tristate
rlabel metal2 s 231766 163200 231822 164000 6 la_output[66]
port 542 nsew signal tristate
rlabel metal2 s 235262 163200 235318 164000 6 la_output[67]
port 543 nsew signal tristate
rlabel metal2 s 238758 163200 238814 164000 6 la_output[68]
port 544 nsew signal tristate
rlabel metal2 s 242162 163200 242218 164000 6 la_output[69]
port 545 nsew signal tristate
rlabel metal2 s 23754 163200 23810 164000 6 la_output[6]
port 546 nsew signal tristate
rlabel metal2 s 245658 163200 245714 164000 6 la_output[70]
port 547 nsew signal tristate
rlabel metal2 s 249154 163200 249210 164000 6 la_output[71]
port 548 nsew signal tristate
rlabel metal2 s 252558 163200 252614 164000 6 la_output[72]
port 549 nsew signal tristate
rlabel metal2 s 256054 163200 256110 164000 6 la_output[73]
port 550 nsew signal tristate
rlabel metal2 s 259550 163200 259606 164000 6 la_output[74]
port 551 nsew signal tristate
rlabel metal2 s 262954 163200 263010 164000 6 la_output[75]
port 552 nsew signal tristate
rlabel metal2 s 266450 163200 266506 164000 6 la_output[76]
port 553 nsew signal tristate
rlabel metal2 s 269946 163200 270002 164000 6 la_output[77]
port 554 nsew signal tristate
rlabel metal2 s 273350 163200 273406 164000 6 la_output[78]
port 555 nsew signal tristate
rlabel metal2 s 276846 163200 276902 164000 6 la_output[79]
port 556 nsew signal tristate
rlabel metal2 s 27250 163200 27306 164000 6 la_output[7]
port 557 nsew signal tristate
rlabel metal2 s 280342 163200 280398 164000 6 la_output[80]
port 558 nsew signal tristate
rlabel metal2 s 283838 163200 283894 164000 6 la_output[81]
port 559 nsew signal tristate
rlabel metal2 s 287242 163200 287298 164000 6 la_output[82]
port 560 nsew signal tristate
rlabel metal2 s 290738 163200 290794 164000 6 la_output[83]
port 561 nsew signal tristate
rlabel metal2 s 294234 163200 294290 164000 6 la_output[84]
port 562 nsew signal tristate
rlabel metal2 s 297638 163200 297694 164000 6 la_output[85]
port 563 nsew signal tristate
rlabel metal2 s 301134 163200 301190 164000 6 la_output[86]
port 564 nsew signal tristate
rlabel metal2 s 304630 163200 304686 164000 6 la_output[87]
port 565 nsew signal tristate
rlabel metal2 s 308034 163200 308090 164000 6 la_output[88]
port 566 nsew signal tristate
rlabel metal2 s 311530 163200 311586 164000 6 la_output[89]
port 567 nsew signal tristate
rlabel metal2 s 30654 163200 30710 164000 6 la_output[8]
port 568 nsew signal tristate
rlabel metal2 s 315026 163200 315082 164000 6 la_output[90]
port 569 nsew signal tristate
rlabel metal2 s 318430 163200 318486 164000 6 la_output[91]
port 570 nsew signal tristate
rlabel metal2 s 321926 163200 321982 164000 6 la_output[92]
port 571 nsew signal tristate
rlabel metal2 s 325422 163200 325478 164000 6 la_output[93]
port 572 nsew signal tristate
rlabel metal2 s 328826 163200 328882 164000 6 la_output[94]
port 573 nsew signal tristate
rlabel metal2 s 332322 163200 332378 164000 6 la_output[95]
port 574 nsew signal tristate
rlabel metal2 s 335818 163200 335874 164000 6 la_output[96]
port 575 nsew signal tristate
rlabel metal2 s 339314 163200 339370 164000 6 la_output[97]
port 576 nsew signal tristate
rlabel metal2 s 342718 163200 342774 164000 6 la_output[98]
port 577 nsew signal tristate
rlabel metal2 s 346214 163200 346270 164000 6 la_output[99]
port 578 nsew signal tristate
rlabel metal2 s 34150 163200 34206 164000 6 la_output[9]
port 579 nsew signal tristate
rlabel metal2 s 444194 163200 444250 164000 6 mprj_ack_i
port 580 nsew signal input
rlabel metal2 s 448518 163200 448574 164000 6 mprj_adr_o[0]
port 581 nsew signal tristate
rlabel metal2 s 477958 163200 478014 164000 6 mprj_adr_o[10]
port 582 nsew signal tristate
rlabel metal2 s 480534 163200 480590 164000 6 mprj_adr_o[11]
port 583 nsew signal tristate
rlabel metal2 s 483202 163200 483258 164000 6 mprj_adr_o[12]
port 584 nsew signal tristate
rlabel metal2 s 485778 163200 485834 164000 6 mprj_adr_o[13]
port 585 nsew signal tristate
rlabel metal2 s 488354 163200 488410 164000 6 mprj_adr_o[14]
port 586 nsew signal tristate
rlabel metal2 s 490930 163200 490986 164000 6 mprj_adr_o[15]
port 587 nsew signal tristate
rlabel metal2 s 493598 163200 493654 164000 6 mprj_adr_o[16]
port 588 nsew signal tristate
rlabel metal2 s 496174 163200 496230 164000 6 mprj_adr_o[17]
port 589 nsew signal tristate
rlabel metal2 s 498750 163200 498806 164000 6 mprj_adr_o[18]
port 590 nsew signal tristate
rlabel metal2 s 501418 163200 501474 164000 6 mprj_adr_o[19]
port 591 nsew signal tristate
rlabel metal2 s 451922 163200 451978 164000 6 mprj_adr_o[1]
port 592 nsew signal tristate
rlabel metal2 s 503994 163200 504050 164000 6 mprj_adr_o[20]
port 593 nsew signal tristate
rlabel metal2 s 506570 163200 506626 164000 6 mprj_adr_o[21]
port 594 nsew signal tristate
rlabel metal2 s 509146 163200 509202 164000 6 mprj_adr_o[22]
port 595 nsew signal tristate
rlabel metal2 s 511814 163200 511870 164000 6 mprj_adr_o[23]
port 596 nsew signal tristate
rlabel metal2 s 514390 163200 514446 164000 6 mprj_adr_o[24]
port 597 nsew signal tristate
rlabel metal2 s 516966 163200 517022 164000 6 mprj_adr_o[25]
port 598 nsew signal tristate
rlabel metal2 s 519542 163200 519598 164000 6 mprj_adr_o[26]
port 599 nsew signal tristate
rlabel metal2 s 522210 163200 522266 164000 6 mprj_adr_o[27]
port 600 nsew signal tristate
rlabel metal2 s 524786 163200 524842 164000 6 mprj_adr_o[28]
port 601 nsew signal tristate
rlabel metal2 s 527362 163200 527418 164000 6 mprj_adr_o[29]
port 602 nsew signal tristate
rlabel metal2 s 455418 163200 455474 164000 6 mprj_adr_o[2]
port 603 nsew signal tristate
rlabel metal2 s 529938 163200 529994 164000 6 mprj_adr_o[30]
port 604 nsew signal tristate
rlabel metal2 s 532606 163200 532662 164000 6 mprj_adr_o[31]
port 605 nsew signal tristate
rlabel metal2 s 458914 163200 458970 164000 6 mprj_adr_o[3]
port 606 nsew signal tristate
rlabel metal2 s 462410 163200 462466 164000 6 mprj_adr_o[4]
port 607 nsew signal tristate
rlabel metal2 s 464986 163200 465042 164000 6 mprj_adr_o[5]
port 608 nsew signal tristate
rlabel metal2 s 467562 163200 467618 164000 6 mprj_adr_o[6]
port 609 nsew signal tristate
rlabel metal2 s 470138 163200 470194 164000 6 mprj_adr_o[7]
port 610 nsew signal tristate
rlabel metal2 s 472806 163200 472862 164000 6 mprj_adr_o[8]
port 611 nsew signal tristate
rlabel metal2 s 475382 163200 475438 164000 6 mprj_adr_o[9]
port 612 nsew signal tristate
rlabel metal2 s 445022 163200 445078 164000 6 mprj_cyc_o
port 613 nsew signal tristate
rlabel metal2 s 449346 163200 449402 164000 6 mprj_dat_i[0]
port 614 nsew signal input
rlabel metal2 s 478878 163200 478934 164000 6 mprj_dat_i[10]
port 615 nsew signal input
rlabel metal2 s 481454 163200 481510 164000 6 mprj_dat_i[11]
port 616 nsew signal input
rlabel metal2 s 484030 163200 484086 164000 6 mprj_dat_i[12]
port 617 nsew signal input
rlabel metal2 s 486606 163200 486662 164000 6 mprj_dat_i[13]
port 618 nsew signal input
rlabel metal2 s 489274 163200 489330 164000 6 mprj_dat_i[14]
port 619 nsew signal input
rlabel metal2 s 491850 163200 491906 164000 6 mprj_dat_i[15]
port 620 nsew signal input
rlabel metal2 s 494426 163200 494482 164000 6 mprj_dat_i[16]
port 621 nsew signal input
rlabel metal2 s 497002 163200 497058 164000 6 mprj_dat_i[17]
port 622 nsew signal input
rlabel metal2 s 499670 163200 499726 164000 6 mprj_dat_i[18]
port 623 nsew signal input
rlabel metal2 s 502246 163200 502302 164000 6 mprj_dat_i[19]
port 624 nsew signal input
rlabel metal2 s 452842 163200 452898 164000 6 mprj_dat_i[1]
port 625 nsew signal input
rlabel metal2 s 504822 163200 504878 164000 6 mprj_dat_i[20]
port 626 nsew signal input
rlabel metal2 s 507398 163200 507454 164000 6 mprj_dat_i[21]
port 627 nsew signal input
rlabel metal2 s 510066 163200 510122 164000 6 mprj_dat_i[22]
port 628 nsew signal input
rlabel metal2 s 512642 163200 512698 164000 6 mprj_dat_i[23]
port 629 nsew signal input
rlabel metal2 s 515218 163200 515274 164000 6 mprj_dat_i[24]
port 630 nsew signal input
rlabel metal2 s 517886 163200 517942 164000 6 mprj_dat_i[25]
port 631 nsew signal input
rlabel metal2 s 520462 163200 520518 164000 6 mprj_dat_i[26]
port 632 nsew signal input
rlabel metal2 s 523038 163200 523094 164000 6 mprj_dat_i[27]
port 633 nsew signal input
rlabel metal2 s 525614 163200 525670 164000 6 mprj_dat_i[28]
port 634 nsew signal input
rlabel metal2 s 528282 163200 528338 164000 6 mprj_dat_i[29]
port 635 nsew signal input
rlabel metal2 s 456338 163200 456394 164000 6 mprj_dat_i[2]
port 636 nsew signal input
rlabel metal2 s 530858 163200 530914 164000 6 mprj_dat_i[30]
port 637 nsew signal input
rlabel metal2 s 533434 163200 533490 164000 6 mprj_dat_i[31]
port 638 nsew signal input
rlabel metal2 s 459742 163200 459798 164000 6 mprj_dat_i[3]
port 639 nsew signal input
rlabel metal2 s 463238 163200 463294 164000 6 mprj_dat_i[4]
port 640 nsew signal input
rlabel metal2 s 465814 163200 465870 164000 6 mprj_dat_i[5]
port 641 nsew signal input
rlabel metal2 s 468390 163200 468446 164000 6 mprj_dat_i[6]
port 642 nsew signal input
rlabel metal2 s 471058 163200 471114 164000 6 mprj_dat_i[7]
port 643 nsew signal input
rlabel metal2 s 473634 163200 473690 164000 6 mprj_dat_i[8]
port 644 nsew signal input
rlabel metal2 s 476210 163200 476266 164000 6 mprj_dat_i[9]
port 645 nsew signal input
rlabel metal2 s 450266 163200 450322 164000 6 mprj_dat_o[0]
port 646 nsew signal tristate
rlabel metal2 s 479706 163200 479762 164000 6 mprj_dat_o[10]
port 647 nsew signal tristate
rlabel metal2 s 482282 163200 482338 164000 6 mprj_dat_o[11]
port 648 nsew signal tristate
rlabel metal2 s 484858 163200 484914 164000 6 mprj_dat_o[12]
port 649 nsew signal tristate
rlabel metal2 s 487526 163200 487582 164000 6 mprj_dat_o[13]
port 650 nsew signal tristate
rlabel metal2 s 490102 163200 490158 164000 6 mprj_dat_o[14]
port 651 nsew signal tristate
rlabel metal2 s 492678 163200 492734 164000 6 mprj_dat_o[15]
port 652 nsew signal tristate
rlabel metal2 s 495346 163200 495402 164000 6 mprj_dat_o[16]
port 653 nsew signal tristate
rlabel metal2 s 497922 163200 497978 164000 6 mprj_dat_o[17]
port 654 nsew signal tristate
rlabel metal2 s 500498 163200 500554 164000 6 mprj_dat_o[18]
port 655 nsew signal tristate
rlabel metal2 s 503074 163200 503130 164000 6 mprj_dat_o[19]
port 656 nsew signal tristate
rlabel metal2 s 453670 163200 453726 164000 6 mprj_dat_o[1]
port 657 nsew signal tristate
rlabel metal2 s 505742 163200 505798 164000 6 mprj_dat_o[20]
port 658 nsew signal tristate
rlabel metal2 s 508318 163200 508374 164000 6 mprj_dat_o[21]
port 659 nsew signal tristate
rlabel metal2 s 510894 163200 510950 164000 6 mprj_dat_o[22]
port 660 nsew signal tristate
rlabel metal2 s 513470 163200 513526 164000 6 mprj_dat_o[23]
port 661 nsew signal tristate
rlabel metal2 s 516138 163200 516194 164000 6 mprj_dat_o[24]
port 662 nsew signal tristate
rlabel metal2 s 518714 163200 518770 164000 6 mprj_dat_o[25]
port 663 nsew signal tristate
rlabel metal2 s 521290 163200 521346 164000 6 mprj_dat_o[26]
port 664 nsew signal tristate
rlabel metal2 s 523866 163200 523922 164000 6 mprj_dat_o[27]
port 665 nsew signal tristate
rlabel metal2 s 526534 163200 526590 164000 6 mprj_dat_o[28]
port 666 nsew signal tristate
rlabel metal2 s 529110 163200 529166 164000 6 mprj_dat_o[29]
port 667 nsew signal tristate
rlabel metal2 s 457166 163200 457222 164000 6 mprj_dat_o[2]
port 668 nsew signal tristate
rlabel metal2 s 531686 163200 531742 164000 6 mprj_dat_o[30]
port 669 nsew signal tristate
rlabel metal2 s 534354 163200 534410 164000 6 mprj_dat_o[31]
port 670 nsew signal tristate
rlabel metal2 s 460662 163200 460718 164000 6 mprj_dat_o[3]
port 671 nsew signal tristate
rlabel metal2 s 464066 163200 464122 164000 6 mprj_dat_o[4]
port 672 nsew signal tristate
rlabel metal2 s 466734 163200 466790 164000 6 mprj_dat_o[5]
port 673 nsew signal tristate
rlabel metal2 s 469310 163200 469366 164000 6 mprj_dat_o[6]
port 674 nsew signal tristate
rlabel metal2 s 471886 163200 471942 164000 6 mprj_dat_o[7]
port 675 nsew signal tristate
rlabel metal2 s 474462 163200 474518 164000 6 mprj_dat_o[8]
port 676 nsew signal tristate
rlabel metal2 s 477130 163200 477186 164000 6 mprj_dat_o[9]
port 677 nsew signal tristate
rlabel metal2 s 451094 163200 451150 164000 6 mprj_sel_o[0]
port 678 nsew signal tristate
rlabel metal2 s 454590 163200 454646 164000 6 mprj_sel_o[1]
port 679 nsew signal tristate
rlabel metal2 s 457994 163200 458050 164000 6 mprj_sel_o[2]
port 680 nsew signal tristate
rlabel metal2 s 461490 163200 461546 164000 6 mprj_sel_o[3]
port 681 nsew signal tristate
rlabel metal2 s 445850 163200 445906 164000 6 mprj_stb_o
port 682 nsew signal tristate
rlabel metal2 s 446770 163200 446826 164000 6 mprj_wb_iena
port 683 nsew signal tristate
rlabel metal2 s 447598 163200 447654 164000 6 mprj_we_o
port 684 nsew signal tristate
rlabel metal3 s 539200 90176 540000 90296 6 qspi_enabled
port 685 nsew signal tristate
rlabel metal3 s 539200 84192 540000 84312 6 ser_rx
port 686 nsew signal input
rlabel metal3 s 539200 85688 540000 85808 6 ser_tx
port 687 nsew signal tristate
rlabel metal3 s 539200 81064 540000 81184 6 spi_csb
port 688 nsew signal tristate
rlabel metal3 s 539200 87184 540000 87304 6 spi_enabled
port 689 nsew signal tristate
rlabel metal3 s 539200 79568 540000 79688 6 spi_sck
port 690 nsew signal tristate
rlabel metal3 s 539200 82696 540000 82816 6 spi_sdi
port 691 nsew signal input
rlabel metal3 s 539200 78072 540000 78192 6 spi_sdo
port 692 nsew signal tristate
rlabel metal3 s 539200 76576 540000 76696 6 spi_sdoenb
port 693 nsew signal tristate
rlabel metal3 s 539200 2184 540000 2304 6 sram_ro_addr[0]
port 694 nsew signal input
rlabel metal3 s 539200 3680 540000 3800 6 sram_ro_addr[1]
port 695 nsew signal input
rlabel metal3 s 539200 5176 540000 5296 6 sram_ro_addr[2]
port 696 nsew signal input
rlabel metal3 s 539200 6672 540000 6792 6 sram_ro_addr[3]
port 697 nsew signal input
rlabel metal3 s 539200 8168 540000 8288 6 sram_ro_addr[4]
port 698 nsew signal input
rlabel metal3 s 539200 9800 540000 9920 6 sram_ro_addr[5]
port 699 nsew signal input
rlabel metal3 s 539200 11296 540000 11416 6 sram_ro_addr[6]
port 700 nsew signal input
rlabel metal3 s 539200 12792 540000 12912 6 sram_ro_addr[7]
port 701 nsew signal input
rlabel metal3 s 539200 14288 540000 14408 6 sram_ro_clk
port 702 nsew signal input
rlabel metal3 s 539200 688 540000 808 6 sram_ro_csb
port 703 nsew signal input
rlabel metal3 s 539200 15784 540000 15904 6 sram_ro_data[0]
port 704 nsew signal tristate
rlabel metal3 s 539200 31016 540000 31136 6 sram_ro_data[10]
port 705 nsew signal tristate
rlabel metal3 s 539200 32512 540000 32632 6 sram_ro_data[11]
port 706 nsew signal tristate
rlabel metal3 s 539200 34008 540000 34128 6 sram_ro_data[12]
port 707 nsew signal tristate
rlabel metal3 s 539200 35504 540000 35624 6 sram_ro_data[13]
port 708 nsew signal tristate
rlabel metal3 s 539200 37136 540000 37256 6 sram_ro_data[14]
port 709 nsew signal tristate
rlabel metal3 s 539200 38632 540000 38752 6 sram_ro_data[15]
port 710 nsew signal tristate
rlabel metal3 s 539200 40128 540000 40248 6 sram_ro_data[16]
port 711 nsew signal tristate
rlabel metal3 s 539200 41624 540000 41744 6 sram_ro_data[17]
port 712 nsew signal tristate
rlabel metal3 s 539200 43120 540000 43240 6 sram_ro_data[18]
port 713 nsew signal tristate
rlabel metal3 s 539200 44616 540000 44736 6 sram_ro_data[19]
port 714 nsew signal tristate
rlabel metal3 s 539200 17280 540000 17400 6 sram_ro_data[1]
port 715 nsew signal tristate
rlabel metal3 s 539200 46248 540000 46368 6 sram_ro_data[20]
port 716 nsew signal tristate
rlabel metal3 s 539200 47744 540000 47864 6 sram_ro_data[21]
port 717 nsew signal tristate
rlabel metal3 s 539200 49240 540000 49360 6 sram_ro_data[22]
port 718 nsew signal tristate
rlabel metal3 s 539200 50736 540000 50856 6 sram_ro_data[23]
port 719 nsew signal tristate
rlabel metal3 s 539200 52232 540000 52352 6 sram_ro_data[24]
port 720 nsew signal tristate
rlabel metal3 s 539200 53728 540000 53848 6 sram_ro_data[25]
port 721 nsew signal tristate
rlabel metal3 s 539200 55360 540000 55480 6 sram_ro_data[26]
port 722 nsew signal tristate
rlabel metal3 s 539200 56856 540000 56976 6 sram_ro_data[27]
port 723 nsew signal tristate
rlabel metal3 s 539200 58352 540000 58472 6 sram_ro_data[28]
port 724 nsew signal tristate
rlabel metal3 s 539200 59848 540000 59968 6 sram_ro_data[29]
port 725 nsew signal tristate
rlabel metal3 s 539200 18912 540000 19032 6 sram_ro_data[2]
port 726 nsew signal tristate
rlabel metal3 s 539200 61344 540000 61464 6 sram_ro_data[30]
port 727 nsew signal tristate
rlabel metal3 s 539200 62840 540000 62960 6 sram_ro_data[31]
port 728 nsew signal tristate
rlabel metal3 s 539200 20408 540000 20528 6 sram_ro_data[3]
port 729 nsew signal tristate
rlabel metal3 s 539200 21904 540000 22024 6 sram_ro_data[4]
port 730 nsew signal tristate
rlabel metal3 s 539200 23400 540000 23520 6 sram_ro_data[5]
port 731 nsew signal tristate
rlabel metal3 s 539200 24896 540000 25016 6 sram_ro_data[6]
port 732 nsew signal tristate
rlabel metal3 s 539200 26392 540000 26512 6 sram_ro_data[7]
port 733 nsew signal tristate
rlabel metal3 s 539200 28024 540000 28144 6 sram_ro_data[8]
port 734 nsew signal tristate
rlabel metal3 s 539200 29520 540000 29640 6 sram_ro_data[9]
port 735 nsew signal tristate
rlabel metal3 s 539200 70456 540000 70576 6 trap
port 736 nsew signal tristate
rlabel metal3 s 539200 88680 540000 88800 6 uart_enabled
port 737 nsew signal tristate
rlabel metal2 s 535182 163200 535238 164000 6 user_irq_ena[0]
port 738 nsew signal tristate
rlabel metal2 s 536010 163200 536066 164000 6 user_irq_ena[1]
port 739 nsew signal tristate
rlabel metal2 s 536930 163200 536986 164000 6 user_irq_ena[2]
port 740 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 540000 164000
<< end >>
